// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 11 2017 17:30:03

// File Generated:     Apr 22 2019 18:24:35

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "Pc2drone" view "INTERFACE"

module Pc2drone (
    uart_input_pc,
    debug_CH5_31B,
    debug_CH3_20A,
    debug_CH0_16A,
    uart_input_drone,
    ppm_output,
    debug_CH6_5B,
    debug_CH2_18A,
    debug_CH4_2A,
    debug_CH1_0A,
    clk_system);

    input uart_input_pc;
    output debug_CH5_31B;
    output debug_CH3_20A;
    output debug_CH0_16A;
    input uart_input_drone;
    output ppm_output;
    output debug_CH6_5B;
    output debug_CH2_18A;
    output debug_CH4_2A;
    output debug_CH1_0A;
    input clk_system;

    wire N__47736;
    wire N__47735;
    wire N__47734;
    wire N__47725;
    wire N__47724;
    wire N__47723;
    wire N__47716;
    wire N__47715;
    wire N__47714;
    wire N__47707;
    wire N__47706;
    wire N__47705;
    wire N__47698;
    wire N__47697;
    wire N__47696;
    wire N__47689;
    wire N__47688;
    wire N__47687;
    wire N__47680;
    wire N__47679;
    wire N__47678;
    wire N__47671;
    wire N__47670;
    wire N__47669;
    wire N__47662;
    wire N__47661;
    wire N__47660;
    wire N__47653;
    wire N__47652;
    wire N__47651;
    wire N__47644;
    wire N__47643;
    wire N__47642;
    wire N__47625;
    wire N__47622;
    wire N__47619;
    wire N__47616;
    wire N__47613;
    wire N__47610;
    wire N__47607;
    wire N__47604;
    wire N__47601;
    wire N__47598;
    wire N__47595;
    wire N__47592;
    wire N__47589;
    wire N__47586;
    wire N__47583;
    wire N__47580;
    wire N__47577;
    wire N__47576;
    wire N__47571;
    wire N__47568;
    wire N__47565;
    wire N__47562;
    wire N__47559;
    wire N__47556;
    wire N__47553;
    wire N__47550;
    wire N__47547;
    wire N__47544;
    wire N__47541;
    wire N__47538;
    wire N__47535;
    wire N__47532;
    wire N__47529;
    wire N__47526;
    wire N__47523;
    wire N__47520;
    wire N__47517;
    wire N__47514;
    wire N__47511;
    wire N__47508;
    wire N__47505;
    wire N__47502;
    wire N__47499;
    wire N__47496;
    wire N__47493;
    wire N__47490;
    wire N__47487;
    wire N__47484;
    wire N__47481;
    wire N__47478;
    wire N__47477;
    wire N__47476;
    wire N__47475;
    wire N__47474;
    wire N__47473;
    wire N__47472;
    wire N__47471;
    wire N__47470;
    wire N__47469;
    wire N__47468;
    wire N__47467;
    wire N__47466;
    wire N__47465;
    wire N__47464;
    wire N__47463;
    wire N__47462;
    wire N__47461;
    wire N__47460;
    wire N__47459;
    wire N__47458;
    wire N__47457;
    wire N__47456;
    wire N__47455;
    wire N__47454;
    wire N__47453;
    wire N__47452;
    wire N__47451;
    wire N__47450;
    wire N__47449;
    wire N__47448;
    wire N__47447;
    wire N__47446;
    wire N__47445;
    wire N__47444;
    wire N__47443;
    wire N__47442;
    wire N__47441;
    wire N__47440;
    wire N__47439;
    wire N__47438;
    wire N__47437;
    wire N__47436;
    wire N__47435;
    wire N__47434;
    wire N__47433;
    wire N__47432;
    wire N__47431;
    wire N__47430;
    wire N__47429;
    wire N__47428;
    wire N__47427;
    wire N__47426;
    wire N__47425;
    wire N__47424;
    wire N__47423;
    wire N__47422;
    wire N__47421;
    wire N__47420;
    wire N__47419;
    wire N__47418;
    wire N__47417;
    wire N__47416;
    wire N__47415;
    wire N__47414;
    wire N__47413;
    wire N__47412;
    wire N__47411;
    wire N__47410;
    wire N__47409;
    wire N__47408;
    wire N__47407;
    wire N__47406;
    wire N__47405;
    wire N__47404;
    wire N__47403;
    wire N__47402;
    wire N__47401;
    wire N__47400;
    wire N__47399;
    wire N__47398;
    wire N__47397;
    wire N__47396;
    wire N__47395;
    wire N__47394;
    wire N__47393;
    wire N__47392;
    wire N__47391;
    wire N__47390;
    wire N__47389;
    wire N__47388;
    wire N__47387;
    wire N__47386;
    wire N__47385;
    wire N__47384;
    wire N__47383;
    wire N__47382;
    wire N__47381;
    wire N__47380;
    wire N__47379;
    wire N__47378;
    wire N__47377;
    wire N__47376;
    wire N__47375;
    wire N__47374;
    wire N__47373;
    wire N__47372;
    wire N__47371;
    wire N__47370;
    wire N__47369;
    wire N__47368;
    wire N__47367;
    wire N__47366;
    wire N__47365;
    wire N__47364;
    wire N__47363;
    wire N__47362;
    wire N__47361;
    wire N__47360;
    wire N__47359;
    wire N__47358;
    wire N__47357;
    wire N__47356;
    wire N__47355;
    wire N__47354;
    wire N__47353;
    wire N__47352;
    wire N__47351;
    wire N__47350;
    wire N__47349;
    wire N__47348;
    wire N__47347;
    wire N__47346;
    wire N__47345;
    wire N__47344;
    wire N__47343;
    wire N__47342;
    wire N__47341;
    wire N__47340;
    wire N__47339;
    wire N__47338;
    wire N__47337;
    wire N__47336;
    wire N__47335;
    wire N__47334;
    wire N__47333;
    wire N__47332;
    wire N__47331;
    wire N__47330;
    wire N__47329;
    wire N__47328;
    wire N__47327;
    wire N__47326;
    wire N__47325;
    wire N__47324;
    wire N__47323;
    wire N__47322;
    wire N__47321;
    wire N__47320;
    wire N__47319;
    wire N__47318;
    wire N__47317;
    wire N__47316;
    wire N__47315;
    wire N__47314;
    wire N__47313;
    wire N__47312;
    wire N__47311;
    wire N__47310;
    wire N__47309;
    wire N__47308;
    wire N__47307;
    wire N__47306;
    wire N__47305;
    wire N__47304;
    wire N__47303;
    wire N__47302;
    wire N__47301;
    wire N__47300;
    wire N__47299;
    wire N__47298;
    wire N__47297;
    wire N__47296;
    wire N__47295;
    wire N__47294;
    wire N__47293;
    wire N__47292;
    wire N__47291;
    wire N__47290;
    wire N__47289;
    wire N__47288;
    wire N__47287;
    wire N__47286;
    wire N__47285;
    wire N__47284;
    wire N__47283;
    wire N__47282;
    wire N__47281;
    wire N__47280;
    wire N__47279;
    wire N__47278;
    wire N__47277;
    wire N__47276;
    wire N__47275;
    wire N__47274;
    wire N__47273;
    wire N__47272;
    wire N__47271;
    wire N__47270;
    wire N__47269;
    wire N__47268;
    wire N__47267;
    wire N__47266;
    wire N__47265;
    wire N__47264;
    wire N__47263;
    wire N__46830;
    wire N__46827;
    wire N__46824;
    wire N__46823;
    wire N__46822;
    wire N__46821;
    wire N__46820;
    wire N__46819;
    wire N__46818;
    wire N__46817;
    wire N__46816;
    wire N__46815;
    wire N__46814;
    wire N__46813;
    wire N__46812;
    wire N__46811;
    wire N__46810;
    wire N__46809;
    wire N__46808;
    wire N__46807;
    wire N__46806;
    wire N__46805;
    wire N__46804;
    wire N__46803;
    wire N__46802;
    wire N__46801;
    wire N__46800;
    wire N__46799;
    wire N__46798;
    wire N__46797;
    wire N__46796;
    wire N__46795;
    wire N__46794;
    wire N__46793;
    wire N__46792;
    wire N__46791;
    wire N__46790;
    wire N__46789;
    wire N__46788;
    wire N__46787;
    wire N__46786;
    wire N__46785;
    wire N__46784;
    wire N__46783;
    wire N__46782;
    wire N__46695;
    wire N__46692;
    wire N__46689;
    wire N__46688;
    wire N__46687;
    wire N__46686;
    wire N__46685;
    wire N__46684;
    wire N__46683;
    wire N__46682;
    wire N__46681;
    wire N__46680;
    wire N__46679;
    wire N__46678;
    wire N__46677;
    wire N__46676;
    wire N__46675;
    wire N__46674;
    wire N__46671;
    wire N__46668;
    wire N__46663;
    wire N__46658;
    wire N__46655;
    wire N__46652;
    wire N__46649;
    wire N__46646;
    wire N__46643;
    wire N__46640;
    wire N__46635;
    wire N__46632;
    wire N__46629;
    wire N__46628;
    wire N__46627;
    wire N__46626;
    wire N__46625;
    wire N__46624;
    wire N__46623;
    wire N__46622;
    wire N__46621;
    wire N__46620;
    wire N__46619;
    wire N__46618;
    wire N__46617;
    wire N__46616;
    wire N__46615;
    wire N__46614;
    wire N__46613;
    wire N__46612;
    wire N__46611;
    wire N__46610;
    wire N__46609;
    wire N__46608;
    wire N__46607;
    wire N__46606;
    wire N__46605;
    wire N__46604;
    wire N__46603;
    wire N__46602;
    wire N__46601;
    wire N__46600;
    wire N__46599;
    wire N__46598;
    wire N__46597;
    wire N__46596;
    wire N__46595;
    wire N__46594;
    wire N__46593;
    wire N__46592;
    wire N__46591;
    wire N__46590;
    wire N__46589;
    wire N__46588;
    wire N__46587;
    wire N__46586;
    wire N__46585;
    wire N__46582;
    wire N__46579;
    wire N__46576;
    wire N__46573;
    wire N__46570;
    wire N__46567;
    wire N__46564;
    wire N__46561;
    wire N__46558;
    wire N__46555;
    wire N__46552;
    wire N__46549;
    wire N__46546;
    wire N__46431;
    wire N__46428;
    wire N__46425;
    wire N__46422;
    wire N__46421;
    wire N__46418;
    wire N__46415;
    wire N__46412;
    wire N__46409;
    wire N__46406;
    wire N__46403;
    wire N__46398;
    wire N__46395;
    wire N__46392;
    wire N__46389;
    wire N__46388;
    wire N__46385;
    wire N__46382;
    wire N__46379;
    wire N__46376;
    wire N__46373;
    wire N__46370;
    wire N__46365;
    wire N__46362;
    wire N__46359;
    wire N__46356;
    wire N__46353;
    wire N__46350;
    wire N__46347;
    wire N__46344;
    wire N__46343;
    wire N__46340;
    wire N__46337;
    wire N__46334;
    wire N__46331;
    wire N__46328;
    wire N__46325;
    wire N__46320;
    wire N__46317;
    wire N__46314;
    wire N__46311;
    wire N__46310;
    wire N__46307;
    wire N__46304;
    wire N__46301;
    wire N__46298;
    wire N__46295;
    wire N__46292;
    wire N__46287;
    wire N__46284;
    wire N__46281;
    wire N__46278;
    wire N__46277;
    wire N__46274;
    wire N__46271;
    wire N__46268;
    wire N__46265;
    wire N__46262;
    wire N__46259;
    wire N__46254;
    wire N__46251;
    wire N__46248;
    wire N__46245;
    wire N__46242;
    wire N__46239;
    wire N__46236;
    wire N__46233;
    wire N__46230;
    wire N__46227;
    wire N__46224;
    wire N__46221;
    wire N__46218;
    wire N__46215;
    wire N__46212;
    wire N__46209;
    wire N__46206;
    wire N__46203;
    wire N__46200;
    wire N__46197;
    wire N__46194;
    wire N__46191;
    wire N__46188;
    wire N__46185;
    wire N__46182;
    wire N__46179;
    wire N__46176;
    wire N__46173;
    wire N__46172;
    wire N__46169;
    wire N__46166;
    wire N__46163;
    wire N__46160;
    wire N__46157;
    wire N__46154;
    wire N__46149;
    wire N__46146;
    wire N__46143;
    wire N__46140;
    wire N__46137;
    wire N__46136;
    wire N__46133;
    wire N__46130;
    wire N__46127;
    wire N__46124;
    wire N__46121;
    wire N__46118;
    wire N__46113;
    wire N__46110;
    wire N__46107;
    wire N__46104;
    wire N__46101;
    wire N__46098;
    wire N__46095;
    wire N__46094;
    wire N__46091;
    wire N__46088;
    wire N__46085;
    wire N__46082;
    wire N__46079;
    wire N__46076;
    wire N__46071;
    wire N__46068;
    wire N__46065;
    wire N__46062;
    wire N__46059;
    wire N__46056;
    wire N__46055;
    wire N__46052;
    wire N__46049;
    wire N__46046;
    wire N__46043;
    wire N__46040;
    wire N__46037;
    wire N__46032;
    wire N__46029;
    wire N__46026;
    wire N__46023;
    wire N__46020;
    wire N__46019;
    wire N__46016;
    wire N__46013;
    wire N__46010;
    wire N__46007;
    wire N__46004;
    wire N__46001;
    wire N__45996;
    wire N__45993;
    wire N__45990;
    wire N__45987;
    wire N__45984;
    wire N__45983;
    wire N__45980;
    wire N__45977;
    wire N__45974;
    wire N__45971;
    wire N__45968;
    wire N__45965;
    wire N__45962;
    wire N__45959;
    wire N__45954;
    wire N__45951;
    wire N__45948;
    wire N__45945;
    wire N__45942;
    wire N__45939;
    wire N__45936;
    wire N__45935;
    wire N__45932;
    wire N__45929;
    wire N__45926;
    wire N__45923;
    wire N__45920;
    wire N__45917;
    wire N__45914;
    wire N__45911;
    wire N__45906;
    wire N__45903;
    wire N__45900;
    wire N__45897;
    wire N__45894;
    wire N__45893;
    wire N__45890;
    wire N__45887;
    wire N__45884;
    wire N__45881;
    wire N__45878;
    wire N__45875;
    wire N__45870;
    wire N__45867;
    wire N__45864;
    wire N__45861;
    wire N__45860;
    wire N__45857;
    wire N__45854;
    wire N__45851;
    wire N__45848;
    wire N__45845;
    wire N__45842;
    wire N__45837;
    wire N__45834;
    wire N__45831;
    wire N__45828;
    wire N__45825;
    wire N__45822;
    wire N__45819;
    wire N__45816;
    wire N__45813;
    wire N__45810;
    wire N__45807;
    wire N__45804;
    wire N__45801;
    wire N__45798;
    wire N__45795;
    wire N__45792;
    wire N__45789;
    wire N__45786;
    wire N__45785;
    wire N__45782;
    wire N__45779;
    wire N__45776;
    wire N__45773;
    wire N__45770;
    wire N__45767;
    wire N__45762;
    wire N__45759;
    wire N__45756;
    wire N__45753;
    wire N__45750;
    wire N__45747;
    wire N__45744;
    wire N__45741;
    wire N__45738;
    wire N__45735;
    wire N__45734;
    wire N__45731;
    wire N__45728;
    wire N__45725;
    wire N__45722;
    wire N__45717;
    wire N__45714;
    wire N__45711;
    wire N__45708;
    wire N__45705;
    wire N__45702;
    wire N__45699;
    wire N__45698;
    wire N__45697;
    wire N__45696;
    wire N__45695;
    wire N__45694;
    wire N__45693;
    wire N__45692;
    wire N__45691;
    wire N__45690;
    wire N__45687;
    wire N__45678;
    wire N__45667;
    wire N__45664;
    wire N__45659;
    wire N__45656;
    wire N__45653;
    wire N__45650;
    wire N__45647;
    wire N__45644;
    wire N__45641;
    wire N__45636;
    wire N__45635;
    wire N__45634;
    wire N__45633;
    wire N__45632;
    wire N__45631;
    wire N__45630;
    wire N__45629;
    wire N__45628;
    wire N__45619;
    wire N__45608;
    wire N__45603;
    wire N__45600;
    wire N__45597;
    wire N__45596;
    wire N__45593;
    wire N__45590;
    wire N__45587;
    wire N__45584;
    wire N__45581;
    wire N__45578;
    wire N__45575;
    wire N__45572;
    wire N__45567;
    wire N__45564;
    wire N__45561;
    wire N__45558;
    wire N__45557;
    wire N__45554;
    wire N__45551;
    wire N__45548;
    wire N__45545;
    wire N__45542;
    wire N__45539;
    wire N__45534;
    wire N__45531;
    wire N__45528;
    wire N__45525;
    wire N__45522;
    wire N__45519;
    wire N__45516;
    wire N__45513;
    wire N__45510;
    wire N__45507;
    wire N__45504;
    wire N__45501;
    wire N__45498;
    wire N__45495;
    wire N__45494;
    wire N__45493;
    wire N__45490;
    wire N__45485;
    wire N__45482;
    wire N__45479;
    wire N__45476;
    wire N__45473;
    wire N__45468;
    wire N__45465;
    wire N__45462;
    wire N__45459;
    wire N__45456;
    wire N__45453;
    wire N__45452;
    wire N__45449;
    wire N__45446;
    wire N__45443;
    wire N__45440;
    wire N__45437;
    wire N__45434;
    wire N__45429;
    wire N__45426;
    wire N__45423;
    wire N__45420;
    wire N__45417;
    wire N__45414;
    wire N__45411;
    wire N__45408;
    wire N__45405;
    wire N__45402;
    wire N__45399;
    wire N__45396;
    wire N__45393;
    wire N__45390;
    wire N__45387;
    wire N__45384;
    wire N__45381;
    wire N__45378;
    wire N__45375;
    wire N__45372;
    wire N__45369;
    wire N__45366;
    wire N__45363;
    wire N__45362;
    wire N__45359;
    wire N__45358;
    wire N__45355;
    wire N__45352;
    wire N__45351;
    wire N__45350;
    wire N__45347;
    wire N__45344;
    wire N__45341;
    wire N__45338;
    wire N__45335;
    wire N__45332;
    wire N__45331;
    wire N__45330;
    wire N__45327;
    wire N__45324;
    wire N__45321;
    wire N__45318;
    wire N__45315;
    wire N__45314;
    wire N__45313;
    wire N__45310;
    wire N__45307;
    wire N__45302;
    wire N__45299;
    wire N__45298;
    wire N__45297;
    wire N__45296;
    wire N__45293;
    wire N__45290;
    wire N__45287;
    wire N__45284;
    wire N__45275;
    wire N__45274;
    wire N__45271;
    wire N__45268;
    wire N__45265;
    wire N__45260;
    wire N__45253;
    wire N__45250;
    wire N__45237;
    wire N__45234;
    wire N__45231;
    wire N__45228;
    wire N__45225;
    wire N__45224;
    wire N__45221;
    wire N__45218;
    wire N__45215;
    wire N__45214;
    wire N__45213;
    wire N__45212;
    wire N__45211;
    wire N__45208;
    wire N__45205;
    wire N__45204;
    wire N__45201;
    wire N__45200;
    wire N__45197;
    wire N__45194;
    wire N__45191;
    wire N__45190;
    wire N__45187;
    wire N__45186;
    wire N__45183;
    wire N__45180;
    wire N__45177;
    wire N__45176;
    wire N__45173;
    wire N__45168;
    wire N__45165;
    wire N__45162;
    wire N__45161;
    wire N__45158;
    wire N__45155;
    wire N__45150;
    wire N__45147;
    wire N__45144;
    wire N__45141;
    wire N__45134;
    wire N__45131;
    wire N__45130;
    wire N__45127;
    wire N__45124;
    wire N__45121;
    wire N__45118;
    wire N__45115;
    wire N__45112;
    wire N__45109;
    wire N__45106;
    wire N__45103;
    wire N__45096;
    wire N__45091;
    wire N__45078;
    wire N__45075;
    wire N__45072;
    wire N__45069;
    wire N__45066;
    wire N__45063;
    wire N__45060;
    wire N__45057;
    wire N__45054;
    wire N__45051;
    wire N__45050;
    wire N__45047;
    wire N__45044;
    wire N__45041;
    wire N__45038;
    wire N__45033;
    wire N__45030;
    wire N__45027;
    wire N__45024;
    wire N__45021;
    wire N__45018;
    wire N__45015;
    wire N__45014;
    wire N__45013;
    wire N__45012;
    wire N__45009;
    wire N__45006;
    wire N__45005;
    wire N__45002;
    wire N__45001;
    wire N__44998;
    wire N__44995;
    wire N__44992;
    wire N__44989;
    wire N__44988;
    wire N__44985;
    wire N__44984;
    wire N__44983;
    wire N__44982;
    wire N__44979;
    wire N__44976;
    wire N__44973;
    wire N__44970;
    wire N__44967;
    wire N__44964;
    wire N__44961;
    wire N__44958;
    wire N__44955;
    wire N__44954;
    wire N__44953;
    wire N__44950;
    wire N__44947;
    wire N__44946;
    wire N__44941;
    wire N__44934;
    wire N__44931;
    wire N__44926;
    wire N__44923;
    wire N__44920;
    wire N__44915;
    wire N__44914;
    wire N__44911;
    wire N__44908;
    wire N__44903;
    wire N__44898;
    wire N__44893;
    wire N__44890;
    wire N__44877;
    wire N__44874;
    wire N__44871;
    wire N__44868;
    wire N__44865;
    wire N__44864;
    wire N__44861;
    wire N__44860;
    wire N__44857;
    wire N__44856;
    wire N__44853;
    wire N__44850;
    wire N__44849;
    wire N__44846;
    wire N__44843;
    wire N__44838;
    wire N__44835;
    wire N__44832;
    wire N__44829;
    wire N__44828;
    wire N__44825;
    wire N__44822;
    wire N__44821;
    wire N__44816;
    wire N__44813;
    wire N__44808;
    wire N__44805;
    wire N__44800;
    wire N__44795;
    wire N__44792;
    wire N__44789;
    wire N__44786;
    wire N__44783;
    wire N__44780;
    wire N__44777;
    wire N__44772;
    wire N__44769;
    wire N__44766;
    wire N__44763;
    wire N__44760;
    wire N__44757;
    wire N__44754;
    wire N__44751;
    wire N__44748;
    wire N__44745;
    wire N__44742;
    wire N__44739;
    wire N__44736;
    wire N__44733;
    wire N__44730;
    wire N__44727;
    wire N__44724;
    wire N__44721;
    wire N__44718;
    wire N__44715;
    wire N__44712;
    wire N__44709;
    wire N__44706;
    wire N__44703;
    wire N__44700;
    wire N__44697;
    wire N__44694;
    wire N__44691;
    wire N__44688;
    wire N__44685;
    wire N__44682;
    wire N__44679;
    wire N__44676;
    wire N__44673;
    wire N__44670;
    wire N__44667;
    wire N__44666;
    wire N__44665;
    wire N__44662;
    wire N__44661;
    wire N__44656;
    wire N__44653;
    wire N__44650;
    wire N__44647;
    wire N__44642;
    wire N__44639;
    wire N__44634;
    wire N__44631;
    wire N__44628;
    wire N__44625;
    wire N__44622;
    wire N__44621;
    wire N__44620;
    wire N__44617;
    wire N__44614;
    wire N__44611;
    wire N__44608;
    wire N__44601;
    wire N__44598;
    wire N__44595;
    wire N__44592;
    wire N__44589;
    wire N__44586;
    wire N__44585;
    wire N__44584;
    wire N__44581;
    wire N__44578;
    wire N__44575;
    wire N__44572;
    wire N__44565;
    wire N__44562;
    wire N__44559;
    wire N__44556;
    wire N__44553;
    wire N__44552;
    wire N__44549;
    wire N__44548;
    wire N__44545;
    wire N__44542;
    wire N__44541;
    wire N__44540;
    wire N__44539;
    wire N__44538;
    wire N__44537;
    wire N__44532;
    wire N__44529;
    wire N__44526;
    wire N__44523;
    wire N__44520;
    wire N__44515;
    wire N__44512;
    wire N__44499;
    wire N__44496;
    wire N__44495;
    wire N__44492;
    wire N__44489;
    wire N__44486;
    wire N__44485;
    wire N__44482;
    wire N__44479;
    wire N__44476;
    wire N__44469;
    wire N__44468;
    wire N__44465;
    wire N__44462;
    wire N__44461;
    wire N__44458;
    wire N__44455;
    wire N__44452;
    wire N__44451;
    wire N__44448;
    wire N__44445;
    wire N__44442;
    wire N__44439;
    wire N__44436;
    wire N__44429;
    wire N__44424;
    wire N__44423;
    wire N__44422;
    wire N__44421;
    wire N__44420;
    wire N__44415;
    wire N__44410;
    wire N__44407;
    wire N__44406;
    wire N__44405;
    wire N__44398;
    wire N__44393;
    wire N__44392;
    wire N__44391;
    wire N__44386;
    wire N__44383;
    wire N__44382;
    wire N__44379;
    wire N__44378;
    wire N__44375;
    wire N__44372;
    wire N__44369;
    wire N__44366;
    wire N__44363;
    wire N__44360;
    wire N__44355;
    wire N__44352;
    wire N__44343;
    wire N__44340;
    wire N__44337;
    wire N__44334;
    wire N__44331;
    wire N__44330;
    wire N__44327;
    wire N__44324;
    wire N__44321;
    wire N__44318;
    wire N__44313;
    wire N__44310;
    wire N__44307;
    wire N__44304;
    wire N__44301;
    wire N__44298;
    wire N__44295;
    wire N__44292;
    wire N__44291;
    wire N__44290;
    wire N__44287;
    wire N__44284;
    wire N__44283;
    wire N__44280;
    wire N__44275;
    wire N__44272;
    wire N__44271;
    wire N__44270;
    wire N__44267;
    wire N__44264;
    wire N__44263;
    wire N__44262;
    wire N__44259;
    wire N__44258;
    wire N__44255;
    wire N__44254;
    wire N__44251;
    wire N__44250;
    wire N__44249;
    wire N__44244;
    wire N__44241;
    wire N__44240;
    wire N__44237;
    wire N__44234;
    wire N__44227;
    wire N__44224;
    wire N__44221;
    wire N__44218;
    wire N__44213;
    wire N__44210;
    wire N__44207;
    wire N__44206;
    wire N__44205;
    wire N__44202;
    wire N__44199;
    wire N__44190;
    wire N__44187;
    wire N__44184;
    wire N__44181;
    wire N__44178;
    wire N__44175;
    wire N__44172;
    wire N__44169;
    wire N__44154;
    wire N__44151;
    wire N__44148;
    wire N__44145;
    wire N__44142;
    wire N__44139;
    wire N__44138;
    wire N__44137;
    wire N__44136;
    wire N__44135;
    wire N__44132;
    wire N__44129;
    wire N__44128;
    wire N__44127;
    wire N__44126;
    wire N__44125;
    wire N__44124;
    wire N__44123;
    wire N__44122;
    wire N__44119;
    wire N__44118;
    wire N__44117;
    wire N__44116;
    wire N__44113;
    wire N__44112;
    wire N__44111;
    wire N__44110;
    wire N__44109;
    wire N__44108;
    wire N__44107;
    wire N__44106;
    wire N__44105;
    wire N__44104;
    wire N__44103;
    wire N__44102;
    wire N__44101;
    wire N__44100;
    wire N__44099;
    wire N__44098;
    wire N__44097;
    wire N__44096;
    wire N__44093;
    wire N__44092;
    wire N__44091;
    wire N__44090;
    wire N__44089;
    wire N__44088;
    wire N__44087;
    wire N__44086;
    wire N__44085;
    wire N__44084;
    wire N__44083;
    wire N__44082;
    wire N__44081;
    wire N__44080;
    wire N__44079;
    wire N__44078;
    wire N__44077;
    wire N__44076;
    wire N__44075;
    wire N__44074;
    wire N__44073;
    wire N__44072;
    wire N__44071;
    wire N__44070;
    wire N__44069;
    wire N__44068;
    wire N__44067;
    wire N__44066;
    wire N__44065;
    wire N__44060;
    wire N__44057;
    wire N__44052;
    wire N__44049;
    wire N__44046;
    wire N__44043;
    wire N__44040;
    wire N__44037;
    wire N__44034;
    wire N__44031;
    wire N__44022;
    wire N__44019;
    wire N__44014;
    wire N__44009;
    wire N__44004;
    wire N__43999;
    wire N__43996;
    wire N__43993;
    wire N__43990;
    wire N__43983;
    wire N__43980;
    wire N__43977;
    wire N__43974;
    wire N__43971;
    wire N__43968;
    wire N__43965;
    wire N__43960;
    wire N__43957;
    wire N__43954;
    wire N__43951;
    wire N__43948;
    wire N__43941;
    wire N__43938;
    wire N__43933;
    wire N__43930;
    wire N__43927;
    wire N__43922;
    wire N__43919;
    wire N__43916;
    wire N__43913;
    wire N__43908;
    wire N__43905;
    wire N__43902;
    wire N__43901;
    wire N__43900;
    wire N__43899;
    wire N__43898;
    wire N__43897;
    wire N__43896;
    wire N__43895;
    wire N__43894;
    wire N__43893;
    wire N__43892;
    wire N__43891;
    wire N__43890;
    wire N__43889;
    wire N__43888;
    wire N__43887;
    wire N__43886;
    wire N__43885;
    wire N__43884;
    wire N__43883;
    wire N__43882;
    wire N__43881;
    wire N__43880;
    wire N__43879;
    wire N__43878;
    wire N__43877;
    wire N__43876;
    wire N__43875;
    wire N__43874;
    wire N__43873;
    wire N__43872;
    wire N__43871;
    wire N__43870;
    wire N__43869;
    wire N__43868;
    wire N__43867;
    wire N__43866;
    wire N__43865;
    wire N__43864;
    wire N__43863;
    wire N__43862;
    wire N__43861;
    wire N__43860;
    wire N__43859;
    wire N__43858;
    wire N__43857;
    wire N__43856;
    wire N__43855;
    wire N__43854;
    wire N__43853;
    wire N__43852;
    wire N__43851;
    wire N__43850;
    wire N__43849;
    wire N__43848;
    wire N__43847;
    wire N__43846;
    wire N__43845;
    wire N__43844;
    wire N__43843;
    wire N__43842;
    wire N__43841;
    wire N__43840;
    wire N__43839;
    wire N__43838;
    wire N__43837;
    wire N__43836;
    wire N__43835;
    wire N__43834;
    wire N__43833;
    wire N__43832;
    wire N__43831;
    wire N__43830;
    wire N__43829;
    wire N__43828;
    wire N__43827;
    wire N__43826;
    wire N__43825;
    wire N__43824;
    wire N__43823;
    wire N__43822;
    wire N__43821;
    wire N__43820;
    wire N__43819;
    wire N__43818;
    wire N__43817;
    wire N__43816;
    wire N__43815;
    wire N__43814;
    wire N__43813;
    wire N__43812;
    wire N__43811;
    wire N__43810;
    wire N__43809;
    wire N__43808;
    wire N__43807;
    wire N__43806;
    wire N__43805;
    wire N__43804;
    wire N__43803;
    wire N__43802;
    wire N__43801;
    wire N__43800;
    wire N__43799;
    wire N__43796;
    wire N__43793;
    wire N__43790;
    wire N__43787;
    wire N__43784;
    wire N__43781;
    wire N__43778;
    wire N__43775;
    wire N__43772;
    wire N__43769;
    wire N__43766;
    wire N__43763;
    wire N__43760;
    wire N__43757;
    wire N__43754;
    wire N__43751;
    wire N__43748;
    wire N__43745;
    wire N__43742;
    wire N__43739;
    wire N__43736;
    wire N__43733;
    wire N__43730;
    wire N__43727;
    wire N__43724;
    wire N__43721;
    wire N__43718;
    wire N__43715;
    wire N__43712;
    wire N__43709;
    wire N__43706;
    wire N__43703;
    wire N__43700;
    wire N__43697;
    wire N__43694;
    wire N__43691;
    wire N__43688;
    wire N__43685;
    wire N__43682;
    wire N__43679;
    wire N__43676;
    wire N__43673;
    wire N__43670;
    wire N__43377;
    wire N__43374;
    wire N__43371;
    wire N__43368;
    wire N__43365;
    wire N__43364;
    wire N__43361;
    wire N__43358;
    wire N__43355;
    wire N__43354;
    wire N__43353;
    wire N__43350;
    wire N__43349;
    wire N__43346;
    wire N__43343;
    wire N__43342;
    wire N__43341;
    wire N__43340;
    wire N__43339;
    wire N__43336;
    wire N__43333;
    wire N__43330;
    wire N__43325;
    wire N__43322;
    wire N__43319;
    wire N__43316;
    wire N__43313;
    wire N__43312;
    wire N__43309;
    wire N__43308;
    wire N__43305;
    wire N__43298;
    wire N__43293;
    wire N__43290;
    wire N__43287;
    wire N__43286;
    wire N__43283;
    wire N__43280;
    wire N__43277;
    wire N__43274;
    wire N__43267;
    wire N__43266;
    wire N__43263;
    wire N__43258;
    wire N__43253;
    wire N__43250;
    wire N__43247;
    wire N__43244;
    wire N__43239;
    wire N__43230;
    wire N__43227;
    wire N__43224;
    wire N__43221;
    wire N__43218;
    wire N__43215;
    wire N__43212;
    wire N__43209;
    wire N__43206;
    wire N__43203;
    wire N__43200;
    wire N__43197;
    wire N__43194;
    wire N__43191;
    wire N__43188;
    wire N__43185;
    wire N__43182;
    wire N__43179;
    wire N__43176;
    wire N__43173;
    wire N__43170;
    wire N__43167;
    wire N__43164;
    wire N__43161;
    wire N__43158;
    wire N__43155;
    wire N__43152;
    wire N__43149;
    wire N__43146;
    wire N__43143;
    wire N__43140;
    wire N__43139;
    wire N__43138;
    wire N__43135;
    wire N__43132;
    wire N__43131;
    wire N__43130;
    wire N__43129;
    wire N__43128;
    wire N__43127;
    wire N__43126;
    wire N__43125;
    wire N__43124;
    wire N__43123;
    wire N__43122;
    wire N__43119;
    wire N__43118;
    wire N__43117;
    wire N__43116;
    wire N__43111;
    wire N__43110;
    wire N__43107;
    wire N__43104;
    wire N__43101;
    wire N__43098;
    wire N__43093;
    wire N__43088;
    wire N__43087;
    wire N__43086;
    wire N__43085;
    wire N__43082;
    wire N__43081;
    wire N__43078;
    wire N__43075;
    wire N__43074;
    wire N__43071;
    wire N__43070;
    wire N__43069;
    wire N__43068;
    wire N__43065;
    wire N__43062;
    wire N__43059;
    wire N__43056;
    wire N__43055;
    wire N__43054;
    wire N__43053;
    wire N__43052;
    wire N__43051;
    wire N__43050;
    wire N__43047;
    wire N__43042;
    wire N__43035;
    wire N__43030;
    wire N__43027;
    wire N__43024;
    wire N__43021;
    wire N__43020;
    wire N__43017;
    wire N__43014;
    wire N__43009;
    wire N__43008;
    wire N__43007;
    wire N__43004;
    wire N__43003;
    wire N__43000;
    wire N__42999;
    wire N__42996;
    wire N__42995;
    wire N__42994;
    wire N__42989;
    wire N__42984;
    wire N__42979;
    wire N__42976;
    wire N__42971;
    wire N__42968;
    wire N__42963;
    wire N__42956;
    wire N__42953;
    wire N__42950;
    wire N__42947;
    wire N__42944;
    wire N__42939;
    wire N__42924;
    wire N__42923;
    wire N__42920;
    wire N__42917;
    wire N__42916;
    wire N__42913;
    wire N__42908;
    wire N__42903;
    wire N__42900;
    wire N__42895;
    wire N__42890;
    wire N__42887;
    wire N__42886;
    wire N__42885;
    wire N__42882;
    wire N__42877;
    wire N__42870;
    wire N__42867;
    wire N__42862;
    wire N__42859;
    wire N__42856;
    wire N__42853;
    wire N__42848;
    wire N__42845;
    wire N__42842;
    wire N__42841;
    wire N__42838;
    wire N__42835;
    wire N__42832;
    wire N__42829;
    wire N__42824;
    wire N__42821;
    wire N__42816;
    wire N__42813;
    wire N__42810;
    wire N__42807;
    wire N__42802;
    wire N__42797;
    wire N__42788;
    wire N__42785;
    wire N__42782;
    wire N__42771;
    wire N__42768;
    wire N__42765;
    wire N__42762;
    wire N__42759;
    wire N__42756;
    wire N__42753;
    wire N__42750;
    wire N__42747;
    wire N__42744;
    wire N__42741;
    wire N__42740;
    wire N__42737;
    wire N__42736;
    wire N__42733;
    wire N__42730;
    wire N__42727;
    wire N__42720;
    wire N__42717;
    wire N__42714;
    wire N__42711;
    wire N__42708;
    wire N__42707;
    wire N__42706;
    wire N__42703;
    wire N__42700;
    wire N__42697;
    wire N__42692;
    wire N__42687;
    wire N__42684;
    wire N__42681;
    wire N__42678;
    wire N__42675;
    wire N__42672;
    wire N__42669;
    wire N__42666;
    wire N__42663;
    wire N__42660;
    wire N__42657;
    wire N__42654;
    wire N__42651;
    wire N__42648;
    wire N__42645;
    wire N__42642;
    wire N__42639;
    wire N__42636;
    wire N__42633;
    wire N__42630;
    wire N__42627;
    wire N__42624;
    wire N__42621;
    wire N__42618;
    wire N__42617;
    wire N__42616;
    wire N__42613;
    wire N__42612;
    wire N__42611;
    wire N__42610;
    wire N__42609;
    wire N__42608;
    wire N__42607;
    wire N__42606;
    wire N__42605;
    wire N__42604;
    wire N__42603;
    wire N__42600;
    wire N__42599;
    wire N__42598;
    wire N__42591;
    wire N__42580;
    wire N__42573;
    wire N__42564;
    wire N__42555;
    wire N__42552;
    wire N__42549;
    wire N__42546;
    wire N__42543;
    wire N__42540;
    wire N__42539;
    wire N__42538;
    wire N__42535;
    wire N__42532;
    wire N__42531;
    wire N__42528;
    wire N__42525;
    wire N__42522;
    wire N__42519;
    wire N__42516;
    wire N__42513;
    wire N__42510;
    wire N__42507;
    wire N__42504;
    wire N__42501;
    wire N__42496;
    wire N__42489;
    wire N__42486;
    wire N__42485;
    wire N__42484;
    wire N__42481;
    wire N__42478;
    wire N__42475;
    wire N__42472;
    wire N__42465;
    wire N__42462;
    wire N__42459;
    wire N__42456;
    wire N__42453;
    wire N__42450;
    wire N__42447;
    wire N__42446;
    wire N__42445;
    wire N__42442;
    wire N__42439;
    wire N__42436;
    wire N__42433;
    wire N__42426;
    wire N__42423;
    wire N__42420;
    wire N__42417;
    wire N__42414;
    wire N__42411;
    wire N__42408;
    wire N__42405;
    wire N__42402;
    wire N__42399;
    wire N__42396;
    wire N__42393;
    wire N__42390;
    wire N__42387;
    wire N__42384;
    wire N__42381;
    wire N__42378;
    wire N__42375;
    wire N__42372;
    wire N__42369;
    wire N__42366;
    wire N__42363;
    wire N__42362;
    wire N__42361;
    wire N__42358;
    wire N__42353;
    wire N__42348;
    wire N__42347;
    wire N__42346;
    wire N__42343;
    wire N__42338;
    wire N__42337;
    wire N__42334;
    wire N__42331;
    wire N__42328;
    wire N__42327;
    wire N__42326;
    wire N__42325;
    wire N__42324;
    wire N__42323;
    wire N__42320;
    wire N__42317;
    wire N__42314;
    wire N__42311;
    wire N__42302;
    wire N__42291;
    wire N__42290;
    wire N__42289;
    wire N__42288;
    wire N__42287;
    wire N__42286;
    wire N__42285;
    wire N__42284;
    wire N__42281;
    wire N__42278;
    wire N__42277;
    wire N__42276;
    wire N__42275;
    wire N__42274;
    wire N__42273;
    wire N__42272;
    wire N__42271;
    wire N__42270;
    wire N__42267;
    wire N__42260;
    wire N__42259;
    wire N__42258;
    wire N__42255;
    wire N__42254;
    wire N__42251;
    wire N__42250;
    wire N__42249;
    wire N__42248;
    wire N__42247;
    wire N__42238;
    wire N__42235;
    wire N__42234;
    wire N__42233;
    wire N__42232;
    wire N__42231;
    wire N__42230;
    wire N__42229;
    wire N__42228;
    wire N__42225;
    wire N__42222;
    wire N__42219;
    wire N__42214;
    wire N__42209;
    wire N__42204;
    wire N__42195;
    wire N__42188;
    wire N__42185;
    wire N__42182;
    wire N__42179;
    wire N__42176;
    wire N__42173;
    wire N__42172;
    wire N__42171;
    wire N__42168;
    wire N__42167;
    wire N__42166;
    wire N__42165;
    wire N__42164;
    wire N__42163;
    wire N__42162;
    wire N__42159;
    wire N__42158;
    wire N__42155;
    wire N__42152;
    wire N__42151;
    wire N__42148;
    wire N__42133;
    wire N__42130;
    wire N__42127;
    wire N__42122;
    wire N__42115;
    wire N__42114;
    wire N__42111;
    wire N__42106;
    wire N__42097;
    wire N__42092;
    wire N__42089;
    wire N__42084;
    wire N__42077;
    wire N__42070;
    wire N__42067;
    wire N__42048;
    wire N__42047;
    wire N__42044;
    wire N__42043;
    wire N__42042;
    wire N__42041;
    wire N__42040;
    wire N__42039;
    wire N__42038;
    wire N__42037;
    wire N__42036;
    wire N__42035;
    wire N__42034;
    wire N__42031;
    wire N__42024;
    wire N__42023;
    wire N__42022;
    wire N__42021;
    wire N__42020;
    wire N__42019;
    wire N__42018;
    wire N__42015;
    wire N__42012;
    wire N__42011;
    wire N__42010;
    wire N__42009;
    wire N__42008;
    wire N__42007;
    wire N__42004;
    wire N__42003;
    wire N__42002;
    wire N__41999;
    wire N__41998;
    wire N__41997;
    wire N__41996;
    wire N__41995;
    wire N__41994;
    wire N__41993;
    wire N__41992;
    wire N__41991;
    wire N__41988;
    wire N__41985;
    wire N__41984;
    wire N__41979;
    wire N__41978;
    wire N__41977;
    wire N__41976;
    wire N__41975;
    wire N__41972;
    wire N__41969;
    wire N__41964;
    wire N__41955;
    wire N__41948;
    wire N__41947;
    wire N__41946;
    wire N__41945;
    wire N__41944;
    wire N__41943;
    wire N__41942;
    wire N__41941;
    wire N__41940;
    wire N__41939;
    wire N__41938;
    wire N__41937;
    wire N__41936;
    wire N__41933;
    wire N__41930;
    wire N__41925;
    wire N__41924;
    wire N__41923;
    wire N__41922;
    wire N__41921;
    wire N__41916;
    wire N__41913;
    wire N__41910;
    wire N__41905;
    wire N__41900;
    wire N__41893;
    wire N__41892;
    wire N__41883;
    wire N__41880;
    wire N__41871;
    wire N__41864;
    wire N__41859;
    wire N__41848;
    wire N__41841;
    wire N__41840;
    wire N__41837;
    wire N__41830;
    wire N__41827;
    wire N__41822;
    wire N__41817;
    wire N__41816;
    wire N__41815;
    wire N__41814;
    wire N__41811;
    wire N__41808;
    wire N__41795;
    wire N__41792;
    wire N__41785;
    wire N__41778;
    wire N__41777;
    wire N__41776;
    wire N__41775;
    wire N__41774;
    wire N__41773;
    wire N__41772;
    wire N__41771;
    wire N__41770;
    wire N__41767;
    wire N__41764;
    wire N__41759;
    wire N__41752;
    wire N__41747;
    wire N__41744;
    wire N__41741;
    wire N__41736;
    wire N__41729;
    wire N__41726;
    wire N__41723;
    wire N__41710;
    wire N__41701;
    wire N__41698;
    wire N__41691;
    wire N__41688;
    wire N__41673;
    wire N__41670;
    wire N__41667;
    wire N__41664;
    wire N__41661;
    wire N__41658;
    wire N__41655;
    wire N__41652;
    wire N__41651;
    wire N__41648;
    wire N__41645;
    wire N__41642;
    wire N__41641;
    wire N__41638;
    wire N__41635;
    wire N__41632;
    wire N__41627;
    wire N__41624;
    wire N__41619;
    wire N__41618;
    wire N__41617;
    wire N__41616;
    wire N__41615;
    wire N__41614;
    wire N__41613;
    wire N__41612;
    wire N__41611;
    wire N__41610;
    wire N__41609;
    wire N__41608;
    wire N__41607;
    wire N__41606;
    wire N__41603;
    wire N__41602;
    wire N__41601;
    wire N__41600;
    wire N__41599;
    wire N__41596;
    wire N__41595;
    wire N__41590;
    wire N__41587;
    wire N__41584;
    wire N__41579;
    wire N__41576;
    wire N__41573;
    wire N__41566;
    wire N__41557;
    wire N__41552;
    wire N__41547;
    wire N__41542;
    wire N__41537;
    wire N__41534;
    wire N__41529;
    wire N__41514;
    wire N__41511;
    wire N__41508;
    wire N__41505;
    wire N__41502;
    wire N__41501;
    wire N__41500;
    wire N__41499;
    wire N__41498;
    wire N__41497;
    wire N__41496;
    wire N__41493;
    wire N__41490;
    wire N__41487;
    wire N__41484;
    wire N__41481;
    wire N__41478;
    wire N__41475;
    wire N__41474;
    wire N__41473;
    wire N__41466;
    wire N__41463;
    wire N__41458;
    wire N__41455;
    wire N__41452;
    wire N__41449;
    wire N__41448;
    wire N__41447;
    wire N__41446;
    wire N__41445;
    wire N__41444;
    wire N__41435;
    wire N__41430;
    wire N__41427;
    wire N__41424;
    wire N__41423;
    wire N__41420;
    wire N__41419;
    wire N__41416;
    wire N__41413;
    wire N__41412;
    wire N__41411;
    wire N__41406;
    wire N__41403;
    wire N__41400;
    wire N__41393;
    wire N__41390;
    wire N__41387;
    wire N__41384;
    wire N__41381;
    wire N__41380;
    wire N__41377;
    wire N__41370;
    wire N__41365;
    wire N__41360;
    wire N__41357;
    wire N__41346;
    wire N__41343;
    wire N__41340;
    wire N__41337;
    wire N__41336;
    wire N__41333;
    wire N__41332;
    wire N__41329;
    wire N__41326;
    wire N__41323;
    wire N__41320;
    wire N__41317;
    wire N__41314;
    wire N__41307;
    wire N__41304;
    wire N__41301;
    wire N__41298;
    wire N__41295;
    wire N__41292;
    wire N__41289;
    wire N__41286;
    wire N__41283;
    wire N__41280;
    wire N__41277;
    wire N__41274;
    wire N__41271;
    wire N__41268;
    wire N__41265;
    wire N__41262;
    wire N__41259;
    wire N__41256;
    wire N__41253;
    wire N__41250;
    wire N__41247;
    wire N__41246;
    wire N__41243;
    wire N__41242;
    wire N__41239;
    wire N__41236;
    wire N__41233;
    wire N__41230;
    wire N__41227;
    wire N__41222;
    wire N__41217;
    wire N__41214;
    wire N__41211;
    wire N__41208;
    wire N__41205;
    wire N__41202;
    wire N__41199;
    wire N__41196;
    wire N__41193;
    wire N__41190;
    wire N__41187;
    wire N__41184;
    wire N__41183;
    wire N__41180;
    wire N__41177;
    wire N__41172;
    wire N__41169;
    wire N__41166;
    wire N__41163;
    wire N__41160;
    wire N__41159;
    wire N__41158;
    wire N__41151;
    wire N__41148;
    wire N__41147;
    wire N__41146;
    wire N__41145;
    wire N__41142;
    wire N__41141;
    wire N__41138;
    wire N__41133;
    wire N__41132;
    wire N__41129;
    wire N__41128;
    wire N__41125;
    wire N__41124;
    wire N__41123;
    wire N__41122;
    wire N__41121;
    wire N__41118;
    wire N__41115;
    wire N__41112;
    wire N__41109;
    wire N__41106;
    wire N__41103;
    wire N__41098;
    wire N__41095;
    wire N__41094;
    wire N__41091;
    wire N__41084;
    wire N__41079;
    wire N__41074;
    wire N__41071;
    wire N__41068;
    wire N__41065;
    wire N__41064;
    wire N__41063;
    wire N__41062;
    wire N__41059;
    wire N__41054;
    wire N__41051;
    wire N__41046;
    wire N__41041;
    wire N__41038;
    wire N__41025;
    wire N__41022;
    wire N__41021;
    wire N__41018;
    wire N__41015;
    wire N__41012;
    wire N__41009;
    wire N__41006;
    wire N__41003;
    wire N__41000;
    wire N__40997;
    wire N__40992;
    wire N__40991;
    wire N__40990;
    wire N__40989;
    wire N__40988;
    wire N__40985;
    wire N__40984;
    wire N__40983;
    wire N__40982;
    wire N__40979;
    wire N__40978;
    wire N__40977;
    wire N__40974;
    wire N__40971;
    wire N__40968;
    wire N__40965;
    wire N__40962;
    wire N__40959;
    wire N__40958;
    wire N__40955;
    wire N__40952;
    wire N__40949;
    wire N__40948;
    wire N__40945;
    wire N__40936;
    wire N__40931;
    wire N__40930;
    wire N__40929;
    wire N__40928;
    wire N__40927;
    wire N__40926;
    wire N__40923;
    wire N__40918;
    wire N__40915;
    wire N__40910;
    wire N__40909;
    wire N__40904;
    wire N__40901;
    wire N__40898;
    wire N__40895;
    wire N__40892;
    wire N__40889;
    wire N__40888;
    wire N__40879;
    wire N__40876;
    wire N__40873;
    wire N__40870;
    wire N__40867;
    wire N__40864;
    wire N__40861;
    wire N__40858;
    wire N__40855;
    wire N__40852;
    wire N__40849;
    wire N__40840;
    wire N__40837;
    wire N__40824;
    wire N__40821;
    wire N__40818;
    wire N__40815;
    wire N__40812;
    wire N__40809;
    wire N__40806;
    wire N__40803;
    wire N__40800;
    wire N__40799;
    wire N__40798;
    wire N__40795;
    wire N__40792;
    wire N__40789;
    wire N__40782;
    wire N__40779;
    wire N__40776;
    wire N__40773;
    wire N__40770;
    wire N__40767;
    wire N__40764;
    wire N__40761;
    wire N__40758;
    wire N__40755;
    wire N__40754;
    wire N__40751;
    wire N__40748;
    wire N__40745;
    wire N__40742;
    wire N__40741;
    wire N__40738;
    wire N__40735;
    wire N__40732;
    wire N__40729;
    wire N__40722;
    wire N__40719;
    wire N__40716;
    wire N__40713;
    wire N__40710;
    wire N__40709;
    wire N__40708;
    wire N__40701;
    wire N__40698;
    wire N__40695;
    wire N__40692;
    wire N__40691;
    wire N__40690;
    wire N__40687;
    wire N__40684;
    wire N__40681;
    wire N__40678;
    wire N__40675;
    wire N__40672;
    wire N__40669;
    wire N__40666;
    wire N__40659;
    wire N__40656;
    wire N__40653;
    wire N__40650;
    wire N__40647;
    wire N__40644;
    wire N__40641;
    wire N__40640;
    wire N__40639;
    wire N__40636;
    wire N__40633;
    wire N__40630;
    wire N__40623;
    wire N__40622;
    wire N__40619;
    wire N__40616;
    wire N__40613;
    wire N__40610;
    wire N__40607;
    wire N__40604;
    wire N__40599;
    wire N__40596;
    wire N__40593;
    wire N__40590;
    wire N__40587;
    wire N__40584;
    wire N__40581;
    wire N__40578;
    wire N__40575;
    wire N__40574;
    wire N__40571;
    wire N__40568;
    wire N__40565;
    wire N__40562;
    wire N__40559;
    wire N__40554;
    wire N__40553;
    wire N__40552;
    wire N__40545;
    wire N__40542;
    wire N__40539;
    wire N__40536;
    wire N__40535;
    wire N__40532;
    wire N__40531;
    wire N__40528;
    wire N__40525;
    wire N__40522;
    wire N__40515;
    wire N__40512;
    wire N__40509;
    wire N__40506;
    wire N__40503;
    wire N__40500;
    wire N__40497;
    wire N__40494;
    wire N__40491;
    wire N__40490;
    wire N__40489;
    wire N__40486;
    wire N__40485;
    wire N__40482;
    wire N__40479;
    wire N__40476;
    wire N__40473;
    wire N__40472;
    wire N__40471;
    wire N__40468;
    wire N__40465;
    wire N__40460;
    wire N__40455;
    wire N__40454;
    wire N__40451;
    wire N__40448;
    wire N__40443;
    wire N__40440;
    wire N__40437;
    wire N__40432;
    wire N__40425;
    wire N__40422;
    wire N__40421;
    wire N__40418;
    wire N__40415;
    wire N__40412;
    wire N__40409;
    wire N__40408;
    wire N__40407;
    wire N__40406;
    wire N__40403;
    wire N__40400;
    wire N__40397;
    wire N__40392;
    wire N__40383;
    wire N__40380;
    wire N__40379;
    wire N__40378;
    wire N__40377;
    wire N__40374;
    wire N__40373;
    wire N__40370;
    wire N__40367;
    wire N__40364;
    wire N__40363;
    wire N__40362;
    wire N__40359;
    wire N__40352;
    wire N__40349;
    wire N__40346;
    wire N__40343;
    wire N__40340;
    wire N__40337;
    wire N__40326;
    wire N__40325;
    wire N__40322;
    wire N__40321;
    wire N__40318;
    wire N__40315;
    wire N__40312;
    wire N__40309;
    wire N__40306;
    wire N__40303;
    wire N__40302;
    wire N__40301;
    wire N__40300;
    wire N__40299;
    wire N__40296;
    wire N__40291;
    wire N__40282;
    wire N__40275;
    wire N__40272;
    wire N__40269;
    wire N__40266;
    wire N__40263;
    wire N__40260;
    wire N__40257;
    wire N__40254;
    wire N__40251;
    wire N__40248;
    wire N__40247;
    wire N__40244;
    wire N__40241;
    wire N__40238;
    wire N__40235;
    wire N__40230;
    wire N__40227;
    wire N__40224;
    wire N__40221;
    wire N__40218;
    wire N__40215;
    wire N__40212;
    wire N__40209;
    wire N__40206;
    wire N__40203;
    wire N__40200;
    wire N__40197;
    wire N__40194;
    wire N__40191;
    wire N__40188;
    wire N__40185;
    wire N__40182;
    wire N__40179;
    wire N__40176;
    wire N__40173;
    wire N__40170;
    wire N__40167;
    wire N__40164;
    wire N__40161;
    wire N__40158;
    wire N__40155;
    wire N__40152;
    wire N__40149;
    wire N__40146;
    wire N__40143;
    wire N__40140;
    wire N__40137;
    wire N__40136;
    wire N__40135;
    wire N__40134;
    wire N__40133;
    wire N__40132;
    wire N__40131;
    wire N__40130;
    wire N__40129;
    wire N__40128;
    wire N__40127;
    wire N__40126;
    wire N__40125;
    wire N__40122;
    wire N__40121;
    wire N__40118;
    wire N__40115;
    wire N__40114;
    wire N__40113;
    wire N__40110;
    wire N__40105;
    wire N__40102;
    wire N__40099;
    wire N__40096;
    wire N__40093;
    wire N__40092;
    wire N__40091;
    wire N__40088;
    wire N__40083;
    wire N__40080;
    wire N__40077;
    wire N__40072;
    wire N__40069;
    wire N__40066;
    wire N__40059;
    wire N__40056;
    wire N__40055;
    wire N__40052;
    wire N__40049;
    wire N__40044;
    wire N__40041;
    wire N__40036;
    wire N__40033;
    wire N__40022;
    wire N__40019;
    wire N__40014;
    wire N__40007;
    wire N__40002;
    wire N__39993;
    wire N__39992;
    wire N__39991;
    wire N__39988;
    wire N__39985;
    wire N__39982;
    wire N__39981;
    wire N__39976;
    wire N__39975;
    wire N__39974;
    wire N__39971;
    wire N__39968;
    wire N__39965;
    wire N__39960;
    wire N__39951;
    wire N__39948;
    wire N__39945;
    wire N__39942;
    wire N__39939;
    wire N__39936;
    wire N__39933;
    wire N__39930;
    wire N__39927;
    wire N__39924;
    wire N__39921;
    wire N__39918;
    wire N__39915;
    wire N__39912;
    wire N__39909;
    wire N__39906;
    wire N__39903;
    wire N__39900;
    wire N__39897;
    wire N__39894;
    wire N__39891;
    wire N__39888;
    wire N__39885;
    wire N__39882;
    wire N__39879;
    wire N__39876;
    wire N__39873;
    wire N__39870;
    wire N__39867;
    wire N__39864;
    wire N__39861;
    wire N__39858;
    wire N__39855;
    wire N__39852;
    wire N__39849;
    wire N__39846;
    wire N__39843;
    wire N__39840;
    wire N__39837;
    wire N__39834;
    wire N__39831;
    wire N__39828;
    wire N__39825;
    wire N__39822;
    wire N__39819;
    wire N__39816;
    wire N__39813;
    wire N__39810;
    wire N__39807;
    wire N__39804;
    wire N__39801;
    wire N__39798;
    wire N__39795;
    wire N__39792;
    wire N__39789;
    wire N__39786;
    wire N__39783;
    wire N__39780;
    wire N__39777;
    wire N__39774;
    wire N__39773;
    wire N__39770;
    wire N__39767;
    wire N__39764;
    wire N__39759;
    wire N__39756;
    wire N__39755;
    wire N__39750;
    wire N__39747;
    wire N__39746;
    wire N__39743;
    wire N__39742;
    wire N__39739;
    wire N__39738;
    wire N__39731;
    wire N__39728;
    wire N__39725;
    wire N__39722;
    wire N__39719;
    wire N__39716;
    wire N__39713;
    wire N__39710;
    wire N__39707;
    wire N__39704;
    wire N__39699;
    wire N__39698;
    wire N__39697;
    wire N__39694;
    wire N__39689;
    wire N__39684;
    wire N__39683;
    wire N__39682;
    wire N__39679;
    wire N__39676;
    wire N__39673;
    wire N__39670;
    wire N__39667;
    wire N__39660;
    wire N__39659;
    wire N__39656;
    wire N__39655;
    wire N__39652;
    wire N__39647;
    wire N__39642;
    wire N__39641;
    wire N__39638;
    wire N__39635;
    wire N__39630;
    wire N__39627;
    wire N__39624;
    wire N__39623;
    wire N__39620;
    wire N__39617;
    wire N__39612;
    wire N__39611;
    wire N__39610;
    wire N__39607;
    wire N__39604;
    wire N__39601;
    wire N__39594;
    wire N__39591;
    wire N__39588;
    wire N__39585;
    wire N__39582;
    wire N__39581;
    wire N__39578;
    wire N__39575;
    wire N__39572;
    wire N__39569;
    wire N__39566;
    wire N__39561;
    wire N__39558;
    wire N__39555;
    wire N__39552;
    wire N__39549;
    wire N__39546;
    wire N__39543;
    wire N__39540;
    wire N__39537;
    wire N__39534;
    wire N__39531;
    wire N__39530;
    wire N__39527;
    wire N__39524;
    wire N__39519;
    wire N__39518;
    wire N__39517;
    wire N__39516;
    wire N__39513;
    wire N__39512;
    wire N__39509;
    wire N__39504;
    wire N__39503;
    wire N__39502;
    wire N__39497;
    wire N__39496;
    wire N__39495;
    wire N__39494;
    wire N__39491;
    wire N__39488;
    wire N__39483;
    wire N__39480;
    wire N__39477;
    wire N__39474;
    wire N__39471;
    wire N__39468;
    wire N__39463;
    wire N__39458;
    wire N__39447;
    wire N__39444;
    wire N__39441;
    wire N__39438;
    wire N__39435;
    wire N__39432;
    wire N__39429;
    wire N__39426;
    wire N__39423;
    wire N__39420;
    wire N__39417;
    wire N__39414;
    wire N__39411;
    wire N__39408;
    wire N__39405;
    wire N__39402;
    wire N__39399;
    wire N__39396;
    wire N__39393;
    wire N__39390;
    wire N__39387;
    wire N__39386;
    wire N__39385;
    wire N__39382;
    wire N__39381;
    wire N__39378;
    wire N__39373;
    wire N__39370;
    wire N__39363;
    wire N__39360;
    wire N__39357;
    wire N__39356;
    wire N__39355;
    wire N__39354;
    wire N__39351;
    wire N__39346;
    wire N__39343;
    wire N__39336;
    wire N__39333;
    wire N__39330;
    wire N__39327;
    wire N__39324;
    wire N__39321;
    wire N__39318;
    wire N__39315;
    wire N__39312;
    wire N__39309;
    wire N__39306;
    wire N__39303;
    wire N__39300;
    wire N__39297;
    wire N__39294;
    wire N__39293;
    wire N__39290;
    wire N__39289;
    wire N__39286;
    wire N__39283;
    wire N__39280;
    wire N__39273;
    wire N__39270;
    wire N__39267;
    wire N__39264;
    wire N__39263;
    wire N__39262;
    wire N__39259;
    wire N__39256;
    wire N__39253;
    wire N__39246;
    wire N__39245;
    wire N__39244;
    wire N__39241;
    wire N__39238;
    wire N__39235;
    wire N__39228;
    wire N__39227;
    wire N__39224;
    wire N__39219;
    wire N__39216;
    wire N__39213;
    wire N__39210;
    wire N__39207;
    wire N__39204;
    wire N__39201;
    wire N__39198;
    wire N__39195;
    wire N__39192;
    wire N__39189;
    wire N__39186;
    wire N__39183;
    wire N__39180;
    wire N__39177;
    wire N__39174;
    wire N__39171;
    wire N__39168;
    wire N__39165;
    wire N__39162;
    wire N__39159;
    wire N__39156;
    wire N__39153;
    wire N__39150;
    wire N__39147;
    wire N__39144;
    wire N__39141;
    wire N__39138;
    wire N__39135;
    wire N__39132;
    wire N__39131;
    wire N__39130;
    wire N__39127;
    wire N__39126;
    wire N__39125;
    wire N__39124;
    wire N__39115;
    wire N__39112;
    wire N__39111;
    wire N__39108;
    wire N__39107;
    wire N__39104;
    wire N__39095;
    wire N__39090;
    wire N__39087;
    wire N__39084;
    wire N__39081;
    wire N__39078;
    wire N__39075;
    wire N__39072;
    wire N__39069;
    wire N__39066;
    wire N__39063;
    wire N__39060;
    wire N__39059;
    wire N__39056;
    wire N__39051;
    wire N__39048;
    wire N__39045;
    wire N__39042;
    wire N__39039;
    wire N__39036;
    wire N__39033;
    wire N__39030;
    wire N__39029;
    wire N__39026;
    wire N__39023;
    wire N__39020;
    wire N__39017;
    wire N__39014;
    wire N__39011;
    wire N__39006;
    wire N__39005;
    wire N__39002;
    wire N__39001;
    wire N__38998;
    wire N__38995;
    wire N__38992;
    wire N__38985;
    wire N__38984;
    wire N__38983;
    wire N__38980;
    wire N__38977;
    wire N__38976;
    wire N__38975;
    wire N__38974;
    wire N__38973;
    wire N__38972;
    wire N__38971;
    wire N__38968;
    wire N__38965;
    wire N__38958;
    wire N__38953;
    wire N__38950;
    wire N__38949;
    wire N__38948;
    wire N__38947;
    wire N__38946;
    wire N__38945;
    wire N__38942;
    wire N__38939;
    wire N__38932;
    wire N__38929;
    wire N__38926;
    wire N__38925;
    wire N__38922;
    wire N__38919;
    wire N__38918;
    wire N__38917;
    wire N__38916;
    wire N__38913;
    wire N__38910;
    wire N__38907;
    wire N__38898;
    wire N__38895;
    wire N__38892;
    wire N__38889;
    wire N__38886;
    wire N__38879;
    wire N__38876;
    wire N__38869;
    wire N__38864;
    wire N__38861;
    wire N__38860;
    wire N__38859;
    wire N__38858;
    wire N__38857;
    wire N__38852;
    wire N__38849;
    wire N__38844;
    wire N__38841;
    wire N__38834;
    wire N__38823;
    wire N__38820;
    wire N__38817;
    wire N__38814;
    wire N__38811;
    wire N__38808;
    wire N__38805;
    wire N__38802;
    wire N__38801;
    wire N__38800;
    wire N__38797;
    wire N__38792;
    wire N__38787;
    wire N__38784;
    wire N__38781;
    wire N__38778;
    wire N__38775;
    wire N__38772;
    wire N__38769;
    wire N__38766;
    wire N__38763;
    wire N__38760;
    wire N__38757;
    wire N__38754;
    wire N__38751;
    wire N__38748;
    wire N__38745;
    wire N__38742;
    wire N__38739;
    wire N__38736;
    wire N__38733;
    wire N__38730;
    wire N__38727;
    wire N__38724;
    wire N__38721;
    wire N__38718;
    wire N__38715;
    wire N__38712;
    wire N__38709;
    wire N__38706;
    wire N__38703;
    wire N__38700;
    wire N__38697;
    wire N__38694;
    wire N__38691;
    wire N__38688;
    wire N__38685;
    wire N__38682;
    wire N__38679;
    wire N__38676;
    wire N__38673;
    wire N__38670;
    wire N__38667;
    wire N__38664;
    wire N__38661;
    wire N__38658;
    wire N__38655;
    wire N__38652;
    wire N__38649;
    wire N__38646;
    wire N__38643;
    wire N__38640;
    wire N__38637;
    wire N__38634;
    wire N__38631;
    wire N__38628;
    wire N__38625;
    wire N__38622;
    wire N__38619;
    wire N__38616;
    wire N__38613;
    wire N__38610;
    wire N__38607;
    wire N__38604;
    wire N__38601;
    wire N__38598;
    wire N__38595;
    wire N__38592;
    wire N__38589;
    wire N__38586;
    wire N__38583;
    wire N__38580;
    wire N__38577;
    wire N__38574;
    wire N__38571;
    wire N__38568;
    wire N__38565;
    wire N__38562;
    wire N__38559;
    wire N__38556;
    wire N__38553;
    wire N__38550;
    wire N__38547;
    wire N__38544;
    wire N__38541;
    wire N__38538;
    wire N__38535;
    wire N__38532;
    wire N__38529;
    wire N__38526;
    wire N__38523;
    wire N__38520;
    wire N__38517;
    wire N__38514;
    wire N__38511;
    wire N__38508;
    wire N__38505;
    wire N__38502;
    wire N__38499;
    wire N__38496;
    wire N__38493;
    wire N__38490;
    wire N__38487;
    wire N__38484;
    wire N__38481;
    wire N__38478;
    wire N__38475;
    wire N__38472;
    wire N__38469;
    wire N__38466;
    wire N__38463;
    wire N__38460;
    wire N__38457;
    wire N__38454;
    wire N__38451;
    wire N__38448;
    wire N__38445;
    wire N__38442;
    wire N__38439;
    wire N__38436;
    wire N__38433;
    wire N__38430;
    wire N__38427;
    wire N__38424;
    wire N__38421;
    wire N__38418;
    wire N__38415;
    wire N__38412;
    wire N__38409;
    wire N__38406;
    wire N__38405;
    wire N__38402;
    wire N__38401;
    wire N__38398;
    wire N__38395;
    wire N__38392;
    wire N__38387;
    wire N__38384;
    wire N__38379;
    wire N__38376;
    wire N__38373;
    wire N__38372;
    wire N__38369;
    wire N__38366;
    wire N__38363;
    wire N__38358;
    wire N__38355;
    wire N__38352;
    wire N__38349;
    wire N__38346;
    wire N__38343;
    wire N__38340;
    wire N__38337;
    wire N__38334;
    wire N__38331;
    wire N__38328;
    wire N__38325;
    wire N__38322;
    wire N__38319;
    wire N__38316;
    wire N__38313;
    wire N__38310;
    wire N__38307;
    wire N__38304;
    wire N__38301;
    wire N__38298;
    wire N__38295;
    wire N__38292;
    wire N__38289;
    wire N__38286;
    wire N__38283;
    wire N__38280;
    wire N__38277;
    wire N__38274;
    wire N__38271;
    wire N__38268;
    wire N__38265;
    wire N__38262;
    wire N__38259;
    wire N__38256;
    wire N__38253;
    wire N__38250;
    wire N__38247;
    wire N__38244;
    wire N__38241;
    wire N__38238;
    wire N__38235;
    wire N__38232;
    wire N__38229;
    wire N__38226;
    wire N__38223;
    wire N__38220;
    wire N__38217;
    wire N__38214;
    wire N__38211;
    wire N__38208;
    wire N__38205;
    wire N__38202;
    wire N__38199;
    wire N__38196;
    wire N__38193;
    wire N__38190;
    wire N__38187;
    wire N__38184;
    wire N__38181;
    wire N__38178;
    wire N__38175;
    wire N__38172;
    wire N__38169;
    wire N__38166;
    wire N__38163;
    wire N__38160;
    wire N__38157;
    wire N__38154;
    wire N__38151;
    wire N__38148;
    wire N__38145;
    wire N__38144;
    wire N__38141;
    wire N__38138;
    wire N__38135;
    wire N__38132;
    wire N__38129;
    wire N__38124;
    wire N__38121;
    wire N__38118;
    wire N__38115;
    wire N__38112;
    wire N__38109;
    wire N__38106;
    wire N__38103;
    wire N__38100;
    wire N__38097;
    wire N__38096;
    wire N__38093;
    wire N__38090;
    wire N__38087;
    wire N__38084;
    wire N__38081;
    wire N__38076;
    wire N__38073;
    wire N__38070;
    wire N__38067;
    wire N__38064;
    wire N__38061;
    wire N__38058;
    wire N__38055;
    wire N__38052;
    wire N__38049;
    wire N__38046;
    wire N__38045;
    wire N__38042;
    wire N__38039;
    wire N__38036;
    wire N__38031;
    wire N__38028;
    wire N__38025;
    wire N__38022;
    wire N__38019;
    wire N__38016;
    wire N__38013;
    wire N__38010;
    wire N__38007;
    wire N__38004;
    wire N__38001;
    wire N__38000;
    wire N__37997;
    wire N__37994;
    wire N__37991;
    wire N__37986;
    wire N__37983;
    wire N__37980;
    wire N__37977;
    wire N__37974;
    wire N__37973;
    wire N__37970;
    wire N__37967;
    wire N__37964;
    wire N__37961;
    wire N__37958;
    wire N__37953;
    wire N__37950;
    wire N__37947;
    wire N__37944;
    wire N__37941;
    wire N__37938;
    wire N__37935;
    wire N__37932;
    wire N__37929;
    wire N__37928;
    wire N__37925;
    wire N__37922;
    wire N__37917;
    wire N__37914;
    wire N__37911;
    wire N__37908;
    wire N__37905;
    wire N__37902;
    wire N__37899;
    wire N__37898;
    wire N__37895;
    wire N__37892;
    wire N__37887;
    wire N__37884;
    wire N__37881;
    wire N__37878;
    wire N__37875;
    wire N__37872;
    wire N__37869;
    wire N__37866;
    wire N__37865;
    wire N__37862;
    wire N__37859;
    wire N__37856;
    wire N__37851;
    wire N__37848;
    wire N__37845;
    wire N__37842;
    wire N__37839;
    wire N__37836;
    wire N__37833;
    wire N__37832;
    wire N__37829;
    wire N__37826;
    wire N__37823;
    wire N__37820;
    wire N__37817;
    wire N__37814;
    wire N__37809;
    wire N__37806;
    wire N__37803;
    wire N__37800;
    wire N__37797;
    wire N__37794;
    wire N__37791;
    wire N__37788;
    wire N__37787;
    wire N__37784;
    wire N__37781;
    wire N__37778;
    wire N__37773;
    wire N__37770;
    wire N__37767;
    wire N__37764;
    wire N__37763;
    wire N__37762;
    wire N__37757;
    wire N__37754;
    wire N__37751;
    wire N__37746;
    wire N__37743;
    wire N__37740;
    wire N__37739;
    wire N__37738;
    wire N__37735;
    wire N__37730;
    wire N__37725;
    wire N__37722;
    wire N__37719;
    wire N__37718;
    wire N__37717;
    wire N__37714;
    wire N__37713;
    wire N__37712;
    wire N__37705;
    wire N__37704;
    wire N__37703;
    wire N__37700;
    wire N__37697;
    wire N__37694;
    wire N__37691;
    wire N__37688;
    wire N__37687;
    wire N__37686;
    wire N__37683;
    wire N__37680;
    wire N__37675;
    wire N__37670;
    wire N__37667;
    wire N__37662;
    wire N__37653;
    wire N__37652;
    wire N__37651;
    wire N__37650;
    wire N__37647;
    wire N__37642;
    wire N__37639;
    wire N__37632;
    wire N__37631;
    wire N__37630;
    wire N__37627;
    wire N__37624;
    wire N__37621;
    wire N__37618;
    wire N__37615;
    wire N__37612;
    wire N__37609;
    wire N__37604;
    wire N__37601;
    wire N__37596;
    wire N__37593;
    wire N__37592;
    wire N__37591;
    wire N__37590;
    wire N__37587;
    wire N__37584;
    wire N__37583;
    wire N__37582;
    wire N__37581;
    wire N__37578;
    wire N__37575;
    wire N__37574;
    wire N__37569;
    wire N__37568;
    wire N__37565;
    wire N__37562;
    wire N__37559;
    wire N__37554;
    wire N__37553;
    wire N__37552;
    wire N__37551;
    wire N__37550;
    wire N__37549;
    wire N__37548;
    wire N__37545;
    wire N__37542;
    wire N__37539;
    wire N__37530;
    wire N__37525;
    wire N__37518;
    wire N__37515;
    wire N__37512;
    wire N__37497;
    wire N__37494;
    wire N__37491;
    wire N__37488;
    wire N__37487;
    wire N__37486;
    wire N__37483;
    wire N__37480;
    wire N__37477;
    wire N__37470;
    wire N__37469;
    wire N__37468;
    wire N__37461;
    wire N__37458;
    wire N__37455;
    wire N__37454;
    wire N__37451;
    wire N__37448;
    wire N__37443;
    wire N__37440;
    wire N__37437;
    wire N__37434;
    wire N__37431;
    wire N__37428;
    wire N__37427;
    wire N__37426;
    wire N__37419;
    wire N__37416;
    wire N__37413;
    wire N__37412;
    wire N__37409;
    wire N__37406;
    wire N__37401;
    wire N__37398;
    wire N__37395;
    wire N__37392;
    wire N__37389;
    wire N__37386;
    wire N__37385;
    wire N__37384;
    wire N__37381;
    wire N__37376;
    wire N__37371;
    wire N__37370;
    wire N__37367;
    wire N__37364;
    wire N__37359;
    wire N__37358;
    wire N__37355;
    wire N__37352;
    wire N__37347;
    wire N__37344;
    wire N__37343;
    wire N__37340;
    wire N__37337;
    wire N__37332;
    wire N__37331;
    wire N__37328;
    wire N__37325;
    wire N__37320;
    wire N__37319;
    wire N__37318;
    wire N__37317;
    wire N__37314;
    wire N__37311;
    wire N__37308;
    wire N__37305;
    wire N__37302;
    wire N__37299;
    wire N__37294;
    wire N__37291;
    wire N__37288;
    wire N__37285;
    wire N__37282;
    wire N__37275;
    wire N__37272;
    wire N__37269;
    wire N__37266;
    wire N__37263;
    wire N__37262;
    wire N__37261;
    wire N__37260;
    wire N__37259;
    wire N__37258;
    wire N__37257;
    wire N__37256;
    wire N__37255;
    wire N__37254;
    wire N__37251;
    wire N__37250;
    wire N__37247;
    wire N__37244;
    wire N__37243;
    wire N__37242;
    wire N__37241;
    wire N__37240;
    wire N__37237;
    wire N__37234;
    wire N__37233;
    wire N__37232;
    wire N__37231;
    wire N__37228;
    wire N__37227;
    wire N__37226;
    wire N__37225;
    wire N__37224;
    wire N__37221;
    wire N__37218;
    wire N__37215;
    wire N__37214;
    wire N__37207;
    wire N__37204;
    wire N__37203;
    wire N__37200;
    wire N__37197;
    wire N__37194;
    wire N__37193;
    wire N__37192;
    wire N__37191;
    wire N__37188;
    wire N__37181;
    wire N__37172;
    wire N__37169;
    wire N__37166;
    wire N__37165;
    wire N__37158;
    wire N__37151;
    wire N__37150;
    wire N__37149;
    wire N__37148;
    wire N__37147;
    wire N__37142;
    wire N__37139;
    wire N__37136;
    wire N__37129;
    wire N__37122;
    wire N__37117;
    wire N__37110;
    wire N__37105;
    wire N__37104;
    wire N__37103;
    wire N__37102;
    wire N__37099;
    wire N__37096;
    wire N__37093;
    wire N__37092;
    wire N__37091;
    wire N__37090;
    wire N__37089;
    wire N__37086;
    wire N__37083;
    wire N__37080;
    wire N__37071;
    wire N__37068;
    wire N__37065;
    wire N__37054;
    wire N__37047;
    wire N__37040;
    wire N__37037;
    wire N__37032;
    wire N__37029;
    wire N__37026;
    wire N__37021;
    wire N__37012;
    wire N__37009;
    wire N__37006;
    wire N__37003;
    wire N__36996;
    wire N__36993;
    wire N__36992;
    wire N__36989;
    wire N__36988;
    wire N__36985;
    wire N__36982;
    wire N__36979;
    wire N__36976;
    wire N__36971;
    wire N__36966;
    wire N__36965;
    wire N__36964;
    wire N__36963;
    wire N__36960;
    wire N__36957;
    wire N__36952;
    wire N__36945;
    wire N__36942;
    wire N__36941;
    wire N__36940;
    wire N__36939;
    wire N__36936;
    wire N__36933;
    wire N__36928;
    wire N__36921;
    wire N__36918;
    wire N__36915;
    wire N__36912;
    wire N__36909;
    wire N__36906;
    wire N__36903;
    wire N__36902;
    wire N__36901;
    wire N__36894;
    wire N__36891;
    wire N__36888;
    wire N__36887;
    wire N__36884;
    wire N__36881;
    wire N__36880;
    wire N__36877;
    wire N__36874;
    wire N__36873;
    wire N__36872;
    wire N__36871;
    wire N__36868;
    wire N__36867;
    wire N__36866;
    wire N__36865;
    wire N__36864;
    wire N__36861;
    wire N__36858;
    wire N__36857;
    wire N__36856;
    wire N__36855;
    wire N__36852;
    wire N__36849;
    wire N__36846;
    wire N__36843;
    wire N__36840;
    wire N__36839;
    wire N__36838;
    wire N__36835;
    wire N__36832;
    wire N__36829;
    wire N__36826;
    wire N__36823;
    wire N__36820;
    wire N__36819;
    wire N__36816;
    wire N__36813;
    wire N__36810;
    wire N__36807;
    wire N__36802;
    wire N__36799;
    wire N__36792;
    wire N__36781;
    wire N__36778;
    wire N__36769;
    wire N__36766;
    wire N__36759;
    wire N__36750;
    wire N__36747;
    wire N__36744;
    wire N__36741;
    wire N__36738;
    wire N__36735;
    wire N__36732;
    wire N__36729;
    wire N__36726;
    wire N__36723;
    wire N__36720;
    wire N__36717;
    wire N__36714;
    wire N__36711;
    wire N__36710;
    wire N__36707;
    wire N__36704;
    wire N__36699;
    wire N__36696;
    wire N__36693;
    wire N__36692;
    wire N__36691;
    wire N__36688;
    wire N__36687;
    wire N__36686;
    wire N__36683;
    wire N__36680;
    wire N__36679;
    wire N__36678;
    wire N__36677;
    wire N__36672;
    wire N__36671;
    wire N__36668;
    wire N__36663;
    wire N__36660;
    wire N__36655;
    wire N__36652;
    wire N__36649;
    wire N__36646;
    wire N__36641;
    wire N__36638;
    wire N__36633;
    wire N__36626;
    wire N__36623;
    wire N__36618;
    wire N__36617;
    wire N__36616;
    wire N__36615;
    wire N__36612;
    wire N__36609;
    wire N__36608;
    wire N__36607;
    wire N__36606;
    wire N__36605;
    wire N__36604;
    wire N__36601;
    wire N__36598;
    wire N__36595;
    wire N__36592;
    wire N__36589;
    wire N__36586;
    wire N__36583;
    wire N__36580;
    wire N__36577;
    wire N__36572;
    wire N__36567;
    wire N__36564;
    wire N__36549;
    wire N__36546;
    wire N__36545;
    wire N__36544;
    wire N__36541;
    wire N__36538;
    wire N__36537;
    wire N__36536;
    wire N__36535;
    wire N__36532;
    wire N__36531;
    wire N__36526;
    wire N__36525;
    wire N__36522;
    wire N__36519;
    wire N__36516;
    wire N__36513;
    wire N__36510;
    wire N__36507;
    wire N__36504;
    wire N__36489;
    wire N__36488;
    wire N__36485;
    wire N__36484;
    wire N__36483;
    wire N__36480;
    wire N__36477;
    wire N__36476;
    wire N__36475;
    wire N__36472;
    wire N__36469;
    wire N__36464;
    wire N__36459;
    wire N__36450;
    wire N__36447;
    wire N__36444;
    wire N__36441;
    wire N__36438;
    wire N__36435;
    wire N__36432;
    wire N__36429;
    wire N__36426;
    wire N__36423;
    wire N__36420;
    wire N__36417;
    wire N__36416;
    wire N__36413;
    wire N__36410;
    wire N__36407;
    wire N__36404;
    wire N__36401;
    wire N__36396;
    wire N__36393;
    wire N__36392;
    wire N__36391;
    wire N__36388;
    wire N__36385;
    wire N__36382;
    wire N__36379;
    wire N__36372;
    wire N__36371;
    wire N__36370;
    wire N__36369;
    wire N__36366;
    wire N__36361;
    wire N__36358;
    wire N__36351;
    wire N__36348;
    wire N__36345;
    wire N__36342;
    wire N__36341;
    wire N__36340;
    wire N__36337;
    wire N__36334;
    wire N__36331;
    wire N__36324;
    wire N__36321;
    wire N__36320;
    wire N__36319;
    wire N__36316;
    wire N__36313;
    wire N__36310;
    wire N__36303;
    wire N__36300;
    wire N__36297;
    wire N__36294;
    wire N__36291;
    wire N__36290;
    wire N__36287;
    wire N__36284;
    wire N__36279;
    wire N__36276;
    wire N__36273;
    wire N__36270;
    wire N__36267;
    wire N__36266;
    wire N__36263;
    wire N__36262;
    wire N__36259;
    wire N__36256;
    wire N__36253;
    wire N__36250;
    wire N__36245;
    wire N__36244;
    wire N__36241;
    wire N__36238;
    wire N__36235;
    wire N__36228;
    wire N__36227;
    wire N__36224;
    wire N__36221;
    wire N__36216;
    wire N__36213;
    wire N__36212;
    wire N__36209;
    wire N__36206;
    wire N__36205;
    wire N__36202;
    wire N__36199;
    wire N__36196;
    wire N__36191;
    wire N__36186;
    wire N__36185;
    wire N__36182;
    wire N__36179;
    wire N__36176;
    wire N__36173;
    wire N__36170;
    wire N__36167;
    wire N__36162;
    wire N__36159;
    wire N__36156;
    wire N__36153;
    wire N__36150;
    wire N__36149;
    wire N__36148;
    wire N__36145;
    wire N__36142;
    wire N__36139;
    wire N__36136;
    wire N__36129;
    wire N__36126;
    wire N__36123;
    wire N__36120;
    wire N__36117;
    wire N__36114;
    wire N__36111;
    wire N__36108;
    wire N__36105;
    wire N__36102;
    wire N__36099;
    wire N__36096;
    wire N__36093;
    wire N__36090;
    wire N__36087;
    wire N__36084;
    wire N__36081;
    wire N__36078;
    wire N__36075;
    wire N__36072;
    wire N__36069;
    wire N__36066;
    wire N__36063;
    wire N__36060;
    wire N__36057;
    wire N__36054;
    wire N__36051;
    wire N__36048;
    wire N__36047;
    wire N__36044;
    wire N__36041;
    wire N__36038;
    wire N__36035;
    wire N__36032;
    wire N__36027;
    wire N__36024;
    wire N__36021;
    wire N__36018;
    wire N__36015;
    wire N__36014;
    wire N__36011;
    wire N__36008;
    wire N__36005;
    wire N__36000;
    wire N__35997;
    wire N__35994;
    wire N__35991;
    wire N__35988;
    wire N__35985;
    wire N__35984;
    wire N__35981;
    wire N__35978;
    wire N__35975;
    wire N__35972;
    wire N__35967;
    wire N__35964;
    wire N__35961;
    wire N__35958;
    wire N__35955;
    wire N__35952;
    wire N__35949;
    wire N__35946;
    wire N__35945;
    wire N__35942;
    wire N__35939;
    wire N__35936;
    wire N__35933;
    wire N__35930;
    wire N__35927;
    wire N__35922;
    wire N__35919;
    wire N__35916;
    wire N__35913;
    wire N__35910;
    wire N__35907;
    wire N__35906;
    wire N__35903;
    wire N__35900;
    wire N__35897;
    wire N__35894;
    wire N__35891;
    wire N__35888;
    wire N__35883;
    wire N__35880;
    wire N__35877;
    wire N__35874;
    wire N__35871;
    wire N__35868;
    wire N__35865;
    wire N__35862;
    wire N__35859;
    wire N__35858;
    wire N__35855;
    wire N__35852;
    wire N__35849;
    wire N__35848;
    wire N__35845;
    wire N__35842;
    wire N__35839;
    wire N__35832;
    wire N__35829;
    wire N__35826;
    wire N__35823;
    wire N__35820;
    wire N__35819;
    wire N__35818;
    wire N__35815;
    wire N__35814;
    wire N__35811;
    wire N__35808;
    wire N__35805;
    wire N__35802;
    wire N__35801;
    wire N__35800;
    wire N__35791;
    wire N__35788;
    wire N__35785;
    wire N__35784;
    wire N__35783;
    wire N__35782;
    wire N__35781;
    wire N__35780;
    wire N__35779;
    wire N__35772;
    wire N__35769;
    wire N__35766;
    wire N__35761;
    wire N__35756;
    wire N__35745;
    wire N__35744;
    wire N__35741;
    wire N__35738;
    wire N__35735;
    wire N__35734;
    wire N__35733;
    wire N__35732;
    wire N__35731;
    wire N__35730;
    wire N__35729;
    wire N__35728;
    wire N__35723;
    wire N__35720;
    wire N__35717;
    wire N__35714;
    wire N__35711;
    wire N__35708;
    wire N__35703;
    wire N__35698;
    wire N__35697;
    wire N__35690;
    wire N__35685;
    wire N__35684;
    wire N__35683;
    wire N__35680;
    wire N__35677;
    wire N__35672;
    wire N__35667;
    wire N__35658;
    wire N__35655;
    wire N__35652;
    wire N__35649;
    wire N__35646;
    wire N__35645;
    wire N__35642;
    wire N__35639;
    wire N__35636;
    wire N__35633;
    wire N__35630;
    wire N__35625;
    wire N__35624;
    wire N__35621;
    wire N__35616;
    wire N__35613;
    wire N__35610;
    wire N__35607;
    wire N__35604;
    wire N__35601;
    wire N__35600;
    wire N__35597;
    wire N__35594;
    wire N__35591;
    wire N__35586;
    wire N__35583;
    wire N__35582;
    wire N__35579;
    wire N__35576;
    wire N__35573;
    wire N__35568;
    wire N__35565;
    wire N__35562;
    wire N__35559;
    wire N__35556;
    wire N__35553;
    wire N__35550;
    wire N__35549;
    wire N__35548;
    wire N__35547;
    wire N__35544;
    wire N__35537;
    wire N__35532;
    wire N__35531;
    wire N__35528;
    wire N__35527;
    wire N__35524;
    wire N__35523;
    wire N__35520;
    wire N__35517;
    wire N__35512;
    wire N__35509;
    wire N__35506;
    wire N__35503;
    wire N__35500;
    wire N__35497;
    wire N__35490;
    wire N__35487;
    wire N__35484;
    wire N__35481;
    wire N__35478;
    wire N__35477;
    wire N__35474;
    wire N__35473;
    wire N__35470;
    wire N__35467;
    wire N__35464;
    wire N__35461;
    wire N__35456;
    wire N__35451;
    wire N__35450;
    wire N__35447;
    wire N__35446;
    wire N__35443;
    wire N__35440;
    wire N__35435;
    wire N__35430;
    wire N__35429;
    wire N__35426;
    wire N__35423;
    wire N__35420;
    wire N__35417;
    wire N__35412;
    wire N__35409;
    wire N__35408;
    wire N__35405;
    wire N__35402;
    wire N__35399;
    wire N__35396;
    wire N__35393;
    wire N__35388;
    wire N__35385;
    wire N__35382;
    wire N__35379;
    wire N__35378;
    wire N__35375;
    wire N__35374;
    wire N__35371;
    wire N__35368;
    wire N__35365;
    wire N__35360;
    wire N__35357;
    wire N__35354;
    wire N__35349;
    wire N__35346;
    wire N__35343;
    wire N__35340;
    wire N__35339;
    wire N__35338;
    wire N__35335;
    wire N__35330;
    wire N__35327;
    wire N__35322;
    wire N__35319;
    wire N__35316;
    wire N__35313;
    wire N__35310;
    wire N__35309;
    wire N__35308;
    wire N__35307;
    wire N__35302;
    wire N__35299;
    wire N__35296;
    wire N__35289;
    wire N__35288;
    wire N__35287;
    wire N__35286;
    wire N__35285;
    wire N__35282;
    wire N__35279;
    wire N__35276;
    wire N__35273;
    wire N__35270;
    wire N__35269;
    wire N__35268;
    wire N__35267;
    wire N__35256;
    wire N__35251;
    wire N__35250;
    wire N__35249;
    wire N__35248;
    wire N__35245;
    wire N__35240;
    wire N__35233;
    wire N__35226;
    wire N__35223;
    wire N__35222;
    wire N__35219;
    wire N__35218;
    wire N__35215;
    wire N__35212;
    wire N__35209;
    wire N__35206;
    wire N__35203;
    wire N__35196;
    wire N__35193;
    wire N__35192;
    wire N__35189;
    wire N__35186;
    wire N__35181;
    wire N__35180;
    wire N__35177;
    wire N__35174;
    wire N__35169;
    wire N__35168;
    wire N__35165;
    wire N__35160;
    wire N__35157;
    wire N__35156;
    wire N__35153;
    wire N__35150;
    wire N__35145;
    wire N__35142;
    wire N__35139;
    wire N__35136;
    wire N__35133;
    wire N__35130;
    wire N__35129;
    wire N__35128;
    wire N__35125;
    wire N__35122;
    wire N__35119;
    wire N__35112;
    wire N__35109;
    wire N__35106;
    wire N__35105;
    wire N__35102;
    wire N__35099;
    wire N__35094;
    wire N__35091;
    wire N__35088;
    wire N__35087;
    wire N__35084;
    wire N__35081;
    wire N__35078;
    wire N__35073;
    wire N__35070;
    wire N__35067;
    wire N__35066;
    wire N__35063;
    wire N__35060;
    wire N__35057;
    wire N__35052;
    wire N__35049;
    wire N__35046;
    wire N__35043;
    wire N__35042;
    wire N__35037;
    wire N__35034;
    wire N__35033;
    wire N__35030;
    wire N__35027;
    wire N__35022;
    wire N__35019;
    wire N__35018;
    wire N__35015;
    wire N__35012;
    wire N__35007;
    wire N__35004;
    wire N__35003;
    wire N__35000;
    wire N__34997;
    wire N__34992;
    wire N__34989;
    wire N__34988;
    wire N__34985;
    wire N__34982;
    wire N__34977;
    wire N__34974;
    wire N__34971;
    wire N__34970;
    wire N__34967;
    wire N__34964;
    wire N__34961;
    wire N__34956;
    wire N__34953;
    wire N__34950;
    wire N__34947;
    wire N__34946;
    wire N__34943;
    wire N__34940;
    wire N__34935;
    wire N__34932;
    wire N__34929;
    wire N__34928;
    wire N__34925;
    wire N__34922;
    wire N__34921;
    wire N__34918;
    wire N__34915;
    wire N__34912;
    wire N__34909;
    wire N__34902;
    wire N__34899;
    wire N__34896;
    wire N__34893;
    wire N__34892;
    wire N__34889;
    wire N__34886;
    wire N__34881;
    wire N__34878;
    wire N__34875;
    wire N__34872;
    wire N__34869;
    wire N__34866;
    wire N__34863;
    wire N__34860;
    wire N__34857;
    wire N__34854;
    wire N__34853;
    wire N__34850;
    wire N__34849;
    wire N__34846;
    wire N__34843;
    wire N__34840;
    wire N__34833;
    wire N__34832;
    wire N__34831;
    wire N__34828;
    wire N__34825;
    wire N__34822;
    wire N__34819;
    wire N__34818;
    wire N__34815;
    wire N__34812;
    wire N__34809;
    wire N__34806;
    wire N__34803;
    wire N__34798;
    wire N__34791;
    wire N__34790;
    wire N__34787;
    wire N__34784;
    wire N__34779;
    wire N__34776;
    wire N__34773;
    wire N__34770;
    wire N__34769;
    wire N__34766;
    wire N__34763;
    wire N__34758;
    wire N__34755;
    wire N__34754;
    wire N__34751;
    wire N__34748;
    wire N__34745;
    wire N__34740;
    wire N__34737;
    wire N__34736;
    wire N__34735;
    wire N__34732;
    wire N__34727;
    wire N__34722;
    wire N__34719;
    wire N__34716;
    wire N__34713;
    wire N__34712;
    wire N__34711;
    wire N__34704;
    wire N__34701;
    wire N__34698;
    wire N__34695;
    wire N__34692;
    wire N__34689;
    wire N__34686;
    wire N__34683;
    wire N__34680;
    wire N__34679;
    wire N__34676;
    wire N__34675;
    wire N__34672;
    wire N__34671;
    wire N__34668;
    wire N__34665;
    wire N__34660;
    wire N__34653;
    wire N__34650;
    wire N__34647;
    wire N__34644;
    wire N__34641;
    wire N__34638;
    wire N__34635;
    wire N__34632;
    wire N__34631;
    wire N__34630;
    wire N__34627;
    wire N__34624;
    wire N__34619;
    wire N__34614;
    wire N__34611;
    wire N__34608;
    wire N__34605;
    wire N__34602;
    wire N__34601;
    wire N__34600;
    wire N__34597;
    wire N__34594;
    wire N__34591;
    wire N__34584;
    wire N__34581;
    wire N__34578;
    wire N__34577;
    wire N__34574;
    wire N__34571;
    wire N__34570;
    wire N__34567;
    wire N__34564;
    wire N__34561;
    wire N__34558;
    wire N__34555;
    wire N__34548;
    wire N__34545;
    wire N__34542;
    wire N__34539;
    wire N__34536;
    wire N__34533;
    wire N__34530;
    wire N__34527;
    wire N__34524;
    wire N__34521;
    wire N__34520;
    wire N__34517;
    wire N__34514;
    wire N__34509;
    wire N__34506;
    wire N__34503;
    wire N__34500;
    wire N__34499;
    wire N__34496;
    wire N__34493;
    wire N__34490;
    wire N__34487;
    wire N__34484;
    wire N__34481;
    wire N__34476;
    wire N__34473;
    wire N__34470;
    wire N__34467;
    wire N__34464;
    wire N__34461;
    wire N__34460;
    wire N__34457;
    wire N__34454;
    wire N__34449;
    wire N__34446;
    wire N__34443;
    wire N__34440;
    wire N__34437;
    wire N__34434;
    wire N__34431;
    wire N__34428;
    wire N__34425;
    wire N__34424;
    wire N__34423;
    wire N__34420;
    wire N__34417;
    wire N__34412;
    wire N__34407;
    wire N__34406;
    wire N__34405;
    wire N__34402;
    wire N__34399;
    wire N__34394;
    wire N__34389;
    wire N__34386;
    wire N__34385;
    wire N__34384;
    wire N__34381;
    wire N__34376;
    wire N__34371;
    wire N__34368;
    wire N__34367;
    wire N__34366;
    wire N__34359;
    wire N__34356;
    wire N__34355;
    wire N__34352;
    wire N__34349;
    wire N__34346;
    wire N__34343;
    wire N__34340;
    wire N__34335;
    wire N__34334;
    wire N__34333;
    wire N__34330;
    wire N__34323;
    wire N__34320;
    wire N__34317;
    wire N__34314;
    wire N__34311;
    wire N__34308;
    wire N__34307;
    wire N__34304;
    wire N__34301;
    wire N__34298;
    wire N__34295;
    wire N__34292;
    wire N__34289;
    wire N__34286;
    wire N__34283;
    wire N__34278;
    wire N__34277;
    wire N__34276;
    wire N__34271;
    wire N__34268;
    wire N__34263;
    wire N__34260;
    wire N__34257;
    wire N__34254;
    wire N__34251;
    wire N__34250;
    wire N__34247;
    wire N__34242;
    wire N__34241;
    wire N__34238;
    wire N__34235;
    wire N__34232;
    wire N__34227;
    wire N__34224;
    wire N__34223;
    wire N__34220;
    wire N__34217;
    wire N__34214;
    wire N__34211;
    wire N__34208;
    wire N__34205;
    wire N__34200;
    wire N__34197;
    wire N__34194;
    wire N__34191;
    wire N__34188;
    wire N__34185;
    wire N__34184;
    wire N__34183;
    wire N__34180;
    wire N__34175;
    wire N__34172;
    wire N__34167;
    wire N__34166;
    wire N__34163;
    wire N__34160;
    wire N__34157;
    wire N__34154;
    wire N__34149;
    wire N__34146;
    wire N__34143;
    wire N__34140;
    wire N__34139;
    wire N__34136;
    wire N__34133;
    wire N__34128;
    wire N__34125;
    wire N__34122;
    wire N__34119;
    wire N__34116;
    wire N__34113;
    wire N__34110;
    wire N__34107;
    wire N__34104;
    wire N__34101;
    wire N__34100;
    wire N__34095;
    wire N__34092;
    wire N__34089;
    wire N__34086;
    wire N__34083;
    wire N__34080;
    wire N__34077;
    wire N__34074;
    wire N__34071;
    wire N__34068;
    wire N__34065;
    wire N__34064;
    wire N__34061;
    wire N__34060;
    wire N__34057;
    wire N__34054;
    wire N__34049;
    wire N__34044;
    wire N__34041;
    wire N__34040;
    wire N__34037;
    wire N__34036;
    wire N__34033;
    wire N__34030;
    wire N__34025;
    wire N__34020;
    wire N__34017;
    wire N__34014;
    wire N__34011;
    wire N__34008;
    wire N__34005;
    wire N__34002;
    wire N__33999;
    wire N__33998;
    wire N__33997;
    wire N__33994;
    wire N__33991;
    wire N__33988;
    wire N__33981;
    wire N__33980;
    wire N__33979;
    wire N__33976;
    wire N__33973;
    wire N__33970;
    wire N__33967;
    wire N__33962;
    wire N__33957;
    wire N__33956;
    wire N__33955;
    wire N__33954;
    wire N__33951;
    wire N__33948;
    wire N__33945;
    wire N__33940;
    wire N__33933;
    wire N__33930;
    wire N__33929;
    wire N__33926;
    wire N__33923;
    wire N__33918;
    wire N__33917;
    wire N__33916;
    wire N__33915;
    wire N__33914;
    wire N__33913;
    wire N__33908;
    wire N__33905;
    wire N__33902;
    wire N__33899;
    wire N__33896;
    wire N__33885;
    wire N__33884;
    wire N__33881;
    wire N__33878;
    wire N__33875;
    wire N__33872;
    wire N__33871;
    wire N__33870;
    wire N__33869;
    wire N__33864;
    wire N__33859;
    wire N__33856;
    wire N__33849;
    wire N__33846;
    wire N__33843;
    wire N__33842;
    wire N__33841;
    wire N__33840;
    wire N__33837;
    wire N__33834;
    wire N__33831;
    wire N__33828;
    wire N__33823;
    wire N__33820;
    wire N__33817;
    wire N__33814;
    wire N__33811;
    wire N__33808;
    wire N__33801;
    wire N__33798;
    wire N__33795;
    wire N__33792;
    wire N__33791;
    wire N__33788;
    wire N__33787;
    wire N__33786;
    wire N__33783;
    wire N__33780;
    wire N__33777;
    wire N__33774;
    wire N__33771;
    wire N__33768;
    wire N__33765;
    wire N__33760;
    wire N__33753;
    wire N__33752;
    wire N__33751;
    wire N__33750;
    wire N__33747;
    wire N__33744;
    wire N__33741;
    wire N__33738;
    wire N__33735;
    wire N__33732;
    wire N__33723;
    wire N__33720;
    wire N__33719;
    wire N__33718;
    wire N__33715;
    wire N__33712;
    wire N__33709;
    wire N__33704;
    wire N__33703;
    wire N__33700;
    wire N__33697;
    wire N__33694;
    wire N__33693;
    wire N__33690;
    wire N__33687;
    wire N__33684;
    wire N__33681;
    wire N__33672;
    wire N__33669;
    wire N__33666;
    wire N__33665;
    wire N__33662;
    wire N__33659;
    wire N__33654;
    wire N__33653;
    wire N__33650;
    wire N__33647;
    wire N__33644;
    wire N__33641;
    wire N__33638;
    wire N__33635;
    wire N__33630;
    wire N__33629;
    wire N__33628;
    wire N__33627;
    wire N__33626;
    wire N__33625;
    wire N__33624;
    wire N__33623;
    wire N__33622;
    wire N__33621;
    wire N__33620;
    wire N__33619;
    wire N__33618;
    wire N__33617;
    wire N__33616;
    wire N__33615;
    wire N__33614;
    wire N__33613;
    wire N__33612;
    wire N__33611;
    wire N__33610;
    wire N__33609;
    wire N__33608;
    wire N__33607;
    wire N__33606;
    wire N__33605;
    wire N__33604;
    wire N__33603;
    wire N__33602;
    wire N__33601;
    wire N__33600;
    wire N__33599;
    wire N__33598;
    wire N__33531;
    wire N__33528;
    wire N__33525;
    wire N__33522;
    wire N__33519;
    wire N__33516;
    wire N__33513;
    wire N__33510;
    wire N__33509;
    wire N__33508;
    wire N__33505;
    wire N__33502;
    wire N__33499;
    wire N__33496;
    wire N__33489;
    wire N__33486;
    wire N__33483;
    wire N__33480;
    wire N__33477;
    wire N__33474;
    wire N__33471;
    wire N__33468;
    wire N__33465;
    wire N__33462;
    wire N__33459;
    wire N__33456;
    wire N__33453;
    wire N__33450;
    wire N__33447;
    wire N__33444;
    wire N__33441;
    wire N__33440;
    wire N__33439;
    wire N__33436;
    wire N__33435;
    wire N__33432;
    wire N__33429;
    wire N__33426;
    wire N__33423;
    wire N__33420;
    wire N__33417;
    wire N__33414;
    wire N__33413;
    wire N__33410;
    wire N__33409;
    wire N__33406;
    wire N__33405;
    wire N__33404;
    wire N__33401;
    wire N__33398;
    wire N__33395;
    wire N__33394;
    wire N__33393;
    wire N__33390;
    wire N__33389;
    wire N__33386;
    wire N__33383;
    wire N__33380;
    wire N__33377;
    wire N__33374;
    wire N__33369;
    wire N__33366;
    wire N__33363;
    wire N__33362;
    wire N__33359;
    wire N__33356;
    wire N__33349;
    wire N__33346;
    wire N__33345;
    wire N__33336;
    wire N__33333;
    wire N__33330;
    wire N__33325;
    wire N__33322;
    wire N__33319;
    wire N__33312;
    wire N__33307;
    wire N__33300;
    wire N__33297;
    wire N__33294;
    wire N__33291;
    wire N__33288;
    wire N__33285;
    wire N__33282;
    wire N__33279;
    wire N__33276;
    wire N__33275;
    wire N__33274;
    wire N__33271;
    wire N__33266;
    wire N__33261;
    wire N__33260;
    wire N__33257;
    wire N__33254;
    wire N__33251;
    wire N__33246;
    wire N__33245;
    wire N__33244;
    wire N__33241;
    wire N__33240;
    wire N__33237;
    wire N__33236;
    wire N__33235;
    wire N__33232;
    wire N__33231;
    wire N__33230;
    wire N__33229;
    wire N__33224;
    wire N__33219;
    wire N__33210;
    wire N__33209;
    wire N__33208;
    wire N__33205;
    wire N__33204;
    wire N__33201;
    wire N__33196;
    wire N__33191;
    wire N__33188;
    wire N__33185;
    wire N__33182;
    wire N__33181;
    wire N__33178;
    wire N__33175;
    wire N__33174;
    wire N__33173;
    wire N__33172;
    wire N__33167;
    wire N__33166;
    wire N__33165;
    wire N__33164;
    wire N__33163;
    wire N__33160;
    wire N__33157;
    wire N__33152;
    wire N__33147;
    wire N__33146;
    wire N__33143;
    wire N__33140;
    wire N__33131;
    wire N__33126;
    wire N__33121;
    wire N__33116;
    wire N__33105;
    wire N__33102;
    wire N__33099;
    wire N__33098;
    wire N__33097;
    wire N__33094;
    wire N__33091;
    wire N__33088;
    wire N__33081;
    wire N__33078;
    wire N__33077;
    wire N__33076;
    wire N__33071;
    wire N__33070;
    wire N__33069;
    wire N__33068;
    wire N__33067;
    wire N__33064;
    wire N__33061;
    wire N__33058;
    wire N__33051;
    wire N__33050;
    wire N__33049;
    wire N__33044;
    wire N__33039;
    wire N__33034;
    wire N__33027;
    wire N__33026;
    wire N__33023;
    wire N__33020;
    wire N__33015;
    wire N__33012;
    wire N__33011;
    wire N__33008;
    wire N__33005;
    wire N__33002;
    wire N__32999;
    wire N__32996;
    wire N__32993;
    wire N__32988;
    wire N__32985;
    wire N__32982;
    wire N__32981;
    wire N__32980;
    wire N__32977;
    wire N__32970;
    wire N__32967;
    wire N__32964;
    wire N__32961;
    wire N__32960;
    wire N__32957;
    wire N__32954;
    wire N__32949;
    wire N__32946;
    wire N__32943;
    wire N__32942;
    wire N__32939;
    wire N__32938;
    wire N__32935;
    wire N__32932;
    wire N__32929;
    wire N__32928;
    wire N__32923;
    wire N__32920;
    wire N__32917;
    wire N__32914;
    wire N__32911;
    wire N__32908;
    wire N__32905;
    wire N__32902;
    wire N__32899;
    wire N__32896;
    wire N__32893;
    wire N__32886;
    wire N__32883;
    wire N__32880;
    wire N__32877;
    wire N__32874;
    wire N__32871;
    wire N__32868;
    wire N__32865;
    wire N__32862;
    wire N__32859;
    wire N__32856;
    wire N__32853;
    wire N__32852;
    wire N__32849;
    wire N__32846;
    wire N__32845;
    wire N__32844;
    wire N__32839;
    wire N__32836;
    wire N__32833;
    wire N__32826;
    wire N__32823;
    wire N__32822;
    wire N__32821;
    wire N__32818;
    wire N__32815;
    wire N__32812;
    wire N__32805;
    wire N__32802;
    wire N__32799;
    wire N__32796;
    wire N__32795;
    wire N__32792;
    wire N__32789;
    wire N__32784;
    wire N__32781;
    wire N__32778;
    wire N__32775;
    wire N__32772;
    wire N__32771;
    wire N__32768;
    wire N__32765;
    wire N__32762;
    wire N__32759;
    wire N__32754;
    wire N__32751;
    wire N__32748;
    wire N__32745;
    wire N__32742;
    wire N__32741;
    wire N__32738;
    wire N__32735;
    wire N__32730;
    wire N__32727;
    wire N__32724;
    wire N__32723;
    wire N__32720;
    wire N__32717;
    wire N__32712;
    wire N__32709;
    wire N__32706;
    wire N__32703;
    wire N__32700;
    wire N__32697;
    wire N__32696;
    wire N__32693;
    wire N__32690;
    wire N__32687;
    wire N__32684;
    wire N__32681;
    wire N__32678;
    wire N__32673;
    wire N__32670;
    wire N__32667;
    wire N__32664;
    wire N__32661;
    wire N__32658;
    wire N__32655;
    wire N__32654;
    wire N__32651;
    wire N__32648;
    wire N__32643;
    wire N__32640;
    wire N__32637;
    wire N__32636;
    wire N__32635;
    wire N__32630;
    wire N__32627;
    wire N__32622;
    wire N__32619;
    wire N__32618;
    wire N__32617;
    wire N__32614;
    wire N__32611;
    wire N__32606;
    wire N__32603;
    wire N__32600;
    wire N__32595;
    wire N__32592;
    wire N__32589;
    wire N__32588;
    wire N__32585;
    wire N__32582;
    wire N__32577;
    wire N__32574;
    wire N__32571;
    wire N__32570;
    wire N__32569;
    wire N__32566;
    wire N__32559;
    wire N__32556;
    wire N__32553;
    wire N__32550;
    wire N__32547;
    wire N__32544;
    wire N__32543;
    wire N__32542;
    wire N__32539;
    wire N__32534;
    wire N__32529;
    wire N__32528;
    wire N__32525;
    wire N__32522;
    wire N__32519;
    wire N__32516;
    wire N__32513;
    wire N__32510;
    wire N__32505;
    wire N__32502;
    wire N__32499;
    wire N__32496;
    wire N__32493;
    wire N__32492;
    wire N__32489;
    wire N__32486;
    wire N__32483;
    wire N__32480;
    wire N__32477;
    wire N__32474;
    wire N__32471;
    wire N__32468;
    wire N__32463;
    wire N__32460;
    wire N__32457;
    wire N__32454;
    wire N__32451;
    wire N__32450;
    wire N__32447;
    wire N__32444;
    wire N__32441;
    wire N__32438;
    wire N__32435;
    wire N__32432;
    wire N__32427;
    wire N__32424;
    wire N__32421;
    wire N__32418;
    wire N__32415;
    wire N__32412;
    wire N__32409;
    wire N__32406;
    wire N__32405;
    wire N__32404;
    wire N__32403;
    wire N__32402;
    wire N__32401;
    wire N__32400;
    wire N__32385;
    wire N__32382;
    wire N__32379;
    wire N__32376;
    wire N__32373;
    wire N__32370;
    wire N__32367;
    wire N__32366;
    wire N__32365;
    wire N__32358;
    wire N__32355;
    wire N__32352;
    wire N__32351;
    wire N__32348;
    wire N__32345;
    wire N__32342;
    wire N__32339;
    wire N__32336;
    wire N__32333;
    wire N__32328;
    wire N__32325;
    wire N__32322;
    wire N__32319;
    wire N__32316;
    wire N__32315;
    wire N__32314;
    wire N__32311;
    wire N__32304;
    wire N__32301;
    wire N__32298;
    wire N__32295;
    wire N__32292;
    wire N__32289;
    wire N__32286;
    wire N__32285;
    wire N__32284;
    wire N__32279;
    wire N__32278;
    wire N__32275;
    wire N__32272;
    wire N__32269;
    wire N__32264;
    wire N__32259;
    wire N__32256;
    wire N__32253;
    wire N__32252;
    wire N__32247;
    wire N__32244;
    wire N__32241;
    wire N__32238;
    wire N__32235;
    wire N__32232;
    wire N__32231;
    wire N__32226;
    wire N__32223;
    wire N__32220;
    wire N__32217;
    wire N__32214;
    wire N__32211;
    wire N__32210;
    wire N__32205;
    wire N__32202;
    wire N__32199;
    wire N__32196;
    wire N__32193;
    wire N__32190;
    wire N__32189;
    wire N__32184;
    wire N__32181;
    wire N__32178;
    wire N__32175;
    wire N__32172;
    wire N__32169;
    wire N__32168;
    wire N__32163;
    wire N__32160;
    wire N__32157;
    wire N__32154;
    wire N__32151;
    wire N__32148;
    wire N__32147;
    wire N__32142;
    wire N__32139;
    wire N__32136;
    wire N__32133;
    wire N__32130;
    wire N__32129;
    wire N__32126;
    wire N__32125;
    wire N__32124;
    wire N__32123;
    wire N__32122;
    wire N__32121;
    wire N__32120;
    wire N__32119;
    wire N__32118;
    wire N__32117;
    wire N__32110;
    wire N__32103;
    wire N__32096;
    wire N__32091;
    wire N__32082;
    wire N__32081;
    wire N__32080;
    wire N__32077;
    wire N__32076;
    wire N__32075;
    wire N__32074;
    wire N__32073;
    wire N__32072;
    wire N__32071;
    wire N__32068;
    wire N__32067;
    wire N__32062;
    wire N__32055;
    wire N__32048;
    wire N__32043;
    wire N__32034;
    wire N__32033;
    wire N__32032;
    wire N__32031;
    wire N__32030;
    wire N__32029;
    wire N__32026;
    wire N__32025;
    wire N__32024;
    wire N__32023;
    wire N__32020;
    wire N__32013;
    wire N__32006;
    wire N__32001;
    wire N__31992;
    wire N__31989;
    wire N__31986;
    wire N__31983;
    wire N__31980;
    wire N__31977;
    wire N__31974;
    wire N__31971;
    wire N__31970;
    wire N__31969;
    wire N__31966;
    wire N__31961;
    wire N__31956;
    wire N__31953;
    wire N__31950;
    wire N__31947;
    wire N__31944;
    wire N__31943;
    wire N__31940;
    wire N__31937;
    wire N__31934;
    wire N__31931;
    wire N__31928;
    wire N__31925;
    wire N__31920;
    wire N__31919;
    wire N__31918;
    wire N__31915;
    wire N__31908;
    wire N__31905;
    wire N__31902;
    wire N__31899;
    wire N__31896;
    wire N__31893;
    wire N__31892;
    wire N__31889;
    wire N__31886;
    wire N__31883;
    wire N__31880;
    wire N__31877;
    wire N__31874;
    wire N__31869;
    wire N__31866;
    wire N__31863;
    wire N__31860;
    wire N__31857;
    wire N__31854;
    wire N__31851;
    wire N__31850;
    wire N__31849;
    wire N__31846;
    wire N__31843;
    wire N__31842;
    wire N__31839;
    wire N__31836;
    wire N__31829;
    wire N__31828;
    wire N__31825;
    wire N__31822;
    wire N__31819;
    wire N__31814;
    wire N__31811;
    wire N__31810;
    wire N__31807;
    wire N__31804;
    wire N__31801;
    wire N__31796;
    wire N__31791;
    wire N__31788;
    wire N__31785;
    wire N__31782;
    wire N__31779;
    wire N__31776;
    wire N__31773;
    wire N__31772;
    wire N__31769;
    wire N__31768;
    wire N__31765;
    wire N__31762;
    wire N__31759;
    wire N__31754;
    wire N__31749;
    wire N__31748;
    wire N__31747;
    wire N__31746;
    wire N__31739;
    wire N__31736;
    wire N__31731;
    wire N__31728;
    wire N__31725;
    wire N__31724;
    wire N__31723;
    wire N__31722;
    wire N__31721;
    wire N__31718;
    wire N__31715;
    wire N__31712;
    wire N__31711;
    wire N__31710;
    wire N__31709;
    wire N__31704;
    wire N__31699;
    wire N__31696;
    wire N__31693;
    wire N__31688;
    wire N__31683;
    wire N__31680;
    wire N__31671;
    wire N__31670;
    wire N__31665;
    wire N__31662;
    wire N__31659;
    wire N__31658;
    wire N__31655;
    wire N__31652;
    wire N__31647;
    wire N__31644;
    wire N__31643;
    wire N__31642;
    wire N__31639;
    wire N__31634;
    wire N__31631;
    wire N__31628;
    wire N__31623;
    wire N__31620;
    wire N__31619;
    wire N__31616;
    wire N__31615;
    wire N__31612;
    wire N__31611;
    wire N__31608;
    wire N__31607;
    wire N__31606;
    wire N__31605;
    wire N__31602;
    wire N__31601;
    wire N__31598;
    wire N__31595;
    wire N__31592;
    wire N__31589;
    wire N__31584;
    wire N__31579;
    wire N__31576;
    wire N__31563;
    wire N__31562;
    wire N__31559;
    wire N__31556;
    wire N__31555;
    wire N__31554;
    wire N__31551;
    wire N__31548;
    wire N__31547;
    wire N__31546;
    wire N__31543;
    wire N__31540;
    wire N__31535;
    wire N__31530;
    wire N__31521;
    wire N__31520;
    wire N__31519;
    wire N__31516;
    wire N__31513;
    wire N__31510;
    wire N__31509;
    wire N__31506;
    wire N__31505;
    wire N__31504;
    wire N__31503;
    wire N__31500;
    wire N__31497;
    wire N__31494;
    wire N__31491;
    wire N__31490;
    wire N__31489;
    wire N__31486;
    wire N__31483;
    wire N__31480;
    wire N__31473;
    wire N__31470;
    wire N__31463;
    wire N__31452;
    wire N__31449;
    wire N__31448;
    wire N__31445;
    wire N__31442;
    wire N__31437;
    wire N__31436;
    wire N__31435;
    wire N__31434;
    wire N__31433;
    wire N__31432;
    wire N__31431;
    wire N__31430;
    wire N__31413;
    wire N__31410;
    wire N__31407;
    wire N__31404;
    wire N__31401;
    wire N__31398;
    wire N__31397;
    wire N__31394;
    wire N__31393;
    wire N__31392;
    wire N__31391;
    wire N__31390;
    wire N__31389;
    wire N__31388;
    wire N__31385;
    wire N__31384;
    wire N__31383;
    wire N__31382;
    wire N__31379;
    wire N__31376;
    wire N__31373;
    wire N__31372;
    wire N__31371;
    wire N__31370;
    wire N__31359;
    wire N__31352;
    wire N__31345;
    wire N__31342;
    wire N__31339;
    wire N__31336;
    wire N__31331;
    wire N__31326;
    wire N__31323;
    wire N__31320;
    wire N__31315;
    wire N__31310;
    wire N__31305;
    wire N__31302;
    wire N__31301;
    wire N__31300;
    wire N__31297;
    wire N__31294;
    wire N__31289;
    wire N__31286;
    wire N__31283;
    wire N__31278;
    wire N__31275;
    wire N__31272;
    wire N__31271;
    wire N__31268;
    wire N__31265;
    wire N__31260;
    wire N__31257;
    wire N__31254;
    wire N__31251;
    wire N__31248;
    wire N__31245;
    wire N__31244;
    wire N__31241;
    wire N__31238;
    wire N__31233;
    wire N__31230;
    wire N__31229;
    wire N__31228;
    wire N__31227;
    wire N__31226;
    wire N__31225;
    wire N__31224;
    wire N__31223;
    wire N__31222;
    wire N__31221;
    wire N__31220;
    wire N__31217;
    wire N__31216;
    wire N__31213;
    wire N__31212;
    wire N__31209;
    wire N__31200;
    wire N__31191;
    wire N__31188;
    wire N__31185;
    wire N__31182;
    wire N__31179;
    wire N__31178;
    wire N__31175;
    wire N__31170;
    wire N__31165;
    wire N__31162;
    wire N__31159;
    wire N__31156;
    wire N__31149;
    wire N__31144;
    wire N__31141;
    wire N__31134;
    wire N__31131;
    wire N__31130;
    wire N__31129;
    wire N__31126;
    wire N__31123;
    wire N__31118;
    wire N__31113;
    wire N__31112;
    wire N__31109;
    wire N__31108;
    wire N__31105;
    wire N__31102;
    wire N__31101;
    wire N__31098;
    wire N__31095;
    wire N__31092;
    wire N__31089;
    wire N__31084;
    wire N__31081;
    wire N__31074;
    wire N__31073;
    wire N__31072;
    wire N__31069;
    wire N__31068;
    wire N__31067;
    wire N__31064;
    wire N__31061;
    wire N__31060;
    wire N__31053;
    wire N__31052;
    wire N__31047;
    wire N__31044;
    wire N__31043;
    wire N__31040;
    wire N__31037;
    wire N__31032;
    wire N__31029;
    wire N__31020;
    wire N__31019;
    wire N__31016;
    wire N__31013;
    wire N__31010;
    wire N__31007;
    wire N__31002;
    wire N__31001;
    wire N__31000;
    wire N__30999;
    wire N__30996;
    wire N__30993;
    wire N__30992;
    wire N__30991;
    wire N__30990;
    wire N__30987;
    wire N__30984;
    wire N__30981;
    wire N__30978;
    wire N__30975;
    wire N__30970;
    wire N__30967;
    wire N__30962;
    wire N__30951;
    wire N__30950;
    wire N__30945;
    wire N__30944;
    wire N__30941;
    wire N__30938;
    wire N__30935;
    wire N__30932;
    wire N__30929;
    wire N__30926;
    wire N__30923;
    wire N__30918;
    wire N__30915;
    wire N__30914;
    wire N__30913;
    wire N__30908;
    wire N__30905;
    wire N__30902;
    wire N__30899;
    wire N__30896;
    wire N__30891;
    wire N__30888;
    wire N__30885;
    wire N__30882;
    wire N__30881;
    wire N__30876;
    wire N__30875;
    wire N__30872;
    wire N__30869;
    wire N__30866;
    wire N__30863;
    wire N__30860;
    wire N__30857;
    wire N__30854;
    wire N__30849;
    wire N__30846;
    wire N__30845;
    wire N__30840;
    wire N__30839;
    wire N__30836;
    wire N__30833;
    wire N__30830;
    wire N__30827;
    wire N__30824;
    wire N__30821;
    wire N__30818;
    wire N__30813;
    wire N__30810;
    wire N__30809;
    wire N__30804;
    wire N__30801;
    wire N__30800;
    wire N__30797;
    wire N__30794;
    wire N__30791;
    wire N__30788;
    wire N__30785;
    wire N__30782;
    wire N__30779;
    wire N__30774;
    wire N__30771;
    wire N__30770;
    wire N__30767;
    wire N__30766;
    wire N__30763;
    wire N__30760;
    wire N__30757;
    wire N__30754;
    wire N__30751;
    wire N__30748;
    wire N__30745;
    wire N__30742;
    wire N__30739;
    wire N__30736;
    wire N__30733;
    wire N__30726;
    wire N__30723;
    wire N__30720;
    wire N__30719;
    wire N__30718;
    wire N__30717;
    wire N__30714;
    wire N__30707;
    wire N__30706;
    wire N__30705;
    wire N__30704;
    wire N__30703;
    wire N__30702;
    wire N__30701;
    wire N__30700;
    wire N__30699;
    wire N__30698;
    wire N__30697;
    wire N__30696;
    wire N__30695;
    wire N__30694;
    wire N__30691;
    wire N__30690;
    wire N__30687;
    wire N__30684;
    wire N__30681;
    wire N__30676;
    wire N__30667;
    wire N__30664;
    wire N__30655;
    wire N__30652;
    wire N__30651;
    wire N__30648;
    wire N__30645;
    wire N__30642;
    wire N__30639;
    wire N__30636;
    wire N__30629;
    wire N__30626;
    wire N__30623;
    wire N__30618;
    wire N__30615;
    wire N__30612;
    wire N__30607;
    wire N__30604;
    wire N__30601;
    wire N__30598;
    wire N__30593;
    wire N__30590;
    wire N__30579;
    wire N__30578;
    wire N__30577;
    wire N__30574;
    wire N__30571;
    wire N__30568;
    wire N__30567;
    wire N__30566;
    wire N__30563;
    wire N__30560;
    wire N__30557;
    wire N__30552;
    wire N__30549;
    wire N__30546;
    wire N__30543;
    wire N__30540;
    wire N__30537;
    wire N__30534;
    wire N__30529;
    wire N__30528;
    wire N__30525;
    wire N__30520;
    wire N__30517;
    wire N__30514;
    wire N__30507;
    wire N__30504;
    wire N__30501;
    wire N__30498;
    wire N__30495;
    wire N__30494;
    wire N__30491;
    wire N__30488;
    wire N__30485;
    wire N__30480;
    wire N__30479;
    wire N__30476;
    wire N__30475;
    wire N__30472;
    wire N__30469;
    wire N__30466;
    wire N__30463;
    wire N__30460;
    wire N__30455;
    wire N__30452;
    wire N__30447;
    wire N__30444;
    wire N__30443;
    wire N__30440;
    wire N__30437;
    wire N__30432;
    wire N__30431;
    wire N__30426;
    wire N__30423;
    wire N__30422;
    wire N__30419;
    wire N__30416;
    wire N__30413;
    wire N__30410;
    wire N__30407;
    wire N__30402;
    wire N__30399;
    wire N__30396;
    wire N__30395;
    wire N__30392;
    wire N__30389;
    wire N__30386;
    wire N__30383;
    wire N__30378;
    wire N__30377;
    wire N__30376;
    wire N__30371;
    wire N__30368;
    wire N__30365;
    wire N__30360;
    wire N__30357;
    wire N__30354;
    wire N__30351;
    wire N__30350;
    wire N__30347;
    wire N__30344;
    wire N__30339;
    wire N__30338;
    wire N__30335;
    wire N__30334;
    wire N__30331;
    wire N__30328;
    wire N__30325;
    wire N__30320;
    wire N__30317;
    wire N__30314;
    wire N__30311;
    wire N__30308;
    wire N__30303;
    wire N__30300;
    wire N__30299;
    wire N__30298;
    wire N__30293;
    wire N__30290;
    wire N__30287;
    wire N__30284;
    wire N__30281;
    wire N__30278;
    wire N__30275;
    wire N__30270;
    wire N__30267;
    wire N__30266;
    wire N__30263;
    wire N__30260;
    wire N__30255;
    wire N__30254;
    wire N__30251;
    wire N__30250;
    wire N__30247;
    wire N__30244;
    wire N__30241;
    wire N__30238;
    wire N__30233;
    wire N__30230;
    wire N__30227;
    wire N__30222;
    wire N__30219;
    wire N__30216;
    wire N__30215;
    wire N__30214;
    wire N__30211;
    wire N__30206;
    wire N__30203;
    wire N__30200;
    wire N__30197;
    wire N__30194;
    wire N__30189;
    wire N__30186;
    wire N__30185;
    wire N__30180;
    wire N__30179;
    wire N__30176;
    wire N__30173;
    wire N__30170;
    wire N__30167;
    wire N__30164;
    wire N__30159;
    wire N__30156;
    wire N__30153;
    wire N__30150;
    wire N__30147;
    wire N__30144;
    wire N__30141;
    wire N__30138;
    wire N__30137;
    wire N__30134;
    wire N__30131;
    wire N__30128;
    wire N__30125;
    wire N__30120;
    wire N__30117;
    wire N__30114;
    wire N__30111;
    wire N__30108;
    wire N__30105;
    wire N__30102;
    wire N__30101;
    wire N__30098;
    wire N__30095;
    wire N__30092;
    wire N__30089;
    wire N__30086;
    wire N__30085;
    wire N__30082;
    wire N__30079;
    wire N__30076;
    wire N__30073;
    wire N__30070;
    wire N__30067;
    wire N__30064;
    wire N__30061;
    wire N__30058;
    wire N__30055;
    wire N__30048;
    wire N__30045;
    wire N__30042;
    wire N__30039;
    wire N__30036;
    wire N__30035;
    wire N__30032;
    wire N__30029;
    wire N__30028;
    wire N__30025;
    wire N__30022;
    wire N__30019;
    wire N__30014;
    wire N__30009;
    wire N__30006;
    wire N__30003;
    wire N__30000;
    wire N__29997;
    wire N__29996;
    wire N__29993;
    wire N__29990;
    wire N__29989;
    wire N__29986;
    wire N__29983;
    wire N__29980;
    wire N__29975;
    wire N__29972;
    wire N__29969;
    wire N__29964;
    wire N__29961;
    wire N__29958;
    wire N__29955;
    wire N__29952;
    wire N__29949;
    wire N__29948;
    wire N__29947;
    wire N__29940;
    wire N__29937;
    wire N__29934;
    wire N__29931;
    wire N__29928;
    wire N__29925;
    wire N__29924;
    wire N__29921;
    wire N__29918;
    wire N__29915;
    wire N__29910;
    wire N__29907;
    wire N__29906;
    wire N__29905;
    wire N__29902;
    wire N__29897;
    wire N__29894;
    wire N__29891;
    wire N__29886;
    wire N__29883;
    wire N__29880;
    wire N__29879;
    wire N__29874;
    wire N__29871;
    wire N__29870;
    wire N__29867;
    wire N__29864;
    wire N__29861;
    wire N__29858;
    wire N__29855;
    wire N__29850;
    wire N__29847;
    wire N__29844;
    wire N__29841;
    wire N__29838;
    wire N__29835;
    wire N__29834;
    wire N__29831;
    wire N__29828;
    wire N__29825;
    wire N__29820;
    wire N__29817;
    wire N__29814;
    wire N__29811;
    wire N__29808;
    wire N__29805;
    wire N__29802;
    wire N__29799;
    wire N__29796;
    wire N__29793;
    wire N__29790;
    wire N__29789;
    wire N__29786;
    wire N__29783;
    wire N__29778;
    wire N__29777;
    wire N__29774;
    wire N__29771;
    wire N__29766;
    wire N__29763;
    wire N__29760;
    wire N__29757;
    wire N__29754;
    wire N__29753;
    wire N__29750;
    wire N__29747;
    wire N__29742;
    wire N__29739;
    wire N__29736;
    wire N__29733;
    wire N__29730;
    wire N__29727;
    wire N__29724;
    wire N__29721;
    wire N__29718;
    wire N__29715;
    wire N__29714;
    wire N__29713;
    wire N__29712;
    wire N__29709;
    wire N__29706;
    wire N__29705;
    wire N__29704;
    wire N__29701;
    wire N__29698;
    wire N__29695;
    wire N__29688;
    wire N__29683;
    wire N__29676;
    wire N__29673;
    wire N__29672;
    wire N__29669;
    wire N__29668;
    wire N__29667;
    wire N__29664;
    wire N__29663;
    wire N__29662;
    wire N__29661;
    wire N__29658;
    wire N__29657;
    wire N__29654;
    wire N__29651;
    wire N__29648;
    wire N__29647;
    wire N__29644;
    wire N__29643;
    wire N__29642;
    wire N__29637;
    wire N__29634;
    wire N__29631;
    wire N__29628;
    wire N__29623;
    wire N__29614;
    wire N__29601;
    wire N__29600;
    wire N__29597;
    wire N__29594;
    wire N__29591;
    wire N__29590;
    wire N__29587;
    wire N__29584;
    wire N__29581;
    wire N__29578;
    wire N__29577;
    wire N__29572;
    wire N__29569;
    wire N__29566;
    wire N__29563;
    wire N__29556;
    wire N__29553;
    wire N__29552;
    wire N__29551;
    wire N__29550;
    wire N__29547;
    wire N__29544;
    wire N__29541;
    wire N__29538;
    wire N__29535;
    wire N__29532;
    wire N__29529;
    wire N__29526;
    wire N__29517;
    wire N__29514;
    wire N__29513;
    wire N__29512;
    wire N__29509;
    wire N__29506;
    wire N__29503;
    wire N__29500;
    wire N__29497;
    wire N__29494;
    wire N__29493;
    wire N__29488;
    wire N__29485;
    wire N__29482;
    wire N__29475;
    wire N__29474;
    wire N__29471;
    wire N__29468;
    wire N__29465;
    wire N__29462;
    wire N__29457;
    wire N__29454;
    wire N__29453;
    wire N__29450;
    wire N__29447;
    wire N__29444;
    wire N__29441;
    wire N__29436;
    wire N__29435;
    wire N__29432;
    wire N__29429;
    wire N__29424;
    wire N__29421;
    wire N__29418;
    wire N__29415;
    wire N__29412;
    wire N__29409;
    wire N__29406;
    wire N__29403;
    wire N__29400;
    wire N__29397;
    wire N__29396;
    wire N__29393;
    wire N__29392;
    wire N__29389;
    wire N__29386;
    wire N__29383;
    wire N__29380;
    wire N__29377;
    wire N__29374;
    wire N__29367;
    wire N__29364;
    wire N__29361;
    wire N__29358;
    wire N__29355;
    wire N__29352;
    wire N__29349;
    wire N__29346;
    wire N__29345;
    wire N__29342;
    wire N__29341;
    wire N__29338;
    wire N__29335;
    wire N__29332;
    wire N__29329;
    wire N__29324;
    wire N__29319;
    wire N__29316;
    wire N__29313;
    wire N__29310;
    wire N__29307;
    wire N__29304;
    wire N__29301;
    wire N__29300;
    wire N__29297;
    wire N__29296;
    wire N__29293;
    wire N__29290;
    wire N__29287;
    wire N__29284;
    wire N__29281;
    wire N__29278;
    wire N__29271;
    wire N__29268;
    wire N__29265;
    wire N__29262;
    wire N__29259;
    wire N__29258;
    wire N__29255;
    wire N__29252;
    wire N__29249;
    wire N__29246;
    wire N__29243;
    wire N__29240;
    wire N__29235;
    wire N__29232;
    wire N__29229;
    wire N__29226;
    wire N__29223;
    wire N__29220;
    wire N__29217;
    wire N__29214;
    wire N__29211;
    wire N__29208;
    wire N__29205;
    wire N__29202;
    wire N__29199;
    wire N__29196;
    wire N__29193;
    wire N__29190;
    wire N__29187;
    wire N__29184;
    wire N__29181;
    wire N__29180;
    wire N__29177;
    wire N__29174;
    wire N__29171;
    wire N__29168;
    wire N__29163;
    wire N__29160;
    wire N__29157;
    wire N__29156;
    wire N__29153;
    wire N__29150;
    wire N__29147;
    wire N__29144;
    wire N__29139;
    wire N__29136;
    wire N__29133;
    wire N__29130;
    wire N__29127;
    wire N__29124;
    wire N__29123;
    wire N__29120;
    wire N__29117;
    wire N__29114;
    wire N__29109;
    wire N__29106;
    wire N__29103;
    wire N__29100;
    wire N__29097;
    wire N__29094;
    wire N__29091;
    wire N__29088;
    wire N__29085;
    wire N__29082;
    wire N__29081;
    wire N__29080;
    wire N__29079;
    wire N__29076;
    wire N__29073;
    wire N__29070;
    wire N__29067;
    wire N__29064;
    wire N__29061;
    wire N__29052;
    wire N__29051;
    wire N__29048;
    wire N__29045;
    wire N__29044;
    wire N__29039;
    wire N__29036;
    wire N__29035;
    wire N__29032;
    wire N__29029;
    wire N__29026;
    wire N__29019;
    wire N__29016;
    wire N__29015;
    wire N__29014;
    wire N__29011;
    wire N__29008;
    wire N__29007;
    wire N__29004;
    wire N__29001;
    wire N__28996;
    wire N__28989;
    wire N__28988;
    wire N__28985;
    wire N__28982;
    wire N__28981;
    wire N__28980;
    wire N__28975;
    wire N__28972;
    wire N__28969;
    wire N__28966;
    wire N__28963;
    wire N__28960;
    wire N__28953;
    wire N__28952;
    wire N__28949;
    wire N__28946;
    wire N__28945;
    wire N__28944;
    wire N__28939;
    wire N__28936;
    wire N__28933;
    wire N__28930;
    wire N__28927;
    wire N__28924;
    wire N__28917;
    wire N__28914;
    wire N__28913;
    wire N__28910;
    wire N__28909;
    wire N__28906;
    wire N__28903;
    wire N__28900;
    wire N__28899;
    wire N__28896;
    wire N__28893;
    wire N__28888;
    wire N__28881;
    wire N__28878;
    wire N__28875;
    wire N__28874;
    wire N__28871;
    wire N__28868;
    wire N__28865;
    wire N__28862;
    wire N__28857;
    wire N__28854;
    wire N__28853;
    wire N__28850;
    wire N__28847;
    wire N__28842;
    wire N__28841;
    wire N__28838;
    wire N__28835;
    wire N__28832;
    wire N__28829;
    wire N__28824;
    wire N__28821;
    wire N__28818;
    wire N__28817;
    wire N__28814;
    wire N__28811;
    wire N__28808;
    wire N__28805;
    wire N__28800;
    wire N__28799;
    wire N__28796;
    wire N__28793;
    wire N__28790;
    wire N__28787;
    wire N__28782;
    wire N__28781;
    wire N__28778;
    wire N__28775;
    wire N__28772;
    wire N__28767;
    wire N__28766;
    wire N__28765;
    wire N__28764;
    wire N__28763;
    wire N__28762;
    wire N__28761;
    wire N__28760;
    wire N__28743;
    wire N__28740;
    wire N__28737;
    wire N__28734;
    wire N__28733;
    wire N__28732;
    wire N__28729;
    wire N__28724;
    wire N__28719;
    wire N__28718;
    wire N__28717;
    wire N__28714;
    wire N__28711;
    wire N__28708;
    wire N__28703;
    wire N__28698;
    wire N__28697;
    wire N__28696;
    wire N__28691;
    wire N__28688;
    wire N__28683;
    wire N__28680;
    wire N__28677;
    wire N__28674;
    wire N__28673;
    wire N__28672;
    wire N__28669;
    wire N__28668;
    wire N__28667;
    wire N__28664;
    wire N__28661;
    wire N__28660;
    wire N__28649;
    wire N__28646;
    wire N__28641;
    wire N__28638;
    wire N__28637;
    wire N__28636;
    wire N__28633;
    wire N__28630;
    wire N__28627;
    wire N__28626;
    wire N__28621;
    wire N__28618;
    wire N__28615;
    wire N__28608;
    wire N__28605;
    wire N__28602;
    wire N__28599;
    wire N__28596;
    wire N__28595;
    wire N__28594;
    wire N__28591;
    wire N__28588;
    wire N__28585;
    wire N__28578;
    wire N__28575;
    wire N__28574;
    wire N__28573;
    wire N__28570;
    wire N__28565;
    wire N__28560;
    wire N__28557;
    wire N__28554;
    wire N__28553;
    wire N__28552;
    wire N__28549;
    wire N__28544;
    wire N__28539;
    wire N__28536;
    wire N__28535;
    wire N__28530;
    wire N__28527;
    wire N__28524;
    wire N__28523;
    wire N__28522;
    wire N__28521;
    wire N__28520;
    wire N__28517;
    wire N__28508;
    wire N__28507;
    wire N__28502;
    wire N__28499;
    wire N__28494;
    wire N__28491;
    wire N__28488;
    wire N__28487;
    wire N__28484;
    wire N__28481;
    wire N__28478;
    wire N__28473;
    wire N__28470;
    wire N__28467;
    wire N__28466;
    wire N__28463;
    wire N__28460;
    wire N__28457;
    wire N__28454;
    wire N__28451;
    wire N__28448;
    wire N__28443;
    wire N__28440;
    wire N__28437;
    wire N__28434;
    wire N__28431;
    wire N__28428;
    wire N__28425;
    wire N__28422;
    wire N__28419;
    wire N__28416;
    wire N__28413;
    wire N__28410;
    wire N__28407;
    wire N__28404;
    wire N__28403;
    wire N__28402;
    wire N__28401;
    wire N__28392;
    wire N__28389;
    wire N__28388;
    wire N__28385;
    wire N__28382;
    wire N__28379;
    wire N__28374;
    wire N__28371;
    wire N__28368;
    wire N__28365;
    wire N__28362;
    wire N__28359;
    wire N__28356;
    wire N__28353;
    wire N__28350;
    wire N__28347;
    wire N__28344;
    wire N__28341;
    wire N__28340;
    wire N__28335;
    wire N__28332;
    wire N__28329;
    wire N__28326;
    wire N__28325;
    wire N__28320;
    wire N__28317;
    wire N__28314;
    wire N__28311;
    wire N__28310;
    wire N__28305;
    wire N__28302;
    wire N__28299;
    wire N__28296;
    wire N__28295;
    wire N__28290;
    wire N__28287;
    wire N__28284;
    wire N__28281;
    wire N__28280;
    wire N__28275;
    wire N__28272;
    wire N__28269;
    wire N__28266;
    wire N__28265;
    wire N__28260;
    wire N__28257;
    wire N__28254;
    wire N__28253;
    wire N__28250;
    wire N__28247;
    wire N__28242;
    wire N__28239;
    wire N__28236;
    wire N__28233;
    wire N__28230;
    wire N__28227;
    wire N__28226;
    wire N__28221;
    wire N__28218;
    wire N__28215;
    wire N__28212;
    wire N__28211;
    wire N__28206;
    wire N__28203;
    wire N__28200;
    wire N__28197;
    wire N__28196;
    wire N__28191;
    wire N__28188;
    wire N__28185;
    wire N__28182;
    wire N__28181;
    wire N__28176;
    wire N__28173;
    wire N__28170;
    wire N__28167;
    wire N__28166;
    wire N__28161;
    wire N__28158;
    wire N__28155;
    wire N__28152;
    wire N__28151;
    wire N__28146;
    wire N__28143;
    wire N__28140;
    wire N__28139;
    wire N__28136;
    wire N__28133;
    wire N__28128;
    wire N__28125;
    wire N__28122;
    wire N__28119;
    wire N__28116;
    wire N__28113;
    wire N__28110;
    wire N__28107;
    wire N__28104;
    wire N__28103;
    wire N__28100;
    wire N__28097;
    wire N__28092;
    wire N__28091;
    wire N__28088;
    wire N__28085;
    wire N__28080;
    wire N__28077;
    wire N__28074;
    wire N__28073;
    wire N__28072;
    wire N__28069;
    wire N__28068;
    wire N__28067;
    wire N__28066;
    wire N__28065;
    wire N__28062;
    wire N__28059;
    wire N__28058;
    wire N__28057;
    wire N__28054;
    wire N__28051;
    wire N__28048;
    wire N__28047;
    wire N__28044;
    wire N__28043;
    wire N__28032;
    wire N__28027;
    wire N__28022;
    wire N__28019;
    wire N__28016;
    wire N__28011;
    wire N__28008;
    wire N__28005;
    wire N__28002;
    wire N__27999;
    wire N__27992;
    wire N__27987;
    wire N__27984;
    wire N__27981;
    wire N__27980;
    wire N__27979;
    wire N__27978;
    wire N__27977;
    wire N__27976;
    wire N__27975;
    wire N__27972;
    wire N__27969;
    wire N__27958;
    wire N__27951;
    wire N__27948;
    wire N__27947;
    wire N__27944;
    wire N__27941;
    wire N__27940;
    wire N__27937;
    wire N__27934;
    wire N__27931;
    wire N__27928;
    wire N__27923;
    wire N__27918;
    wire N__27917;
    wire N__27914;
    wire N__27913;
    wire N__27912;
    wire N__27909;
    wire N__27906;
    wire N__27903;
    wire N__27900;
    wire N__27897;
    wire N__27894;
    wire N__27891;
    wire N__27888;
    wire N__27885;
    wire N__27876;
    wire N__27875;
    wire N__27872;
    wire N__27869;
    wire N__27866;
    wire N__27865;
    wire N__27864;
    wire N__27863;
    wire N__27862;
    wire N__27859;
    wire N__27856;
    wire N__27853;
    wire N__27850;
    wire N__27847;
    wire N__27844;
    wire N__27841;
    wire N__27838;
    wire N__27825;
    wire N__27822;
    wire N__27819;
    wire N__27816;
    wire N__27813;
    wire N__27810;
    wire N__27807;
    wire N__27804;
    wire N__27801;
    wire N__27798;
    wire N__27795;
    wire N__27792;
    wire N__27789;
    wire N__27786;
    wire N__27783;
    wire N__27780;
    wire N__27777;
    wire N__27774;
    wire N__27771;
    wire N__27768;
    wire N__27765;
    wire N__27762;
    wire N__27759;
    wire N__27756;
    wire N__27753;
    wire N__27750;
    wire N__27747;
    wire N__27744;
    wire N__27741;
    wire N__27738;
    wire N__27735;
    wire N__27732;
    wire N__27729;
    wire N__27726;
    wire N__27723;
    wire N__27720;
    wire N__27717;
    wire N__27714;
    wire N__27711;
    wire N__27708;
    wire N__27705;
    wire N__27702;
    wire N__27699;
    wire N__27696;
    wire N__27693;
    wire N__27690;
    wire N__27687;
    wire N__27684;
    wire N__27681;
    wire N__27678;
    wire N__27677;
    wire N__27674;
    wire N__27673;
    wire N__27670;
    wire N__27669;
    wire N__27666;
    wire N__27663;
    wire N__27662;
    wire N__27659;
    wire N__27656;
    wire N__27655;
    wire N__27654;
    wire N__27653;
    wire N__27652;
    wire N__27651;
    wire N__27646;
    wire N__27643;
    wire N__27640;
    wire N__27637;
    wire N__27634;
    wire N__27631;
    wire N__27628;
    wire N__27625;
    wire N__27622;
    wire N__27617;
    wire N__27616;
    wire N__27615;
    wire N__27614;
    wire N__27613;
    wire N__27610;
    wire N__27603;
    wire N__27600;
    wire N__27595;
    wire N__27592;
    wire N__27587;
    wire N__27582;
    wire N__27567;
    wire N__27564;
    wire N__27561;
    wire N__27558;
    wire N__27555;
    wire N__27554;
    wire N__27553;
    wire N__27552;
    wire N__27551;
    wire N__27548;
    wire N__27547;
    wire N__27544;
    wire N__27539;
    wire N__27536;
    wire N__27531;
    wire N__27522;
    wire N__27519;
    wire N__27516;
    wire N__27513;
    wire N__27510;
    wire N__27507;
    wire N__27504;
    wire N__27501;
    wire N__27498;
    wire N__27495;
    wire N__27494;
    wire N__27491;
    wire N__27490;
    wire N__27487;
    wire N__27482;
    wire N__27477;
    wire N__27474;
    wire N__27471;
    wire N__27468;
    wire N__27467;
    wire N__27464;
    wire N__27463;
    wire N__27462;
    wire N__27459;
    wire N__27454;
    wire N__27449;
    wire N__27444;
    wire N__27441;
    wire N__27438;
    wire N__27435;
    wire N__27432;
    wire N__27429;
    wire N__27426;
    wire N__27423;
    wire N__27420;
    wire N__27417;
    wire N__27414;
    wire N__27411;
    wire N__27408;
    wire N__27405;
    wire N__27402;
    wire N__27399;
    wire N__27396;
    wire N__27393;
    wire N__27390;
    wire N__27387;
    wire N__27384;
    wire N__27381;
    wire N__27378;
    wire N__27377;
    wire N__27372;
    wire N__27369;
    wire N__27366;
    wire N__27365;
    wire N__27360;
    wire N__27357;
    wire N__27354;
    wire N__27351;
    wire N__27348;
    wire N__27345;
    wire N__27342;
    wire N__27341;
    wire N__27338;
    wire N__27335;
    wire N__27330;
    wire N__27327;
    wire N__27324;
    wire N__27321;
    wire N__27318;
    wire N__27315;
    wire N__27312;
    wire N__27309;
    wire N__27306;
    wire N__27303;
    wire N__27300;
    wire N__27297;
    wire N__27294;
    wire N__27291;
    wire N__27288;
    wire N__27285;
    wire N__27282;
    wire N__27279;
    wire N__27276;
    wire N__27273;
    wire N__27270;
    wire N__27267;
    wire N__27264;
    wire N__27261;
    wire N__27258;
    wire N__27255;
    wire N__27252;
    wire N__27249;
    wire N__27246;
    wire N__27243;
    wire N__27240;
    wire N__27237;
    wire N__27234;
    wire N__27231;
    wire N__27228;
    wire N__27225;
    wire N__27222;
    wire N__27219;
    wire N__27216;
    wire N__27213;
    wire N__27210;
    wire N__27207;
    wire N__27204;
    wire N__27201;
    wire N__27198;
    wire N__27195;
    wire N__27192;
    wire N__27189;
    wire N__27186;
    wire N__27183;
    wire N__27180;
    wire N__27177;
    wire N__27174;
    wire N__27171;
    wire N__27170;
    wire N__27167;
    wire N__27166;
    wire N__27163;
    wire N__27160;
    wire N__27157;
    wire N__27154;
    wire N__27149;
    wire N__27144;
    wire N__27141;
    wire N__27140;
    wire N__27137;
    wire N__27136;
    wire N__27133;
    wire N__27130;
    wire N__27127;
    wire N__27124;
    wire N__27121;
    wire N__27118;
    wire N__27115;
    wire N__27110;
    wire N__27105;
    wire N__27104;
    wire N__27101;
    wire N__27098;
    wire N__27097;
    wire N__27094;
    wire N__27091;
    wire N__27088;
    wire N__27081;
    wire N__27078;
    wire N__27075;
    wire N__27072;
    wire N__27069;
    wire N__27066;
    wire N__27063;
    wire N__27060;
    wire N__27059;
    wire N__27056;
    wire N__27053;
    wire N__27050;
    wire N__27045;
    wire N__27044;
    wire N__27043;
    wire N__27042;
    wire N__27041;
    wire N__27040;
    wire N__27039;
    wire N__27036;
    wire N__27035;
    wire N__27032;
    wire N__27029;
    wire N__27028;
    wire N__27027;
    wire N__27026;
    wire N__27023;
    wire N__27022;
    wire N__27021;
    wire N__27020;
    wire N__27017;
    wire N__27014;
    wire N__27011;
    wire N__27010;
    wire N__27009;
    wire N__27008;
    wire N__27005;
    wire N__27000;
    wire N__26999;
    wire N__26998;
    wire N__26993;
    wire N__26990;
    wire N__26989;
    wire N__26986;
    wire N__26983;
    wire N__26976;
    wire N__26973;
    wire N__26972;
    wire N__26969;
    wire N__26966;
    wire N__26959;
    wire N__26954;
    wire N__26953;
    wire N__26950;
    wire N__26947;
    wire N__26942;
    wire N__26937;
    wire N__26934;
    wire N__26929;
    wire N__26926;
    wire N__26917;
    wire N__26912;
    wire N__26895;
    wire N__26892;
    wire N__26889;
    wire N__26886;
    wire N__26883;
    wire N__26880;
    wire N__26877;
    wire N__26874;
    wire N__26871;
    wire N__26868;
    wire N__26865;
    wire N__26862;
    wire N__26859;
    wire N__26856;
    wire N__26853;
    wire N__26850;
    wire N__26847;
    wire N__26844;
    wire N__26841;
    wire N__26838;
    wire N__26835;
    wire N__26832;
    wire N__26829;
    wire N__26826;
    wire N__26823;
    wire N__26820;
    wire N__26817;
    wire N__26814;
    wire N__26811;
    wire N__26808;
    wire N__26805;
    wire N__26802;
    wire N__26799;
    wire N__26796;
    wire N__26793;
    wire N__26790;
    wire N__26787;
    wire N__26784;
    wire N__26781;
    wire N__26778;
    wire N__26775;
    wire N__26772;
    wire N__26769;
    wire N__26766;
    wire N__26763;
    wire N__26760;
    wire N__26757;
    wire N__26754;
    wire N__26751;
    wire N__26748;
    wire N__26745;
    wire N__26744;
    wire N__26741;
    wire N__26738;
    wire N__26733;
    wire N__26730;
    wire N__26727;
    wire N__26724;
    wire N__26721;
    wire N__26718;
    wire N__26715;
    wire N__26712;
    wire N__26709;
    wire N__26708;
    wire N__26705;
    wire N__26702;
    wire N__26699;
    wire N__26696;
    wire N__26693;
    wire N__26690;
    wire N__26685;
    wire N__26684;
    wire N__26681;
    wire N__26678;
    wire N__26675;
    wire N__26670;
    wire N__26667;
    wire N__26664;
    wire N__26661;
    wire N__26658;
    wire N__26655;
    wire N__26654;
    wire N__26651;
    wire N__26650;
    wire N__26649;
    wire N__26646;
    wire N__26639;
    wire N__26634;
    wire N__26633;
    wire N__26632;
    wire N__26629;
    wire N__26624;
    wire N__26619;
    wire N__26616;
    wire N__26613;
    wire N__26610;
    wire N__26607;
    wire N__26604;
    wire N__26601;
    wire N__26598;
    wire N__26595;
    wire N__26592;
    wire N__26589;
    wire N__26586;
    wire N__26585;
    wire N__26584;
    wire N__26581;
    wire N__26578;
    wire N__26575;
    wire N__26574;
    wire N__26569;
    wire N__26566;
    wire N__26563;
    wire N__26556;
    wire N__26553;
    wire N__26550;
    wire N__26547;
    wire N__26544;
    wire N__26541;
    wire N__26538;
    wire N__26537;
    wire N__26536;
    wire N__26535;
    wire N__26532;
    wire N__26529;
    wire N__26526;
    wire N__26521;
    wire N__26514;
    wire N__26511;
    wire N__26510;
    wire N__26507;
    wire N__26504;
    wire N__26499;
    wire N__26498;
    wire N__26493;
    wire N__26490;
    wire N__26487;
    wire N__26484;
    wire N__26483;
    wire N__26482;
    wire N__26477;
    wire N__26476;
    wire N__26473;
    wire N__26470;
    wire N__26467;
    wire N__26466;
    wire N__26459;
    wire N__26456;
    wire N__26453;
    wire N__26448;
    wire N__26445;
    wire N__26444;
    wire N__26441;
    wire N__26438;
    wire N__26433;
    wire N__26430;
    wire N__26427;
    wire N__26424;
    wire N__26421;
    wire N__26418;
    wire N__26415;
    wire N__26412;
    wire N__26409;
    wire N__26406;
    wire N__26403;
    wire N__26400;
    wire N__26397;
    wire N__26396;
    wire N__26393;
    wire N__26390;
    wire N__26387;
    wire N__26384;
    wire N__26383;
    wire N__26378;
    wire N__26375;
    wire N__26372;
    wire N__26369;
    wire N__26364;
    wire N__26361;
    wire N__26358;
    wire N__26355;
    wire N__26352;
    wire N__26349;
    wire N__26346;
    wire N__26345;
    wire N__26342;
    wire N__26339;
    wire N__26336;
    wire N__26333;
    wire N__26328;
    wire N__26327;
    wire N__26324;
    wire N__26321;
    wire N__26316;
    wire N__26315;
    wire N__26312;
    wire N__26309;
    wire N__26306;
    wire N__26303;
    wire N__26300;
    wire N__26297;
    wire N__26294;
    wire N__26291;
    wire N__26286;
    wire N__26283;
    wire N__26280;
    wire N__26279;
    wire N__26276;
    wire N__26273;
    wire N__26270;
    wire N__26267;
    wire N__26264;
    wire N__26261;
    wire N__26258;
    wire N__26255;
    wire N__26250;
    wire N__26247;
    wire N__26244;
    wire N__26243;
    wire N__26240;
    wire N__26237;
    wire N__26234;
    wire N__26231;
    wire N__26228;
    wire N__26225;
    wire N__26220;
    wire N__26217;
    wire N__26214;
    wire N__26211;
    wire N__26208;
    wire N__26205;
    wire N__26202;
    wire N__26201;
    wire N__26200;
    wire N__26197;
    wire N__26194;
    wire N__26191;
    wire N__26190;
    wire N__26187;
    wire N__26184;
    wire N__26181;
    wire N__26178;
    wire N__26175;
    wire N__26172;
    wire N__26169;
    wire N__26166;
    wire N__26157;
    wire N__26154;
    wire N__26151;
    wire N__26148;
    wire N__26147;
    wire N__26144;
    wire N__26141;
    wire N__26138;
    wire N__26135;
    wire N__26132;
    wire N__26129;
    wire N__26126;
    wire N__26123;
    wire N__26118;
    wire N__26115;
    wire N__26114;
    wire N__26111;
    wire N__26108;
    wire N__26105;
    wire N__26102;
    wire N__26099;
    wire N__26096;
    wire N__26091;
    wire N__26088;
    wire N__26085;
    wire N__26082;
    wire N__26079;
    wire N__26076;
    wire N__26075;
    wire N__26070;
    wire N__26067;
    wire N__26064;
    wire N__26061;
    wire N__26058;
    wire N__26057;
    wire N__26052;
    wire N__26049;
    wire N__26048;
    wire N__26045;
    wire N__26042;
    wire N__26039;
    wire N__26036;
    wire N__26033;
    wire N__26030;
    wire N__26027;
    wire N__26022;
    wire N__26019;
    wire N__26018;
    wire N__26013;
    wire N__26010;
    wire N__26007;
    wire N__26006;
    wire N__26005;
    wire N__26002;
    wire N__25997;
    wire N__25992;
    wire N__25989;
    wire N__25986;
    wire N__25985;
    wire N__25982;
    wire N__25979;
    wire N__25976;
    wire N__25975;
    wire N__25972;
    wire N__25969;
    wire N__25966;
    wire N__25959;
    wire N__25958;
    wire N__25955;
    wire N__25952;
    wire N__25951;
    wire N__25948;
    wire N__25945;
    wire N__25942;
    wire N__25937;
    wire N__25932;
    wire N__25929;
    wire N__25928;
    wire N__25927;
    wire N__25924;
    wire N__25919;
    wire N__25914;
    wire N__25911;
    wire N__25908;
    wire N__25907;
    wire N__25906;
    wire N__25905;
    wire N__25904;
    wire N__25901;
    wire N__25892;
    wire N__25887;
    wire N__25886;
    wire N__25883;
    wire N__25880;
    wire N__25879;
    wire N__25876;
    wire N__25871;
    wire N__25866;
    wire N__25863;
    wire N__25862;
    wire N__25859;
    wire N__25856;
    wire N__25853;
    wire N__25848;
    wire N__25847;
    wire N__25844;
    wire N__25841;
    wire N__25836;
    wire N__25833;
    wire N__25830;
    wire N__25827;
    wire N__25824;
    wire N__25823;
    wire N__25820;
    wire N__25817;
    wire N__25812;
    wire N__25809;
    wire N__25808;
    wire N__25803;
    wire N__25802;
    wire N__25799;
    wire N__25796;
    wire N__25793;
    wire N__25790;
    wire N__25785;
    wire N__25782;
    wire N__25781;
    wire N__25776;
    wire N__25773;
    wire N__25770;
    wire N__25769;
    wire N__25766;
    wire N__25763;
    wire N__25760;
    wire N__25755;
    wire N__25754;
    wire N__25751;
    wire N__25748;
    wire N__25745;
    wire N__25740;
    wire N__25737;
    wire N__25734;
    wire N__25731;
    wire N__25728;
    wire N__25727;
    wire N__25724;
    wire N__25721;
    wire N__25716;
    wire N__25713;
    wire N__25710;
    wire N__25707;
    wire N__25704;
    wire N__25703;
    wire N__25700;
    wire N__25697;
    wire N__25694;
    wire N__25689;
    wire N__25688;
    wire N__25685;
    wire N__25682;
    wire N__25679;
    wire N__25674;
    wire N__25673;
    wire N__25670;
    wire N__25667;
    wire N__25664;
    wire N__25659;
    wire N__25658;
    wire N__25655;
    wire N__25652;
    wire N__25649;
    wire N__25644;
    wire N__25643;
    wire N__25640;
    wire N__25637;
    wire N__25632;
    wire N__25631;
    wire N__25628;
    wire N__25625;
    wire N__25622;
    wire N__25617;
    wire N__25616;
    wire N__25615;
    wire N__25612;
    wire N__25609;
    wire N__25606;
    wire N__25599;
    wire N__25596;
    wire N__25593;
    wire N__25590;
    wire N__25587;
    wire N__25584;
    wire N__25583;
    wire N__25582;
    wire N__25581;
    wire N__25578;
    wire N__25573;
    wire N__25570;
    wire N__25563;
    wire N__25562;
    wire N__25561;
    wire N__25556;
    wire N__25553;
    wire N__25548;
    wire N__25545;
    wire N__25542;
    wire N__25539;
    wire N__25536;
    wire N__25533;
    wire N__25530;
    wire N__25529;
    wire N__25528;
    wire N__25525;
    wire N__25524;
    wire N__25519;
    wire N__25516;
    wire N__25513;
    wire N__25506;
    wire N__25503;
    wire N__25500;
    wire N__25497;
    wire N__25494;
    wire N__25493;
    wire N__25490;
    wire N__25487;
    wire N__25484;
    wire N__25479;
    wire N__25478;
    wire N__25475;
    wire N__25472;
    wire N__25467;
    wire N__25464;
    wire N__25461;
    wire N__25458;
    wire N__25455;
    wire N__25452;
    wire N__25449;
    wire N__25446;
    wire N__25443;
    wire N__25440;
    wire N__25439;
    wire N__25436;
    wire N__25433;
    wire N__25428;
    wire N__25427;
    wire N__25426;
    wire N__25425;
    wire N__25422;
    wire N__25417;
    wire N__25414;
    wire N__25407;
    wire N__25406;
    wire N__25405;
    wire N__25404;
    wire N__25401;
    wire N__25398;
    wire N__25395;
    wire N__25392;
    wire N__25383;
    wire N__25382;
    wire N__25381;
    wire N__25380;
    wire N__25377;
    wire N__25374;
    wire N__25371;
    wire N__25368;
    wire N__25359;
    wire N__25358;
    wire N__25355;
    wire N__25354;
    wire N__25351;
    wire N__25348;
    wire N__25347;
    wire N__25346;
    wire N__25343;
    wire N__25340;
    wire N__25337;
    wire N__25334;
    wire N__25331;
    wire N__25320;
    wire N__25317;
    wire N__25316;
    wire N__25315;
    wire N__25312;
    wire N__25309;
    wire N__25308;
    wire N__25307;
    wire N__25304;
    wire N__25299;
    wire N__25296;
    wire N__25293;
    wire N__25284;
    wire N__25281;
    wire N__25278;
    wire N__25275;
    wire N__25272;
    wire N__25269;
    wire N__25268;
    wire N__25267;
    wire N__25266;
    wire N__25263;
    wire N__25256;
    wire N__25251;
    wire N__25248;
    wire N__25245;
    wire N__25242;
    wire N__25239;
    wire N__25238;
    wire N__25235;
    wire N__25232;
    wire N__25227;
    wire N__25224;
    wire N__25221;
    wire N__25218;
    wire N__25217;
    wire N__25216;
    wire N__25213;
    wire N__25210;
    wire N__25209;
    wire N__25206;
    wire N__25201;
    wire N__25198;
    wire N__25195;
    wire N__25192;
    wire N__25187;
    wire N__25182;
    wire N__25179;
    wire N__25176;
    wire N__25175;
    wire N__25174;
    wire N__25171;
    wire N__25168;
    wire N__25165;
    wire N__25160;
    wire N__25157;
    wire N__25154;
    wire N__25151;
    wire N__25146;
    wire N__25143;
    wire N__25140;
    wire N__25139;
    wire N__25138;
    wire N__25137;
    wire N__25134;
    wire N__25131;
    wire N__25128;
    wire N__25125;
    wire N__25120;
    wire N__25117;
    wire N__25114;
    wire N__25111;
    wire N__25108;
    wire N__25105;
    wire N__25098;
    wire N__25095;
    wire N__25092;
    wire N__25091;
    wire N__25090;
    wire N__25087;
    wire N__25084;
    wire N__25081;
    wire N__25076;
    wire N__25073;
    wire N__25070;
    wire N__25067;
    wire N__25062;
    wire N__25059;
    wire N__25056;
    wire N__25053;
    wire N__25050;
    wire N__25049;
    wire N__25046;
    wire N__25043;
    wire N__25042;
    wire N__25037;
    wire N__25034;
    wire N__25031;
    wire N__25028;
    wire N__25023;
    wire N__25020;
    wire N__25017;
    wire N__25014;
    wire N__25011;
    wire N__25010;
    wire N__25009;
    wire N__25006;
    wire N__25003;
    wire N__25002;
    wire N__24999;
    wire N__24994;
    wire N__24991;
    wire N__24988;
    wire N__24985;
    wire N__24982;
    wire N__24979;
    wire N__24972;
    wire N__24969;
    wire N__24966;
    wire N__24963;
    wire N__24962;
    wire N__24961;
    wire N__24958;
    wire N__24957;
    wire N__24954;
    wire N__24951;
    wire N__24950;
    wire N__24947;
    wire N__24942;
    wire N__24939;
    wire N__24936;
    wire N__24933;
    wire N__24930;
    wire N__24927;
    wire N__24922;
    wire N__24919;
    wire N__24912;
    wire N__24909;
    wire N__24906;
    wire N__24903;
    wire N__24900;
    wire N__24897;
    wire N__24894;
    wire N__24891;
    wire N__24888;
    wire N__24885;
    wire N__24882;
    wire N__24881;
    wire N__24878;
    wire N__24875;
    wire N__24870;
    wire N__24867;
    wire N__24864;
    wire N__24863;
    wire N__24862;
    wire N__24861;
    wire N__24860;
    wire N__24859;
    wire N__24858;
    wire N__24857;
    wire N__24856;
    wire N__24855;
    wire N__24854;
    wire N__24853;
    wire N__24850;
    wire N__24845;
    wire N__24838;
    wire N__24825;
    wire N__24816;
    wire N__24813;
    wire N__24810;
    wire N__24807;
    wire N__24804;
    wire N__24801;
    wire N__24798;
    wire N__24795;
    wire N__24792;
    wire N__24789;
    wire N__24786;
    wire N__24783;
    wire N__24780;
    wire N__24777;
    wire N__24774;
    wire N__24771;
    wire N__24768;
    wire N__24765;
    wire N__24762;
    wire N__24759;
    wire N__24756;
    wire N__24753;
    wire N__24750;
    wire N__24747;
    wire N__24744;
    wire N__24741;
    wire N__24738;
    wire N__24735;
    wire N__24732;
    wire N__24731;
    wire N__24730;
    wire N__24727;
    wire N__24724;
    wire N__24721;
    wire N__24718;
    wire N__24713;
    wire N__24710;
    wire N__24705;
    wire N__24702;
    wire N__24699;
    wire N__24698;
    wire N__24693;
    wire N__24690;
    wire N__24689;
    wire N__24688;
    wire N__24681;
    wire N__24678;
    wire N__24675;
    wire N__24672;
    wire N__24669;
    wire N__24666;
    wire N__24663;
    wire N__24662;
    wire N__24661;
    wire N__24660;
    wire N__24659;
    wire N__24658;
    wire N__24657;
    wire N__24654;
    wire N__24651;
    wire N__24648;
    wire N__24643;
    wire N__24638;
    wire N__24637;
    wire N__24636;
    wire N__24635;
    wire N__24634;
    wire N__24623;
    wire N__24622;
    wire N__24615;
    wire N__24614;
    wire N__24613;
    wire N__24612;
    wire N__24609;
    wire N__24608;
    wire N__24605;
    wire N__24602;
    wire N__24599;
    wire N__24596;
    wire N__24591;
    wire N__24588;
    wire N__24585;
    wire N__24580;
    wire N__24573;
    wire N__24568;
    wire N__24565;
    wire N__24560;
    wire N__24557;
    wire N__24554;
    wire N__24549;
    wire N__24548;
    wire N__24543;
    wire N__24540;
    wire N__24539;
    wire N__24536;
    wire N__24533;
    wire N__24530;
    wire N__24527;
    wire N__24524;
    wire N__24521;
    wire N__24516;
    wire N__24513;
    wire N__24510;
    wire N__24509;
    wire N__24506;
    wire N__24503;
    wire N__24500;
    wire N__24495;
    wire N__24494;
    wire N__24491;
    wire N__24488;
    wire N__24487;
    wire N__24482;
    wire N__24479;
    wire N__24474;
    wire N__24471;
    wire N__24468;
    wire N__24465;
    wire N__24462;
    wire N__24459;
    wire N__24458;
    wire N__24455;
    wire N__24452;
    wire N__24451;
    wire N__24448;
    wire N__24445;
    wire N__24442;
    wire N__24439;
    wire N__24436;
    wire N__24433;
    wire N__24430;
    wire N__24425;
    wire N__24422;
    wire N__24419;
    wire N__24418;
    wire N__24415;
    wire N__24412;
    wire N__24409;
    wire N__24402;
    wire N__24399;
    wire N__24396;
    wire N__24393;
    wire N__24390;
    wire N__24387;
    wire N__24384;
    wire N__24381;
    wire N__24378;
    wire N__24375;
    wire N__24372;
    wire N__24369;
    wire N__24368;
    wire N__24363;
    wire N__24360;
    wire N__24359;
    wire N__24354;
    wire N__24351;
    wire N__24348;
    wire N__24347;
    wire N__24344;
    wire N__24341;
    wire N__24338;
    wire N__24335;
    wire N__24332;
    wire N__24329;
    wire N__24324;
    wire N__24321;
    wire N__24318;
    wire N__24315;
    wire N__24312;
    wire N__24311;
    wire N__24308;
    wire N__24305;
    wire N__24300;
    wire N__24299;
    wire N__24298;
    wire N__24295;
    wire N__24290;
    wire N__24285;
    wire N__24282;
    wire N__24279;
    wire N__24276;
    wire N__24273;
    wire N__24270;
    wire N__24267;
    wire N__24264;
    wire N__24261;
    wire N__24260;
    wire N__24257;
    wire N__24254;
    wire N__24251;
    wire N__24248;
    wire N__24243;
    wire N__24240;
    wire N__24239;
    wire N__24236;
    wire N__24233;
    wire N__24230;
    wire N__24227;
    wire N__24224;
    wire N__24221;
    wire N__24216;
    wire N__24213;
    wire N__24210;
    wire N__24207;
    wire N__24204;
    wire N__24201;
    wire N__24198;
    wire N__24197;
    wire N__24196;
    wire N__24195;
    wire N__24192;
    wire N__24185;
    wire N__24182;
    wire N__24179;
    wire N__24176;
    wire N__24173;
    wire N__24168;
    wire N__24167;
    wire N__24166;
    wire N__24165;
    wire N__24158;
    wire N__24155;
    wire N__24152;
    wire N__24147;
    wire N__24144;
    wire N__24141;
    wire N__24138;
    wire N__24135;
    wire N__24132;
    wire N__24129;
    wire N__24128;
    wire N__24125;
    wire N__24122;
    wire N__24119;
    wire N__24116;
    wire N__24113;
    wire N__24110;
    wire N__24107;
    wire N__24102;
    wire N__24101;
    wire N__24100;
    wire N__24099;
    wire N__24096;
    wire N__24089;
    wire N__24086;
    wire N__24083;
    wire N__24080;
    wire N__24077;
    wire N__24072;
    wire N__24071;
    wire N__24066;
    wire N__24063;
    wire N__24062;
    wire N__24057;
    wire N__24054;
    wire N__24051;
    wire N__24048;
    wire N__24045;
    wire N__24042;
    wire N__24039;
    wire N__24036;
    wire N__24033;
    wire N__24030;
    wire N__24027;
    wire N__24024;
    wire N__24021;
    wire N__24018;
    wire N__24015;
    wire N__24012;
    wire N__24009;
    wire N__24006;
    wire N__24003;
    wire N__24000;
    wire N__23997;
    wire N__23994;
    wire N__23991;
    wire N__23990;
    wire N__23987;
    wire N__23984;
    wire N__23979;
    wire N__23976;
    wire N__23975;
    wire N__23974;
    wire N__23973;
    wire N__23972;
    wire N__23969;
    wire N__23966;
    wire N__23961;
    wire N__23958;
    wire N__23953;
    wire N__23950;
    wire N__23943;
    wire N__23942;
    wire N__23941;
    wire N__23936;
    wire N__23933;
    wire N__23930;
    wire N__23925;
    wire N__23922;
    wire N__23921;
    wire N__23920;
    wire N__23917;
    wire N__23912;
    wire N__23907;
    wire N__23904;
    wire N__23901;
    wire N__23898;
    wire N__23895;
    wire N__23892;
    wire N__23891;
    wire N__23888;
    wire N__23885;
    wire N__23882;
    wire N__23877;
    wire N__23874;
    wire N__23871;
    wire N__23868;
    wire N__23865;
    wire N__23864;
    wire N__23861;
    wire N__23858;
    wire N__23855;
    wire N__23850;
    wire N__23847;
    wire N__23844;
    wire N__23841;
    wire N__23838;
    wire N__23835;
    wire N__23832;
    wire N__23831;
    wire N__23830;
    wire N__23829;
    wire N__23826;
    wire N__23819;
    wire N__23814;
    wire N__23813;
    wire N__23812;
    wire N__23807;
    wire N__23804;
    wire N__23799;
    wire N__23796;
    wire N__23793;
    wire N__23790;
    wire N__23787;
    wire N__23784;
    wire N__23781;
    wire N__23778;
    wire N__23777;
    wire N__23776;
    wire N__23773;
    wire N__23770;
    wire N__23765;
    wire N__23762;
    wire N__23757;
    wire N__23754;
    wire N__23753;
    wire N__23750;
    wire N__23747;
    wire N__23744;
    wire N__23739;
    wire N__23736;
    wire N__23733;
    wire N__23730;
    wire N__23727;
    wire N__23724;
    wire N__23721;
    wire N__23718;
    wire N__23717;
    wire N__23712;
    wire N__23709;
    wire N__23708;
    wire N__23705;
    wire N__23702;
    wire N__23701;
    wire N__23698;
    wire N__23695;
    wire N__23692;
    wire N__23687;
    wire N__23682;
    wire N__23679;
    wire N__23678;
    wire N__23675;
    wire N__23672;
    wire N__23667;
    wire N__23664;
    wire N__23663;
    wire N__23660;
    wire N__23657;
    wire N__23652;
    wire N__23649;
    wire N__23648;
    wire N__23647;
    wire N__23644;
    wire N__23639;
    wire N__23634;
    wire N__23631;
    wire N__23630;
    wire N__23629;
    wire N__23626;
    wire N__23623;
    wire N__23620;
    wire N__23615;
    wire N__23610;
    wire N__23607;
    wire N__23606;
    wire N__23605;
    wire N__23602;
    wire N__23599;
    wire N__23594;
    wire N__23589;
    wire N__23586;
    wire N__23583;
    wire N__23580;
    wire N__23577;
    wire N__23574;
    wire N__23571;
    wire N__23568;
    wire N__23565;
    wire N__23564;
    wire N__23561;
    wire N__23558;
    wire N__23555;
    wire N__23552;
    wire N__23547;
    wire N__23544;
    wire N__23541;
    wire N__23538;
    wire N__23535;
    wire N__23532;
    wire N__23529;
    wire N__23526;
    wire N__23523;
    wire N__23520;
    wire N__23517;
    wire N__23514;
    wire N__23513;
    wire N__23512;
    wire N__23509;
    wire N__23504;
    wire N__23499;
    wire N__23496;
    wire N__23495;
    wire N__23494;
    wire N__23491;
    wire N__23486;
    wire N__23481;
    wire N__23478;
    wire N__23477;
    wire N__23476;
    wire N__23473;
    wire N__23470;
    wire N__23467;
    wire N__23460;
    wire N__23457;
    wire N__23456;
    wire N__23455;
    wire N__23452;
    wire N__23449;
    wire N__23446;
    wire N__23439;
    wire N__23436;
    wire N__23433;
    wire N__23430;
    wire N__23427;
    wire N__23424;
    wire N__23421;
    wire N__23418;
    wire N__23415;
    wire N__23412;
    wire N__23409;
    wire N__23406;
    wire N__23403;
    wire N__23400;
    wire N__23397;
    wire N__23394;
    wire N__23391;
    wire N__23388;
    wire N__23385;
    wire N__23382;
    wire N__23379;
    wire N__23376;
    wire N__23373;
    wire N__23370;
    wire N__23367;
    wire N__23364;
    wire N__23363;
    wire N__23360;
    wire N__23357;
    wire N__23354;
    wire N__23349;
    wire N__23346;
    wire N__23343;
    wire N__23340;
    wire N__23337;
    wire N__23334;
    wire N__23331;
    wire N__23330;
    wire N__23325;
    wire N__23322;
    wire N__23321;
    wire N__23320;
    wire N__23313;
    wire N__23310;
    wire N__23307;
    wire N__23304;
    wire N__23301;
    wire N__23298;
    wire N__23295;
    wire N__23292;
    wire N__23291;
    wire N__23288;
    wire N__23285;
    wire N__23282;
    wire N__23277;
    wire N__23276;
    wire N__23271;
    wire N__23268;
    wire N__23265;
    wire N__23262;
    wire N__23259;
    wire N__23256;
    wire N__23253;
    wire N__23250;
    wire N__23247;
    wire N__23244;
    wire N__23243;
    wire N__23240;
    wire N__23237;
    wire N__23234;
    wire N__23229;
    wire N__23226;
    wire N__23223;
    wire N__23220;
    wire N__23217;
    wire N__23214;
    wire N__23211;
    wire N__23208;
    wire N__23205;
    wire N__23202;
    wire N__23199;
    wire N__23196;
    wire N__23195;
    wire N__23192;
    wire N__23189;
    wire N__23184;
    wire N__23181;
    wire N__23178;
    wire N__23175;
    wire N__23174;
    wire N__23171;
    wire N__23168;
    wire N__23163;
    wire N__23160;
    wire N__23157;
    wire N__23154;
    wire N__23153;
    wire N__23150;
    wire N__23147;
    wire N__23144;
    wire N__23139;
    wire N__23138;
    wire N__23133;
    wire N__23132;
    wire N__23129;
    wire N__23126;
    wire N__23123;
    wire N__23120;
    wire N__23117;
    wire N__23114;
    wire N__23111;
    wire N__23108;
    wire N__23103;
    wire N__23100;
    wire N__23097;
    wire N__23094;
    wire N__23093;
    wire N__23090;
    wire N__23087;
    wire N__23082;
    wire N__23081;
    wire N__23078;
    wire N__23075;
    wire N__23072;
    wire N__23069;
    wire N__23066;
    wire N__23063;
    wire N__23060;
    wire N__23057;
    wire N__23052;
    wire N__23049;
    wire N__23046;
    wire N__23045;
    wire N__23042;
    wire N__23039;
    wire N__23034;
    wire N__23031;
    wire N__23028;
    wire N__23027;
    wire N__23022;
    wire N__23019;
    wire N__23016;
    wire N__23013;
    wire N__23010;
    wire N__23007;
    wire N__23004;
    wire N__23001;
    wire N__22998;
    wire N__22997;
    wire N__22994;
    wire N__22991;
    wire N__22988;
    wire N__22983;
    wire N__22980;
    wire N__22977;
    wire N__22974;
    wire N__22971;
    wire N__22970;
    wire N__22967;
    wire N__22964;
    wire N__22959;
    wire N__22956;
    wire N__22953;
    wire N__22950;
    wire N__22947;
    wire N__22946;
    wire N__22943;
    wire N__22940;
    wire N__22937;
    wire N__22932;
    wire N__22931;
    wire N__22930;
    wire N__22927;
    wire N__22922;
    wire N__22919;
    wire N__22916;
    wire N__22913;
    wire N__22910;
    wire N__22907;
    wire N__22902;
    wire N__22901;
    wire N__22898;
    wire N__22895;
    wire N__22892;
    wire N__22887;
    wire N__22886;
    wire N__22881;
    wire N__22878;
    wire N__22875;
    wire N__22872;
    wire N__22869;
    wire N__22866;
    wire N__22863;
    wire N__22862;
    wire N__22857;
    wire N__22854;
    wire N__22853;
    wire N__22852;
    wire N__22845;
    wire N__22842;
    wire N__22839;
    wire N__22836;
    wire N__22833;
    wire N__22830;
    wire N__22827;
    wire N__22824;
    wire N__22823;
    wire N__22818;
    wire N__22815;
    wire N__22812;
    wire N__22809;
    wire N__22808;
    wire N__22805;
    wire N__22802;
    wire N__22799;
    wire N__22796;
    wire N__22793;
    wire N__22790;
    wire N__22785;
    wire N__22782;
    wire N__22779;
    wire N__22776;
    wire N__22773;
    wire N__22772;
    wire N__22769;
    wire N__22766;
    wire N__22763;
    wire N__22760;
    wire N__22755;
    wire N__22752;
    wire N__22749;
    wire N__22746;
    wire N__22743;
    wire N__22740;
    wire N__22739;
    wire N__22736;
    wire N__22733;
    wire N__22730;
    wire N__22727;
    wire N__22724;
    wire N__22719;
    wire N__22716;
    wire N__22715;
    wire N__22710;
    wire N__22707;
    wire N__22704;
    wire N__22701;
    wire N__22698;
    wire N__22695;
    wire N__22692;
    wire N__22691;
    wire N__22688;
    wire N__22685;
    wire N__22682;
    wire N__22677;
    wire N__22674;
    wire N__22671;
    wire N__22668;
    wire N__22665;
    wire N__22662;
    wire N__22659;
    wire N__22656;
    wire N__22653;
    wire N__22650;
    wire N__22649;
    wire N__22648;
    wire N__22647;
    wire N__22644;
    wire N__22641;
    wire N__22636;
    wire N__22629;
    wire N__22626;
    wire N__22623;
    wire N__22620;
    wire N__22617;
    wire N__22614;
    wire N__22611;
    wire N__22608;
    wire N__22605;
    wire N__22602;
    wire N__22599;
    wire N__22596;
    wire N__22593;
    wire N__22590;
    wire N__22587;
    wire N__22584;
    wire N__22581;
    wire N__22578;
    wire N__22575;
    wire N__22572;
    wire N__22569;
    wire N__22566;
    wire N__22565;
    wire N__22562;
    wire N__22559;
    wire N__22556;
    wire N__22553;
    wire N__22548;
    wire N__22545;
    wire N__22544;
    wire N__22539;
    wire N__22536;
    wire N__22533;
    wire N__22532;
    wire N__22531;
    wire N__22530;
    wire N__22529;
    wire N__22522;
    wire N__22517;
    wire N__22516;
    wire N__22515;
    wire N__22514;
    wire N__22509;
    wire N__22502;
    wire N__22497;
    wire N__22494;
    wire N__22493;
    wire N__22492;
    wire N__22485;
    wire N__22482;
    wire N__22481;
    wire N__22478;
    wire N__22475;
    wire N__22474;
    wire N__22473;
    wire N__22472;
    wire N__22467;
    wire N__22464;
    wire N__22461;
    wire N__22458;
    wire N__22451;
    wire N__22448;
    wire N__22443;
    wire N__22440;
    wire N__22437;
    wire N__22434;
    wire N__22431;
    wire N__22428;
    wire N__22425;
    wire N__22422;
    wire N__22419;
    wire N__22416;
    wire N__22413;
    wire N__22412;
    wire N__22407;
    wire N__22404;
    wire N__22401;
    wire N__22398;
    wire N__22395;
    wire N__22392;
    wire N__22391;
    wire N__22390;
    wire N__22389;
    wire N__22386;
    wire N__22383;
    wire N__22378;
    wire N__22371;
    wire N__22368;
    wire N__22367;
    wire N__22366;
    wire N__22363;
    wire N__22358;
    wire N__22353;
    wire N__22350;
    wire N__22347;
    wire N__22344;
    wire N__22341;
    wire N__22338;
    wire N__22335;
    wire N__22332;
    wire N__22329;
    wire N__22326;
    wire N__22323;
    wire N__22322;
    wire N__22319;
    wire N__22316;
    wire N__22313;
    wire N__22310;
    wire N__22307;
    wire N__22304;
    wire N__22299;
    wire N__22296;
    wire N__22293;
    wire N__22290;
    wire N__22287;
    wire N__22284;
    wire N__22281;
    wire N__22278;
    wire N__22275;
    wire N__22272;
    wire N__22269;
    wire N__22266;
    wire N__22263;
    wire N__22260;
    wire N__22257;
    wire N__22254;
    wire N__22251;
    wire N__22248;
    wire N__22247;
    wire N__22244;
    wire N__22243;
    wire N__22240;
    wire N__22237;
    wire N__22234;
    wire N__22231;
    wire N__22228;
    wire N__22225;
    wire N__22222;
    wire N__22217;
    wire N__22214;
    wire N__22209;
    wire N__22206;
    wire N__22203;
    wire N__22200;
    wire N__22197;
    wire N__22196;
    wire N__22193;
    wire N__22190;
    wire N__22189;
    wire N__22186;
    wire N__22183;
    wire N__22180;
    wire N__22177;
    wire N__22174;
    wire N__22171;
    wire N__22166;
    wire N__22163;
    wire N__22158;
    wire N__22155;
    wire N__22152;
    wire N__22149;
    wire N__22146;
    wire N__22143;
    wire N__22140;
    wire N__22139;
    wire N__22136;
    wire N__22133;
    wire N__22132;
    wire N__22129;
    wire N__22126;
    wire N__22123;
    wire N__22120;
    wire N__22117;
    wire N__22114;
    wire N__22109;
    wire N__22106;
    wire N__22101;
    wire N__22098;
    wire N__22095;
    wire N__22092;
    wire N__22089;
    wire N__22086;
    wire N__22083;
    wire N__22080;
    wire N__22077;
    wire N__22074;
    wire N__22071;
    wire N__22068;
    wire N__22065;
    wire N__22062;
    wire N__22059;
    wire N__22056;
    wire N__22053;
    wire N__22052;
    wire N__22051;
    wire N__22048;
    wire N__22047;
    wire N__22044;
    wire N__22041;
    wire N__22038;
    wire N__22035;
    wire N__22030;
    wire N__22023;
    wire N__22022;
    wire N__22019;
    wire N__22016;
    wire N__22015;
    wire N__22010;
    wire N__22009;
    wire N__22008;
    wire N__22005;
    wire N__22002;
    wire N__21997;
    wire N__21990;
    wire N__21987;
    wire N__21984;
    wire N__21981;
    wire N__21978;
    wire N__21977;
    wire N__21974;
    wire N__21971;
    wire N__21968;
    wire N__21963;
    wire N__21960;
    wire N__21957;
    wire N__21954;
    wire N__21953;
    wire N__21950;
    wire N__21947;
    wire N__21946;
    wire N__21943;
    wire N__21940;
    wire N__21937;
    wire N__21934;
    wire N__21931;
    wire N__21928;
    wire N__21923;
    wire N__21920;
    wire N__21915;
    wire N__21912;
    wire N__21909;
    wire N__21908;
    wire N__21905;
    wire N__21902;
    wire N__21899;
    wire N__21896;
    wire N__21891;
    wire N__21890;
    wire N__21889;
    wire N__21886;
    wire N__21883;
    wire N__21880;
    wire N__21877;
    wire N__21874;
    wire N__21871;
    wire N__21868;
    wire N__21865;
    wire N__21860;
    wire N__21857;
    wire N__21852;
    wire N__21849;
    wire N__21848;
    wire N__21845;
    wire N__21842;
    wire N__21837;
    wire N__21834;
    wire N__21831;
    wire N__21830;
    wire N__21827;
    wire N__21824;
    wire N__21821;
    wire N__21820;
    wire N__21817;
    wire N__21814;
    wire N__21811;
    wire N__21808;
    wire N__21805;
    wire N__21802;
    wire N__21799;
    wire N__21796;
    wire N__21793;
    wire N__21786;
    wire N__21783;
    wire N__21780;
    wire N__21777;
    wire N__21774;
    wire N__21771;
    wire N__21770;
    wire N__21767;
    wire N__21764;
    wire N__21763;
    wire N__21760;
    wire N__21757;
    wire N__21754;
    wire N__21751;
    wire N__21748;
    wire N__21745;
    wire N__21740;
    wire N__21737;
    wire N__21732;
    wire N__21729;
    wire N__21726;
    wire N__21723;
    wire N__21720;
    wire N__21717;
    wire N__21716;
    wire N__21713;
    wire N__21710;
    wire N__21709;
    wire N__21706;
    wire N__21703;
    wire N__21700;
    wire N__21697;
    wire N__21694;
    wire N__21691;
    wire N__21686;
    wire N__21683;
    wire N__21678;
    wire N__21675;
    wire N__21672;
    wire N__21669;
    wire N__21668;
    wire N__21665;
    wire N__21664;
    wire N__21661;
    wire N__21658;
    wire N__21655;
    wire N__21652;
    wire N__21647;
    wire N__21644;
    wire N__21641;
    wire N__21638;
    wire N__21635;
    wire N__21630;
    wire N__21627;
    wire N__21624;
    wire N__21621;
    wire N__21620;
    wire N__21617;
    wire N__21616;
    wire N__21613;
    wire N__21610;
    wire N__21607;
    wire N__21604;
    wire N__21601;
    wire N__21598;
    wire N__21595;
    wire N__21590;
    wire N__21587;
    wire N__21582;
    wire N__21579;
    wire N__21576;
    wire N__21573;
    wire N__21570;
    wire N__21569;
    wire N__21566;
    wire N__21563;
    wire N__21562;
    wire N__21559;
    wire N__21556;
    wire N__21553;
    wire N__21550;
    wire N__21547;
    wire N__21544;
    wire N__21541;
    wire N__21536;
    wire N__21531;
    wire N__21528;
    wire N__21525;
    wire N__21524;
    wire N__21523;
    wire N__21516;
    wire N__21513;
    wire N__21510;
    wire N__21507;
    wire N__21504;
    wire N__21501;
    wire N__21498;
    wire N__21495;
    wire N__21494;
    wire N__21489;
    wire N__21486;
    wire N__21485;
    wire N__21482;
    wire N__21479;
    wire N__21476;
    wire N__21473;
    wire N__21472;
    wire N__21469;
    wire N__21466;
    wire N__21463;
    wire N__21460;
    wire N__21455;
    wire N__21452;
    wire N__21449;
    wire N__21446;
    wire N__21443;
    wire N__21438;
    wire N__21435;
    wire N__21434;
    wire N__21431;
    wire N__21430;
    wire N__21427;
    wire N__21424;
    wire N__21421;
    wire N__21418;
    wire N__21415;
    wire N__21412;
    wire N__21409;
    wire N__21404;
    wire N__21401;
    wire N__21398;
    wire N__21393;
    wire N__21390;
    wire N__21387;
    wire N__21384;
    wire N__21383;
    wire N__21380;
    wire N__21379;
    wire N__21376;
    wire N__21373;
    wire N__21370;
    wire N__21367;
    wire N__21364;
    wire N__21361;
    wire N__21358;
    wire N__21355;
    wire N__21352;
    wire N__21349;
    wire N__21342;
    wire N__21339;
    wire N__21336;
    wire N__21333;
    wire N__21330;
    wire N__21329;
    wire N__21326;
    wire N__21323;
    wire N__21322;
    wire N__21319;
    wire N__21316;
    wire N__21313;
    wire N__21310;
    wire N__21307;
    wire N__21304;
    wire N__21299;
    wire N__21296;
    wire N__21291;
    wire N__21288;
    wire N__21285;
    wire N__21282;
    wire N__21279;
    wire N__21276;
    wire N__21273;
    wire N__21270;
    wire N__21267;
    wire N__21264;
    wire N__21261;
    wire N__21260;
    wire N__21257;
    wire N__21254;
    wire N__21249;
    wire N__21246;
    wire N__21243;
    wire N__21240;
    wire N__21237;
    wire N__21234;
    wire N__21231;
    wire N__21228;
    wire N__21227;
    wire N__21224;
    wire N__21221;
    wire N__21218;
    wire N__21215;
    wire N__21212;
    wire N__21207;
    wire N__21204;
    wire N__21201;
    wire N__21198;
    wire N__21195;
    wire N__21192;
    wire N__21189;
    wire N__21186;
    wire N__21183;
    wire N__21180;
    wire N__21177;
    wire N__21174;
    wire N__21171;
    wire N__21168;
    wire N__21165;
    wire N__21162;
    wire N__21159;
    wire N__21156;
    wire N__21153;
    wire N__21150;
    wire N__21147;
    wire N__21144;
    wire N__21141;
    wire N__21138;
    wire N__21135;
    wire N__21132;
    wire N__21129;
    wire N__21126;
    wire N__21123;
    wire N__21120;
    wire N__21119;
    wire N__21116;
    wire N__21113;
    wire N__21110;
    wire N__21105;
    wire N__21102;
    wire N__21099;
    wire N__21096;
    wire N__21093;
    wire N__21090;
    wire N__21087;
    wire N__21086;
    wire N__21083;
    wire N__21080;
    wire N__21077;
    wire N__21074;
    wire N__21071;
    wire N__21066;
    wire N__21063;
    wire N__21060;
    wire N__21057;
    wire N__21054;
    wire N__21051;
    wire N__21048;
    wire N__21047;
    wire N__21044;
    wire N__21041;
    wire N__21038;
    wire N__21035;
    wire N__21032;
    wire N__21027;
    wire N__21024;
    wire N__21021;
    wire N__21018;
    wire N__21015;
    wire N__21012;
    wire N__21011;
    wire N__21008;
    wire N__21005;
    wire N__21002;
    wire N__20999;
    wire N__20996;
    wire N__20991;
    wire N__20988;
    wire N__20985;
    wire N__20982;
    wire N__20979;
    wire N__20976;
    wire N__20973;
    wire N__20970;
    wire N__20967;
    wire N__20966;
    wire N__20963;
    wire N__20960;
    wire N__20957;
    wire N__20952;
    wire N__20949;
    wire N__20946;
    wire N__20943;
    wire N__20940;
    wire N__20937;
    wire N__20934;
    wire N__20931;
    wire N__20930;
    wire N__20927;
    wire N__20924;
    wire N__20921;
    wire N__20918;
    wire N__20915;
    wire N__20910;
    wire N__20907;
    wire N__20904;
    wire N__20901;
    wire N__20898;
    wire N__20895;
    wire N__20892;
    wire N__20889;
    wire N__20888;
    wire N__20885;
    wire N__20882;
    wire N__20879;
    wire N__20876;
    wire N__20873;
    wire N__20868;
    wire N__20865;
    wire N__20862;
    wire N__20859;
    wire N__20856;
    wire N__20853;
    wire N__20850;
    wire N__20847;
    wire N__20844;
    wire N__20841;
    wire N__20838;
    wire N__20835;
    wire N__20832;
    wire N__20829;
    wire N__20826;
    wire N__20823;
    wire N__20820;
    wire N__20817;
    wire N__20814;
    wire N__20811;
    wire N__20808;
    wire N__20805;
    wire N__20802;
    wire N__20799;
    wire N__20796;
    wire N__20793;
    wire N__20790;
    wire N__20787;
    wire N__20784;
    wire N__20783;
    wire N__20782;
    wire N__20779;
    wire N__20778;
    wire N__20777;
    wire N__20774;
    wire N__20771;
    wire N__20768;
    wire N__20765;
    wire N__20762;
    wire N__20757;
    wire N__20754;
    wire N__20749;
    wire N__20746;
    wire N__20739;
    wire N__20738;
    wire N__20735;
    wire N__20734;
    wire N__20731;
    wire N__20728;
    wire N__20725;
    wire N__20724;
    wire N__20723;
    wire N__20722;
    wire N__20719;
    wire N__20714;
    wire N__20711;
    wire N__20708;
    wire N__20705;
    wire N__20702;
    wire N__20699;
    wire N__20694;
    wire N__20691;
    wire N__20682;
    wire N__20681;
    wire N__20678;
    wire N__20677;
    wire N__20674;
    wire N__20671;
    wire N__20668;
    wire N__20665;
    wire N__20658;
    wire N__20655;
    wire N__20652;
    wire N__20649;
    wire N__20646;
    wire N__20643;
    wire N__20642;
    wire N__20639;
    wire N__20636;
    wire N__20631;
    wire N__20628;
    wire N__20625;
    wire N__20622;
    wire N__20619;
    wire N__20616;
    wire N__20613;
    wire N__20610;
    wire N__20607;
    wire N__20604;
    wire N__20601;
    wire N__20598;
    wire N__20595;
    wire N__20592;
    wire N__20589;
    wire N__20586;
    wire N__20583;
    wire N__20580;
    wire N__20577;
    wire N__20574;
    wire N__20571;
    wire N__20568;
    wire N__20565;
    wire N__20562;
    wire N__20559;
    wire N__20556;
    wire N__20555;
    wire N__20552;
    wire N__20549;
    wire N__20546;
    wire N__20541;
    wire N__20538;
    wire N__20535;
    wire N__20532;
    wire N__20531;
    wire N__20528;
    wire N__20527;
    wire N__20524;
    wire N__20523;
    wire N__20520;
    wire N__20515;
    wire N__20512;
    wire N__20507;
    wire N__20502;
    wire N__20499;
    wire N__20496;
    wire N__20495;
    wire N__20494;
    wire N__20491;
    wire N__20488;
    wire N__20485;
    wire N__20480;
    wire N__20475;
    wire N__20472;
    wire N__20469;
    wire N__20466;
    wire N__20465;
    wire N__20462;
    wire N__20459;
    wire N__20458;
    wire N__20455;
    wire N__20452;
    wire N__20449;
    wire N__20444;
    wire N__20439;
    wire N__20438;
    wire N__20435;
    wire N__20430;
    wire N__20427;
    wire N__20424;
    wire N__20423;
    wire N__20418;
    wire N__20415;
    wire N__20412;
    wire N__20409;
    wire N__20406;
    wire N__20403;
    wire N__20402;
    wire N__20399;
    wire N__20396;
    wire N__20393;
    wire N__20388;
    wire N__20385;
    wire N__20382;
    wire N__20381;
    wire N__20378;
    wire N__20375;
    wire N__20372;
    wire N__20367;
    wire N__20364;
    wire N__20361;
    wire N__20360;
    wire N__20357;
    wire N__20354;
    wire N__20351;
    wire N__20346;
    wire N__20343;
    wire N__20340;
    wire N__20339;
    wire N__20336;
    wire N__20333;
    wire N__20330;
    wire N__20325;
    wire N__20322;
    wire N__20321;
    wire N__20318;
    wire N__20315;
    wire N__20312;
    wire N__20307;
    wire N__20304;
    wire N__20301;
    wire N__20300;
    wire N__20297;
    wire N__20294;
    wire N__20291;
    wire N__20286;
    wire N__20283;
    wire N__20282;
    wire N__20279;
    wire N__20276;
    wire N__20273;
    wire N__20268;
    wire N__20265;
    wire N__20264;
    wire N__20263;
    wire N__20258;
    wire N__20255;
    wire N__20252;
    wire N__20247;
    wire N__20244;
    wire N__20243;
    wire N__20242;
    wire N__20237;
    wire N__20234;
    wire N__20231;
    wire N__20226;
    wire N__20223;
    wire N__20220;
    wire N__20217;
    wire N__20214;
    wire N__20211;
    wire N__20208;
    wire N__20207;
    wire N__20206;
    wire N__20203;
    wire N__20198;
    wire N__20193;
    wire N__20190;
    wire N__20187;
    wire N__20186;
    wire N__20183;
    wire N__20180;
    wire N__20175;
    wire N__20172;
    wire N__20169;
    wire N__20166;
    wire N__20163;
    wire N__20160;
    wire N__20159;
    wire N__20156;
    wire N__20153;
    wire N__20150;
    wire N__20145;
    wire N__20142;
    wire N__20139;
    wire N__20136;
    wire N__20133;
    wire N__20130;
    wire N__20127;
    wire N__20124;
    wire N__20121;
    wire N__20118;
    wire N__20115;
    wire N__20112;
    wire N__20109;
    wire N__20106;
    wire N__20103;
    wire N__20102;
    wire N__20097;
    wire N__20094;
    wire N__20093;
    wire N__20088;
    wire N__20085;
    wire N__20082;
    wire N__20079;
    wire N__20076;
    wire N__20073;
    wire N__20072;
    wire N__20071;
    wire N__20064;
    wire N__20061;
    wire N__20058;
    wire N__20055;
    wire N__20052;
    wire N__20049;
    wire N__20048;
    wire N__20043;
    wire N__20040;
    wire N__20039;
    wire N__20034;
    wire N__20031;
    wire N__20028;
    wire N__20025;
    wire N__20022;
    wire N__20019;
    wire N__20016;
    wire N__20015;
    wire N__20012;
    wire N__20009;
    wire N__20004;
    wire N__20003;
    wire N__19998;
    wire N__19997;
    wire N__19994;
    wire N__19991;
    wire N__19986;
    wire N__19983;
    wire N__19980;
    wire N__19977;
    wire N__19974;
    wire N__19973;
    wire N__19968;
    wire N__19965;
    wire N__19962;
    wire N__19959;
    wire N__19958;
    wire N__19953;
    wire N__19950;
    wire N__19949;
    wire N__19948;
    wire N__19941;
    wire N__19938;
    wire N__19935;
    wire N__19932;
    wire N__19929;
    wire N__19928;
    wire N__19925;
    wire N__19922;
    wire N__19919;
    wire N__19916;
    wire N__19913;
    wire N__19910;
    wire N__19905;
    wire N__19904;
    wire N__19903;
    wire N__19898;
    wire N__19895;
    wire N__19890;
    wire N__19887;
    wire N__19884;
    wire N__19881;
    wire N__19880;
    wire N__19877;
    wire N__19874;
    wire N__19869;
    wire N__19868;
    wire N__19863;
    wire N__19860;
    wire N__19857;
    wire N__19854;
    wire N__19851;
    wire N__19850;
    wire N__19847;
    wire N__19844;
    wire N__19839;
    wire N__19838;
    wire N__19835;
    wire N__19832;
    wire N__19827;
    wire N__19824;
    wire N__19821;
    wire N__19818;
    wire N__19817;
    wire N__19816;
    wire N__19813;
    wire N__19810;
    wire N__19807;
    wire N__19800;
    wire N__19797;
    wire N__19794;
    wire N__19791;
    wire N__19788;
    wire N__19785;
    wire N__19784;
    wire N__19779;
    wire N__19776;
    wire N__19773;
    wire N__19770;
    wire N__19767;
    wire N__19764;
    wire N__19763;
    wire N__19758;
    wire N__19755;
    wire N__19754;
    wire N__19753;
    wire N__19746;
    wire N__19743;
    wire N__19740;
    wire N__19737;
    wire N__19734;
    wire N__19731;
    wire N__19728;
    wire N__19725;
    wire N__19722;
    wire N__19719;
    wire N__19716;
    wire N__19713;
    wire N__19710;
    wire N__19707;
    wire N__19704;
    wire N__19703;
    wire N__19698;
    wire N__19695;
    wire N__19692;
    wire N__19689;
    wire N__19686;
    wire N__19683;
    wire N__19682;
    wire N__19677;
    wire N__19674;
    wire N__19673;
    wire N__19672;
    wire N__19665;
    wire N__19664;
    wire N__19661;
    wire N__19658;
    wire N__19655;
    wire N__19652;
    wire N__19649;
    wire N__19644;
    wire N__19641;
    wire N__19638;
    wire N__19637;
    wire N__19632;
    wire N__19629;
    wire N__19626;
    wire N__19623;
    wire N__19620;
    wire N__19617;
    wire N__19614;
    wire N__19613;
    wire N__19610;
    wire N__19607;
    wire N__19602;
    wire N__19599;
    wire N__19596;
    wire N__19593;
    wire N__19592;
    wire N__19587;
    wire N__19584;
    wire N__19581;
    wire N__19578;
    wire N__19575;
    wire N__19572;
    wire N__19569;
    wire N__19566;
    wire N__19563;
    wire N__19560;
    wire N__19557;
    wire N__19554;
    wire N__19551;
    wire N__19548;
    wire N__19547;
    wire N__19542;
    wire N__19539;
    wire N__19536;
    wire N__19533;
    wire N__19532;
    wire N__19527;
    wire N__19524;
    wire N__19523;
    wire N__19522;
    wire N__19515;
    wire N__19512;
    wire N__19509;
    wire N__19506;
    wire N__19503;
    wire N__19500;
    wire N__19499;
    wire N__19498;
    wire N__19495;
    wire N__19490;
    wire N__19485;
    wire N__19482;
    wire N__19479;
    wire N__19476;
    wire N__19475;
    wire N__19472;
    wire N__19469;
    wire N__19464;
    wire N__19461;
    wire N__19458;
    wire N__19455;
    wire N__19452;
    wire N__19451;
    wire N__19446;
    wire N__19443;
    wire N__19440;
    wire N__19437;
    wire N__19434;
    wire N__19431;
    wire N__19430;
    wire N__19429;
    wire N__19422;
    wire N__19419;
    wire N__19416;
    wire N__19413;
    wire N__19410;
    wire N__19407;
    wire N__19404;
    wire N__19403;
    wire N__19398;
    wire N__19395;
    wire N__19392;
    wire N__19389;
    wire N__19388;
    wire N__19383;
    wire N__19380;
    wire N__19377;
    wire N__19374;
    wire N__19371;
    wire N__19370;
    wire N__19367;
    wire N__19364;
    wire N__19359;
    wire N__19356;
    wire N__19353;
    wire N__19350;
    wire N__19347;
    wire N__19344;
    wire N__19341;
    wire N__19338;
    wire N__19335;
    wire N__19332;
    wire N__19329;
    wire N__19326;
    wire N__19325;
    wire N__19324;
    wire N__19321;
    wire N__19318;
    wire N__19317;
    wire N__19314;
    wire N__19313;
    wire N__19308;
    wire N__19305;
    wire N__19300;
    wire N__19293;
    wire N__19292;
    wire N__19289;
    wire N__19286;
    wire N__19285;
    wire N__19284;
    wire N__19283;
    wire N__19278;
    wire N__19275;
    wire N__19270;
    wire N__19267;
    wire N__19262;
    wire N__19257;
    wire N__19256;
    wire N__19253;
    wire N__19250;
    wire N__19249;
    wire N__19248;
    wire N__19247;
    wire N__19242;
    wire N__19241;
    wire N__19238;
    wire N__19233;
    wire N__19230;
    wire N__19227;
    wire N__19222;
    wire N__19215;
    wire N__19212;
    wire N__19209;
    wire N__19206;
    wire N__19203;
    wire N__19200;
    wire N__19199;
    wire N__19198;
    wire N__19193;
    wire N__19190;
    wire N__19187;
    wire N__19184;
    wire N__19181;
    wire N__19176;
    wire N__19175;
    wire N__19174;
    wire N__19169;
    wire N__19166;
    wire N__19163;
    wire N__19158;
    wire N__19157;
    wire N__19156;
    wire N__19155;
    wire N__19152;
    wire N__19149;
    wire N__19144;
    wire N__19141;
    wire N__19138;
    wire N__19135;
    wire N__19130;
    wire N__19127;
    wire N__19122;
    wire N__19119;
    wire N__19116;
    wire N__19115;
    wire N__19110;
    wire N__19107;
    wire N__19104;
    wire N__19101;
    wire N__19100;
    wire N__19097;
    wire N__19094;
    wire N__19089;
    wire N__19088;
    wire N__19083;
    wire N__19082;
    wire N__19079;
    wire N__19076;
    wire N__19073;
    wire N__19070;
    wire N__19065;
    wire N__19062;
    wire N__19059;
    wire N__19056;
    wire N__19053;
    wire N__19050;
    wire N__19047;
    wire N__19044;
    wire N__19041;
    wire N__19038;
    wire N__19035;
    wire N__19032;
    wire N__19029;
    wire N__19026;
    wire N__19023;
    wire N__19020;
    wire N__19017;
    wire N__19014;
    wire N__19011;
    wire N__19008;
    wire N__19005;
    wire N__19002;
    wire N__18999;
    wire N__18996;
    wire N__18993;
    wire N__18992;
    wire N__18989;
    wire N__18986;
    wire N__18983;
    wire N__18980;
    wire N__18975;
    wire N__18972;
    wire N__18969;
    wire N__18966;
    wire N__18965;
    wire N__18964;
    wire N__18961;
    wire N__18958;
    wire N__18955;
    wire N__18948;
    wire N__18945;
    wire N__18942;
    wire N__18939;
    wire N__18936;
    wire N__18933;
    wire N__18930;
    wire N__18927;
    wire N__18924;
    wire N__18923;
    wire N__18922;
    wire N__18921;
    wire N__18920;
    wire N__18919;
    wire N__18918;
    wire N__18915;
    wire N__18910;
    wire N__18907;
    wire N__18900;
    wire N__18895;
    wire N__18890;
    wire N__18887;
    wire N__18884;
    wire N__18879;
    wire N__18878;
    wire N__18875;
    wire N__18874;
    wire N__18873;
    wire N__18872;
    wire N__18869;
    wire N__18864;
    wire N__18861;
    wire N__18860;
    wire N__18859;
    wire N__18856;
    wire N__18851;
    wire N__18844;
    wire N__18837;
    wire N__18836;
    wire N__18835;
    wire N__18830;
    wire N__18829;
    wire N__18826;
    wire N__18823;
    wire N__18822;
    wire N__18821;
    wire N__18818;
    wire N__18813;
    wire N__18808;
    wire N__18801;
    wire N__18798;
    wire N__18795;
    wire N__18792;
    wire N__18789;
    wire N__18786;
    wire N__18783;
    wire N__18780;
    wire N__18777;
    wire N__18774;
    wire N__18771;
    wire N__18768;
    wire N__18765;
    wire N__18762;
    wire N__18759;
    wire N__18756;
    wire N__18753;
    wire N__18752;
    wire N__18749;
    wire N__18746;
    wire N__18743;
    wire N__18740;
    wire N__18735;
    wire N__18732;
    wire N__18731;
    wire N__18728;
    wire N__18725;
    wire N__18722;
    wire N__18719;
    wire N__18716;
    wire N__18713;
    wire N__18708;
    wire N__18705;
    wire N__18702;
    wire N__18699;
    wire N__18696;
    wire N__18693;
    wire N__18690;
    wire N__18687;
    wire N__18684;
    wire N__18681;
    wire N__18678;
    wire N__18677;
    wire N__18674;
    wire N__18671;
    wire N__18666;
    wire N__18663;
    wire N__18660;
    wire N__18657;
    wire N__18654;
    wire N__18651;
    wire N__18650;
    wire N__18649;
    wire N__18646;
    wire N__18641;
    wire N__18636;
    wire N__18633;
    wire N__18630;
    wire N__18627;
    wire N__18624;
    wire N__18623;
    wire N__18618;
    wire N__18615;
    wire N__18614;
    wire N__18609;
    wire N__18606;
    wire N__18603;
    wire N__18600;
    wire N__18597;
    wire N__18594;
    wire N__18591;
    wire N__18588;
    wire N__18585;
    wire N__18582;
    wire N__18579;
    wire N__18576;
    wire N__18573;
    wire N__18570;
    wire N__18567;
    wire N__18564;
    wire N__18561;
    wire N__18558;
    wire N__18555;
    wire N__18552;
    wire N__18549;
    wire N__18546;
    wire N__18543;
    wire N__18540;
    wire N__18537;
    wire N__18534;
    wire N__18531;
    wire N__18528;
    wire N__18525;
    wire N__18522;
    wire N__18519;
    wire N__18516;
    wire N__18513;
    wire N__18510;
    wire N__18507;
    wire N__18504;
    wire N__18501;
    wire N__18500;
    wire N__18497;
    wire N__18494;
    wire N__18491;
    wire N__18488;
    wire N__18485;
    wire N__18482;
    wire N__18479;
    wire N__18474;
    wire N__18473;
    wire N__18470;
    wire N__18467;
    wire N__18462;
    wire N__18461;
    wire N__18460;
    wire N__18457;
    wire N__18454;
    wire N__18451;
    wire N__18444;
    wire N__18441;
    wire N__18440;
    wire N__18437;
    wire N__18434;
    wire N__18431;
    wire N__18428;
    wire N__18425;
    wire N__18422;
    wire N__18417;
    wire N__18416;
    wire N__18413;
    wire N__18410;
    wire N__18407;
    wire N__18404;
    wire N__18401;
    wire N__18398;
    wire N__18393;
    wire N__18392;
    wire N__18389;
    wire N__18386;
    wire N__18383;
    wire N__18380;
    wire N__18377;
    wire N__18374;
    wire N__18369;
    wire N__18368;
    wire N__18365;
    wire N__18362;
    wire N__18359;
    wire N__18356;
    wire N__18353;
    wire N__18350;
    wire N__18345;
    wire N__18342;
    wire N__18341;
    wire N__18338;
    wire N__18335;
    wire N__18332;
    wire N__18329;
    wire N__18326;
    wire N__18323;
    wire N__18318;
    wire N__18317;
    wire N__18316;
    wire N__18315;
    wire N__18314;
    wire N__18311;
    wire N__18310;
    wire N__18307;
    wire N__18306;
    wire N__18303;
    wire N__18288;
    wire N__18285;
    wire N__18282;
    wire N__18279;
    wire N__18276;
    wire N__18273;
    wire N__18270;
    wire N__18267;
    wire N__18264;
    wire N__18261;
    wire N__18258;
    wire N__18255;
    wire N__18252;
    wire N__18249;
    wire N__18246;
    wire N__18243;
    wire N__18240;
    wire N__18237;
    wire N__18234;
    wire N__18231;
    wire N__18228;
    wire N__18225;
    wire N__18222;
    wire N__18219;
    wire N__18216;
    wire N__18213;
    wire N__18210;
    wire N__18207;
    wire N__18204;
    wire N__18201;
    wire N__18198;
    wire N__18195;
    wire N__18192;
    wire N__18189;
    wire N__18186;
    wire N__18183;
    wire N__18180;
    wire N__18177;
    wire N__18174;
    wire N__18171;
    wire N__18168;
    wire N__18165;
    wire N__18162;
    wire N__18159;
    wire N__18156;
    wire N__18153;
    wire N__18150;
    wire N__18147;
    wire N__18144;
    wire N__18141;
    wire N__18138;
    wire N__18135;
    wire N__18132;
    wire N__18129;
    wire N__18126;
    wire N__18123;
    wire N__18120;
    wire N__18117;
    wire N__18114;
    wire N__18111;
    wire N__18108;
    wire N__18105;
    wire N__18102;
    wire N__18099;
    wire N__18096;
    wire N__18093;
    wire N__18090;
    wire N__18087;
    wire N__18084;
    wire N__18081;
    wire N__18078;
    wire N__18075;
    wire N__18072;
    wire N__18069;
    wire N__18066;
    wire N__18063;
    wire N__18060;
    wire N__18057;
    wire N__18054;
    wire N__18051;
    wire N__18048;
    wire N__18045;
    wire N__18042;
    wire N__18039;
    wire N__18036;
    wire N__18033;
    wire N__18030;
    wire N__18027;
    wire N__18024;
    wire N__18021;
    wire N__18018;
    wire N__18015;
    wire N__18012;
    wire N__18009;
    wire N__18006;
    wire N__18003;
    wire N__18000;
    wire N__17997;
    wire N__17994;
    wire N__17991;
    wire N__17988;
    wire N__17985;
    wire N__17982;
    wire N__17979;
    wire N__17976;
    wire N__17973;
    wire N__17970;
    wire N__17967;
    wire N__17964;
    wire N__17961;
    wire N__17958;
    wire N__17955;
    wire N__17952;
    wire N__17949;
    wire N__17946;
    wire N__17943;
    wire N__17940;
    wire N__17937;
    wire N__17934;
    wire N__17931;
    wire N__17930;
    wire N__17927;
    wire N__17924;
    wire N__17921;
    wire N__17918;
    wire N__17915;
    wire N__17912;
    wire N__17909;
    wire N__17906;
    wire N__17903;
    wire N__17898;
    wire N__17897;
    wire N__17894;
    wire N__17891;
    wire N__17888;
    wire N__17883;
    wire N__17880;
    wire N__17877;
    wire N__17874;
    wire N__17871;
    wire N__17868;
    wire N__17865;
    wire N__17862;
    wire N__17859;
    wire N__17856;
    wire N__17853;
    wire N__17850;
    wire N__17847;
    wire N__17844;
    wire N__17841;
    wire N__17838;
    wire N__17835;
    wire N__17832;
    wire N__17829;
    wire N__17826;
    wire N__17823;
    wire N__17820;
    wire N__17817;
    wire N__17814;
    wire N__17811;
    wire N__17808;
    wire N__17805;
    wire N__17802;
    wire N__17799;
    wire N__17796;
    wire N__17793;
    wire N__17790;
    wire N__17787;
    wire N__17784;
    wire N__17781;
    wire N__17778;
    wire N__17775;
    wire N__17772;
    wire N__17769;
    wire N__17766;
    wire N__17763;
    wire N__17760;
    wire N__17757;
    wire N__17754;
    wire N__17751;
    wire N__17748;
    wire N__17745;
    wire N__17742;
    wire N__17739;
    wire N__17736;
    wire N__17733;
    wire N__17730;
    wire N__17727;
    wire N__17724;
    wire N__17721;
    wire N__17718;
    wire N__17715;
    wire N__17714;
    wire N__17709;
    wire N__17706;
    wire N__17703;
    wire N__17700;
    wire N__17697;
    wire N__17694;
    wire N__17691;
    wire N__17688;
    wire N__17685;
    wire N__17682;
    wire N__17679;
    wire N__17676;
    wire N__17673;
    wire N__17670;
    wire N__17667;
    wire N__17664;
    wire N__17661;
    wire N__17658;
    wire N__17655;
    wire N__17652;
    wire N__17649;
    wire N__17646;
    wire N__17643;
    wire N__17640;
    wire N__17637;
    wire N__17634;
    wire N__17631;
    wire N__17628;
    wire N__17625;
    wire N__17622;
    wire N__17621;
    wire N__17620;
    wire N__17619;
    wire N__17618;
    wire N__17617;
    wire N__17616;
    wire N__17615;
    wire N__17612;
    wire N__17605;
    wire N__17596;
    wire N__17591;
    wire N__17588;
    wire N__17585;
    wire N__17582;
    wire N__17577;
    wire N__17574;
    wire N__17571;
    wire N__17568;
    wire N__17565;
    wire N__17562;
    wire N__17559;
    wire N__17556;
    wire N__17553;
    wire N__17550;
    wire N__17549;
    wire N__17546;
    wire N__17543;
    wire N__17538;
    wire N__17535;
    wire N__17534;
    wire N__17531;
    wire N__17528;
    wire N__17525;
    wire N__17520;
    wire N__17517;
    wire N__17514;
    wire N__17511;
    wire N__17508;
    wire N__17505;
    wire N__17502;
    wire N__17499;
    wire N__17496;
    wire N__17493;
    wire N__17490;
    wire N__17487;
    wire N__17484;
    wire N__17481;
    wire N__17478;
    wire N__17475;
    wire N__17472;
    wire N__17469;
    wire N__17466;
    wire N__17463;
    wire N__17460;
    wire N__17457;
    wire N__17454;
    wire N__17451;
    wire N__17448;
    wire N__17445;
    wire N__17442;
    wire N__17439;
    wire N__17436;
    wire N__17433;
    wire N__17430;
    wire N__17427;
    wire N__17424;
    wire N__17421;
    wire N__17418;
    wire N__17415;
    wire N__17412;
    wire N__17409;
    wire N__17406;
    wire N__17403;
    wire N__17400;
    wire N__17397;
    wire N__17394;
    wire N__17391;
    wire N__17388;
    wire N__17385;
    wire N__17382;
    wire N__17379;
    wire N__17376;
    wire N__17373;
    wire N__17370;
    wire N__17367;
    wire N__17364;
    wire N__17361;
    wire N__17358;
    wire N__17355;
    wire N__17352;
    wire N__17349;
    wire N__17346;
    wire N__17343;
    wire N__17340;
    wire N__17337;
    wire N__17334;
    wire N__17331;
    wire N__17328;
    wire N__17325;
    wire N__17322;
    wire N__17319;
    wire N__17316;
    wire N__17313;
    wire N__17310;
    wire N__17307;
    wire N__17304;
    wire N__17301;
    wire N__17298;
    wire N__17295;
    wire N__17292;
    wire N__17289;
    wire N__17286;
    wire VCCG0;
    wire GNDG0;
    wire bfn_1_6_0_;
    wire \pid_alt.un1_error_d_reg_2_1 ;
    wire \pid_alt.un1_error_d_reg_1_16 ;
    wire \pid_alt.un1_error_d_reg_add_1_cry_0 ;
    wire \pid_alt.un1_error_d_reg_2_2 ;
    wire \pid_alt.un1_error_d_reg_1_17 ;
    wire \pid_alt.un1_error_d_reg_add_1_cry_1 ;
    wire \pid_alt.un1_error_d_reg_2_3 ;
    wire \pid_alt.un1_error_d_reg_1_18 ;
    wire \pid_alt.un1_error_d_reg_add_1_cry_2 ;
    wire \pid_alt.un1_error_d_reg_2_4 ;
    wire \pid_alt.un1_error_d_reg_1_19 ;
    wire \pid_alt.un1_error_d_reg_add_1_cry_3 ;
    wire \pid_alt.un1_error_d_reg_2_5 ;
    wire \pid_alt.un1_error_d_reg_1_20 ;
    wire \pid_alt.un1_error_d_reg_add_1_cry_4 ;
    wire \pid_alt.un1_error_d_reg_2_6 ;
    wire \pid_alt.un1_error_d_reg_1_21 ;
    wire \pid_alt.un1_error_d_reg_add_1_cry_5 ;
    wire \pid_alt.un1_error_d_reg_1_22 ;
    wire \pid_alt.un1_error_d_reg_2_7 ;
    wire \pid_alt.un1_error_d_reg_add_1_cry_6 ;
    wire \pid_alt.un1_error_d_reg_add_1_cry_7 ;
    wire \pid_alt.un1_error_d_reg_1_23 ;
    wire \pid_alt.un1_error_d_reg_2_8 ;
    wire bfn_1_7_0_;
    wire \pid_alt.un1_error_d_reg_2_9 ;
    wire \pid_alt.un1_error_d_reg_add_1_cry_8 ;
    wire \pid_alt.un1_error_d_reg_2_10 ;
    wire \pid_alt.un1_error_d_reg_add_1_cry_9 ;
    wire \pid_alt.un1_error_d_reg_2_11 ;
    wire \pid_alt.un1_error_d_reg_add_1_cry_10 ;
    wire \pid_alt.un1_error_d_reg_2_12 ;
    wire \pid_alt.un1_error_d_reg_add_1_cry_11 ;
    wire \pid_alt.un1_error_d_reg_2_13 ;
    wire \pid_alt.un1_error_d_reg_add_1_cry_12 ;
    wire \pid_alt.un1_error_d_reg_2_14 ;
    wire \pid_alt.un1_error_d_reg_add_1_cry_13 ;
    wire \pid_alt.un1_error_d_reg_2_15 ;
    wire \pid_alt.un1_error_d_reg_add_1_cry_14 ;
    wire \pid_alt.un1_error_d_reg_add_1_cry_15 ;
    wire \pid_alt.un1_error_d_reg_1_24 ;
    wire \pid_alt.un1_error_d_reg_2_16 ;
    wire bfn_1_8_0_;
    wire \pid_alt.O_10 ;
    wire \pid_alt.un1_error_d_reg_2_0 ;
    wire \pid_alt.un1_error_d_reg_1_15 ;
    wire \pid_alt.O_13 ;
    wire \pid_alt.O_11 ;
    wire \pid_alt.O_5 ;
    wire \pid_alt.O_14 ;
    wire \pid_alt.O_6 ;
    wire \pid_alt.O_12 ;
    wire \pid_alt.O_9 ;
    wire \pid_alt.O_7 ;
    wire \pid_alt.O_1_4 ;
    wire \pid_alt.error_filt_prevZ0Z_0 ;
    wire \pid_alt.error_filt ;
    wire \pid_alt.O_2_5 ;
    wire \pid_alt.error_filt_0 ;
    wire bfn_1_16_0_;
    wire \pid_alt.O_3_6 ;
    wire \pid_alt.O_2_6 ;
    wire \pid_alt.error_filt_cry_0 ;
    wire \pid_alt.O_3_7 ;
    wire \pid_alt.O_2_7 ;
    wire \pid_alt.error_filt_cry_1 ;
    wire \pid_alt.O_3_8 ;
    wire \pid_alt.O_2_8 ;
    wire \pid_alt.error_filt_cry_2 ;
    wire \pid_alt.O_3_9 ;
    wire \pid_alt.O_2_9 ;
    wire \pid_alt.error_filt_cry_3 ;
    wire \pid_alt.O_2_10 ;
    wire \pid_alt.O_3_10 ;
    wire \pid_alt.error_filt_cry_4 ;
    wire \pid_alt.O_3_11 ;
    wire \pid_alt.O_2_11 ;
    wire \pid_alt.error_filt_cry_5 ;
    wire \pid_alt.O_2_12 ;
    wire \pid_alt.O_3_12 ;
    wire \pid_alt.error_filt_cry_6 ;
    wire \pid_alt.error_filt_cry_7 ;
    wire \pid_alt.O_3_13 ;
    wire \pid_alt.O_2_13 ;
    wire bfn_1_17_0_;
    wire \pid_alt.O_3_14 ;
    wire \pid_alt.O_2_14 ;
    wire \pid_alt.error_filt_cry_8 ;
    wire \pid_alt.O_1_15 ;
    wire \pid_alt.error_filt_cry_9 ;
    wire \pid_alt.O_1_16 ;
    wire \pid_alt.error_filt_cry_10 ;
    wire \pid_alt.O_1_17 ;
    wire \pid_alt.error_filt_cry_11 ;
    wire \pid_alt.O_1_18 ;
    wire \pid_alt.error_filt_cry_12 ;
    wire \pid_alt.O_1_19 ;
    wire \pid_alt.error_filt_cry_13 ;
    wire \pid_alt.O_1_20 ;
    wire \pid_alt.error_filt_cry_14 ;
    wire \pid_alt.error_filt_cry_15 ;
    wire bfn_1_18_0_;
    wire \pid_alt.error_filt_cry_16 ;
    wire \pid_alt.error_filt_cry_17 ;
    wire \pid_alt.error_filt_cry_18 ;
    wire \pid_alt.error_filt_cry_19 ;
    wire \pid_alt.error_filt_cry_20 ;
    wire \pid_alt.O_1_21 ;
    wire \pid_alt.error_filt_cry_21 ;
    wire \pid_alt.O_1_11 ;
    wire \pid_alt.O_1_12 ;
    wire \pid_alt.O_1_10 ;
    wire \pid_alt.O_0_17 ;
    wire \pid_alt.O_0_20 ;
    wire \pid_alt.O_0_23 ;
    wire \pid_alt.O_1_13 ;
    wire \pid_alt.O_0_21 ;
    wire \pid_alt.O_0_24 ;
    wire \pid_alt.O_0_18 ;
    wire \pid_alt.O_0_19 ;
    wire \pid_alt.error_p_regZ0Z_17 ;
    wire \pid_alt.error_d_reg_prevZ0Z_17 ;
    wire \pid_alt.error_d_regZ0Z_17 ;
    wire alt_kd_2;
    wire alt_kd_3;
    wire alt_kd_7;
    wire alt_kd_1;
    wire alt_kd_0;
    wire \pid_alt.g0_0_0_cascade_ ;
    wire \pid_alt.error_d_regZ0Z_19 ;
    wire \pid_alt.error_d_reg_prevZ0Z_19 ;
    wire \pid_alt.error_p_regZ0Z_19 ;
    wire \pid_alt.O_1_6 ;
    wire \pid_alt.O_1_5 ;
    wire \pid_alt.O_1_14 ;
    wire alt_kp_3;
    wire alt_kp_1;
    wire alt_kp_7;
    wire alt_kp_2;
    wire \pid_alt.O_0_22 ;
    wire alt_kd_6;
    wire alt_kd_5;
    wire \pid_alt.O_4 ;
    wire \pid_alt.N_1074_0 ;
    wire \pid_alt.N_5_0 ;
    wire \pid_alt.g1_1 ;
    wire \pid_alt.N_1080_0_cascade_ ;
    wire \pid_alt.error_d_reg_fastZ0Z_1 ;
    wire \pid_alt.N_3_0 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI0J511_3Z0Z_2 ;
    wire \pid_alt.error_d_reg_esr_RNITF511_0Z0Z_1_cascade_ ;
    wire \pid_alt.error_p_reg_esr_RNIL2AQ1Z0Z_0 ;
    wire \pid_alt.N_1078_0 ;
    wire \pid_alt.error_p_regZ0Z_1 ;
    wire \pid_alt.error_d_reg_prevZ0Z_1 ;
    wire \pid_alt.error_d_regZ0Z_1 ;
    wire \pid_alt.N_1074_1 ;
    wire \pid_alt.N_3_1_cascade_ ;
    wire \pid_alt.error_d_reg_prev_esr_RNI0J511_1Z0Z_2 ;
    wire \pid_alt.g1_0 ;
    wire \pid_alt.error_d_reg_prevZ0Z_20 ;
    wire \pid_alt.error_d_regZ0Z_20 ;
    wire \pid_alt.O_1_7 ;
    wire alt_kp_0;
    wire alt_kp_6;
    wire alt_kp_5;
    wire \pid_alt.O_0_16 ;
    wire alt_kd_4;
    wire \Commands_frame_decoder.source_alt_kd_1_sqmuxa ;
    wire \pid_alt.g0_4_0 ;
    wire \pid_alt.error_d_reg_prevZ0Z_2 ;
    wire \pid_alt.error_p_regZ0Z_2 ;
    wire \pid_alt.error_d_regZ0Z_2 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI3M511_0Z0Z_3 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI0J511_0Z0Z_2_cascade_ ;
    wire \pid_alt.error_d_reg_prev_esr_RNII5LS3Z0Z_2 ;
    wire \pid_alt.error_p_regZ0Z_3 ;
    wire \pid_alt.error_d_reg_prevZ0Z_3 ;
    wire \pid_alt.error_d_regZ0Z_3 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI53IMZ0Z_18 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI86IM_0Z0Z_19 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI53IMZ0Z_18_cascade_ ;
    wire \pid_alt.error_p_regZ0Z_18 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI53IM_0Z0Z_18_cascade_ ;
    wire \pid_alt.error_d_regZ0Z_18 ;
    wire \pid_alt.error_d_reg_prevZ0Z_18 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI53IM_0Z0Z_18 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI20IMZ0Z_17 ;
    wire \pid_alt.error_p_regZ0Z_13 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIMJHM_0Z0Z_13_cascade_ ;
    wire \pid_alt.error_d_reg_prev_esr_RNIJGHMZ0Z_12 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIMJHM_0Z0Z_13 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIJGHMZ0Z_12_cascade_ ;
    wire \pid_alt.error_p_regZ0Z_12 ;
    wire \pid_alt.error_d_reg_prevZ0Z_12 ;
    wire \pid_alt.error_d_regZ0Z_12 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIJGHM_0Z0Z_12_cascade_ ;
    wire \pid_alt.error_d_regZ0Z_13 ;
    wire \pid_alt.error_d_reg_prevZ0Z_13 ;
    wire \pid_alt.O_0_15 ;
    wire \dron_frame_decoder_1.WDT10lto9_3_cascade_ ;
    wire \dron_frame_decoder_1.WDT10lt12_0_cascade_ ;
    wire \dron_frame_decoder_1.WDT10_0_i_1 ;
    wire \dron_frame_decoder_1.WDT10lt12_0 ;
    wire \dron_frame_decoder_1.WDT10lt14_0 ;
    wire \pid_alt.state_1_0_0 ;
    wire \pid_alt.error_p_regZ0Z_11 ;
    wire \pid_alt.error_d_reg_prevZ0Z_11 ;
    wire \pid_alt.error_d_regZ0Z_11 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI7E8R_0Z0Z_11 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIDAHMZ0Z_10 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI7E8R_0Z0Z_11_cascade_ ;
    wire \pid_alt.error_d_reg_prev_esr_RNIJGHM_0Z0Z_12 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI7E8RZ0Z_11 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIOFGB2Z0Z_10_cascade_ ;
    wire \pid_alt.error_d_reg_prev_esr_RNIVSHMZ0Z_16 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI20IM_0Z0Z_17 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIVSHMZ0Z_16_cascade_ ;
    wire \pid_alt.error_p_regZ0Z_16 ;
    wire \pid_alt.error_d_reg_prevZ0Z_16 ;
    wire \pid_alt.error_d_regZ0Z_16 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIVSHM_0Z0Z_16 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIVSHM_0Z0Z_16_cascade_ ;
    wire \pid_alt.error_d_reg_prev_esr_RNII5611_0Z0Z_8_cascade_ ;
    wire \pid_alt.error_d_reg_prev_esr_RNIF2611Z0Z_7 ;
    wire \pid_alt.error_d_reg_prev_esr_RNII5611_0Z0Z_8 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIF2611Z0Z_7_cascade_ ;
    wire \pid_alt.error_p_regZ0Z_7 ;
    wire \pid_alt.error_d_reg_prevZ0Z_7 ;
    wire \pid_alt.error_d_regZ0Z_7 ;
    wire \pid_alt.error_p_regZ0Z_8 ;
    wire \pid_alt.error_d_regZ0Z_8 ;
    wire \pid_alt.error_d_reg_prevZ0Z_8 ;
    wire \pid_alt.error_d_reg_prev_esr_RNISPHMZ0Z_15 ;
    wire \pid_alt.error_d_reg_prevZ0Z_0 ;
    wire \pid_alt.error_d_reg_prevZ0Z_15 ;
    wire \pid_alt.error_p_regZ0Z_15 ;
    wire \pid_alt.error_d_regZ0Z_15 ;
    wire \pid_alt.error_d_reg_prev_esr_RNISPHM_0Z0Z_15 ;
    wire \pid_alt.error_d_reg_prev_esr_RNISPHM_0Z0Z_15_cascade_ ;
    wire \pid_alt.error_d_reg_prev_esr_RNIPMHMZ0Z_14 ;
    wire \pid_alt.error_p_regZ0Z_14 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIPMHM_0Z0Z_14_cascade_ ;
    wire \pid_alt.error_d_regZ0Z_14 ;
    wire \pid_alt.error_d_reg_prevZ0Z_14 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIMJHMZ0Z_13 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIPMHM_0Z0Z_14 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIMMKM_0Z0Z_23_cascade_ ;
    wire \pid_alt.error_d_reg_prevZ0Z_22 ;
    wire \pid_alt.error_d_regZ0Z_22 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIKKKMZ0Z_22 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIMMKM_0Z0Z_23 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIKKKMZ0Z_22_cascade_ ;
    wire \pid_alt.error_d_regZ0Z_23 ;
    wire \pid_alt.error_d_reg_prevZ0Z_23 ;
    wire \pid_alt.O_1_8 ;
    wire \dron_frame_decoder_1.WDT10_0_i ;
    wire \dron_frame_decoder_1.WDTZ0Z_0 ;
    wire bfn_7_7_0_;
    wire \dron_frame_decoder_1.WDTZ0Z_1 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_0 ;
    wire \dron_frame_decoder_1.WDTZ0Z_2 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_1 ;
    wire \dron_frame_decoder_1.WDTZ0Z_3 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_2 ;
    wire \dron_frame_decoder_1.WDTZ0Z_4 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_3 ;
    wire \dron_frame_decoder_1.WDTZ0Z_5 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_4 ;
    wire \dron_frame_decoder_1.WDTZ0Z_6 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_5 ;
    wire \dron_frame_decoder_1.WDTZ0Z_7 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_6 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_7 ;
    wire \dron_frame_decoder_1.WDTZ0Z_8 ;
    wire bfn_7_8_0_;
    wire \dron_frame_decoder_1.WDTZ0Z_9 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_8 ;
    wire \dron_frame_decoder_1.WDTZ0Z_10 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_9 ;
    wire \dron_frame_decoder_1.WDTZ0Z_11 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_10 ;
    wire \dron_frame_decoder_1.WDTZ0Z_12 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_11 ;
    wire \dron_frame_decoder_1.WDTZ0Z_13 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_12 ;
    wire \dron_frame_decoder_1.WDTZ0Z_14 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_13 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_14 ;
    wire \dron_frame_decoder_1.WDTZ0Z_15 ;
    wire \dron_frame_decoder_1.stateZ0Z_3 ;
    wire \dron_frame_decoder_1.stateZ0Z_2 ;
    wire \dron_frame_decoder_1.N_188_4_cascade_ ;
    wire \dron_frame_decoder_1.state_ns_0_i_a2_0_0_3 ;
    wire \Commands_frame_decoder.source_CH2data_1_sqmuxa_cascade_ ;
    wire \dron_frame_decoder_1.state_ns_0_i_a2_1_0Z0Z_3_cascade_ ;
    wire \dron_frame_decoder_1.N_188_4 ;
    wire \dron_frame_decoder_1.state_ns_0_i_a2_1Z0Z_3_cascade_ ;
    wire \dron_frame_decoder_1.state_RNO_0Z0Z_0_cascade_ ;
    wire \dron_frame_decoder_1.state_ns_0_i_a2_0_0_1Z0Z_1_cascade_ ;
    wire \dron_frame_decoder_1.state_ns_0_i_a2_0_1 ;
    wire \dron_frame_decoder_1.state_ns_0_i_a2_1Z0Z_3 ;
    wire \dron_frame_decoder_1.state_ns_0_i_a2_0_1_cascade_ ;
    wire \pid_alt.error_d_reg_esr_RNITF511_2Z0Z_1 ;
    wire \pid_alt.error_p_regZ0Z_0 ;
    wire \pid_alt.error_d_regZ0Z_0 ;
    wire \dron_frame_decoder_1.stateZ0Z_1 ;
    wire \dron_frame_decoder_1.state_RNO_1Z0Z_0 ;
    wire \pid_alt.error_d_reg_prev_i_0 ;
    wire bfn_7_13_0_;
    wire \pid_alt.error_p_reg_esr_RNI3SMI1Z0Z_0 ;
    wire \pid_alt.un1_pid_prereg_un1_pid_prereg_0_cry_0_c_THRU_CO ;
    wire \pid_alt.error_p_reg_esr_RNIFPN33Z0Z_0 ;
    wire \pid_alt.un1_pid_prereg_0_cry_0 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIF0465Z0Z_2 ;
    wire \pid_alt.un1_pid_prereg_0_cry_1 ;
    wire \pid_alt.error_d_reg_prev_esr_RNILDG87Z0Z_2 ;
    wire \pid_alt.un1_pid_prereg_0_cry_2 ;
    wire \pid_alt.un1_pid_prereg_0_cry_3 ;
    wire \pid_alt.un1_pid_prereg_0_cry_4 ;
    wire \pid_alt.un1_pid_prereg_0_cry_5 ;
    wire \pid_alt.un1_pid_prereg_0_cry_6 ;
    wire bfn_7_14_0_;
    wire \pid_alt.error_d_reg_prev_esr_RNI5G6Q5Z0Z_7 ;
    wire \pid_alt.un1_pid_prereg_0_cry_7 ;
    wire \pid_alt.un1_pid_prereg_0_cry_8 ;
    wire \pid_alt.un1_pid_prereg_0_cry_9 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIKQBI4Z0Z_10 ;
    wire \pid_alt.un1_pid_prereg_0_cry_10 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIP92N4Z0Z_11 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIOFGB2Z0Z_10 ;
    wire \pid_alt.un1_pid_prereg_0_cry_11 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIT4AF4Z0Z_12 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI1QHB2Z0Z_11 ;
    wire \pid_alt.un1_pid_prereg_0_cry_12 ;
    wire \pid_alt.error_d_reg_prev_esr_RNICQF44Z0Z_13 ;
    wire \pid_alt.error_d_reg_prev_esr_RNISAO32Z0Z_12 ;
    wire \pid_alt.un1_pid_prereg_0_cry_13 ;
    wire \pid_alt.un1_pid_prereg_0_cry_14 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI88G14Z0Z_14 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIGFN02Z0Z_13 ;
    wire bfn_7_15_0_;
    wire \pid_alt.error_d_reg_prev_esr_RNIOQI14Z0Z_15 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIOOO02Z0Z_14 ;
    wire \pid_alt.pid_preregZ0Z_16 ;
    wire \pid_alt.un1_pid_prereg_0_cry_15 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI8DL14Z0Z_16 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI02Q02Z0Z_15 ;
    wire \pid_alt.pid_preregZ0Z_17 ;
    wire \pid_alt.un1_pid_prereg_0_cry_16 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIOVN14Z0Z_17 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI8BR02Z0Z_16 ;
    wire \pid_alt.pid_preregZ0Z_18 ;
    wire \pid_alt.un1_pid_prereg_0_cry_17 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI8IQ14Z0Z_18 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIGKS02Z0Z_17 ;
    wire \pid_alt.pid_preregZ0Z_19 ;
    wire \pid_alt.un1_pid_prereg_0_cry_18 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIK3024Z0Z_19 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIOTT02Z0Z_18 ;
    wire \pid_alt.un1_pid_prereg_0_cry_19 ;
    wire \pid_alt.un1_pid_prereg_0_cry_20 ;
    wire \pid_alt.un1_pid_prereg_0_cry_21 ;
    wire \pid_alt.un1_pid_prereg_0_cry_22 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI8IS34Z0Z_22 ;
    wire bfn_7_16_0_;
    wire \pid_alt.un1_pid_prereg_0_cry_23 ;
    wire \pid_alt.un1_pid_prereg_0_cry_24 ;
    wire \pid_alt.un1_pid_prereg_0_cry_25 ;
    wire \pid_alt.un1_pid_prereg_0_cry_26 ;
    wire \pid_alt.un1_pid_prereg_0_cry_27 ;
    wire \pid_alt.un1_pid_prereg_0_cry_28 ;
    wire \pid_alt.un1_pid_prereg_0_cry_29 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI8JT34Z0Z_26 ;
    wire \pid_alt.error_d_reg_prev_esr_RNISSKMZ0Z_26_cascade_ ;
    wire \pid_alt.error_d_reg_prev_esr_RNIMRU12Z0Z_26 ;
    wire \pid_alt.error_d_reg_prev_esr_RNISSKMZ0Z_26 ;
    wire \pid_alt.un1_pid_prereg_296_1_cascade_ ;
    wire \pid_alt.error_d_reg_prev_esr_RNIKQJO2Z0Z_26 ;
    wire \pid_alt.error_d_regZ0Z_27 ;
    wire \pid_alt.error_d_reg_prevZ0Z_27 ;
    wire bfn_7_19_0_;
    wire \pid_alt.error_1 ;
    wire \pid_alt.error_cry_0 ;
    wire \pid_alt.error_2 ;
    wire \pid_alt.error_cry_1 ;
    wire \pid_alt.error_3 ;
    wire \pid_alt.error_cry_2 ;
    wire \pid_alt.error_4 ;
    wire \pid_alt.error_cry_3 ;
    wire alt_command_1;
    wire \pid_alt.error_5 ;
    wire \pid_alt.error_cry_4 ;
    wire alt_command_2;
    wire \pid_alt.error_6 ;
    wire \pid_alt.error_cry_5 ;
    wire alt_command_3;
    wire \pid_alt.error_7 ;
    wire \pid_alt.error_cry_6 ;
    wire \pid_alt.error_cry_7 ;
    wire \pid_alt.error_8 ;
    wire bfn_7_20_0_;
    wire \pid_alt.error_9 ;
    wire \pid_alt.error_cry_8 ;
    wire \pid_alt.error_10 ;
    wire \pid_alt.error_cry_9 ;
    wire \pid_alt.error_11 ;
    wire \pid_alt.error_cry_10 ;
    wire \pid_alt.error_12 ;
    wire \pid_alt.error_cry_11 ;
    wire \pid_alt.error_13 ;
    wire \pid_alt.error_cry_12 ;
    wire \pid_alt.error_14 ;
    wire \pid_alt.error_cry_13 ;
    wire \pid_alt.error_cry_14 ;
    wire \pid_alt.error_15 ;
    wire alt_command_4;
    wire alt_command_5;
    wire alt_command_6;
    wire alt_command_7;
    wire \pid_alt.error_d_reg_prev_esr_RNIOTU12Z0Z_27 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIUUKMZ0Z_27 ;
    wire \pid_alt.un1_pid_prereg_296_1 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIOTU12_0Z0Z_27 ;
    wire \pid_alt.N_410_0 ;
    wire \uart_drone_sync.aux_1__0__0_0 ;
    wire uart_input_drone_c;
    wire \uart_drone_sync.aux_0__0__0_0 ;
    wire \Commands_frame_decoder.WDT8lto13_1_cascade_ ;
    wire \Commands_frame_decoder.WDT_RNI2VDI1Z0Z_10 ;
    wire \Commands_frame_decoder.WDT8lto9_3_cascade_ ;
    wire \Commands_frame_decoder.WDT8lt12_0_cascade_ ;
    wire \Commands_frame_decoder.state_0_sqmuxacf1 ;
    wire \Commands_frame_decoder.WDT_RNII19A1Z0Z_4 ;
    wire \uart_drone_sync.aux_2__0__0_0 ;
    wire \uart_drone_sync.aux_3__0__0_0 ;
    wire \dron_frame_decoder_1.source_data_valid_2_sqmuxa_iZ0 ;
    wire \Commands_frame_decoder.source_offset2data_1_sqmuxa_cascade_ ;
    wire \Commands_frame_decoder.N_322_0_cascade_ ;
    wire \Commands_frame_decoder.state_RNIF38SZ0Z_6 ;
    wire \Commands_frame_decoder.N_354 ;
    wire \Commands_frame_decoder.source_offset2data_1_sqmuxa ;
    wire \Commands_frame_decoder.stateZ0Z_8 ;
    wire \dron_frame_decoder_1.un1_sink_data_valid_5_i_0 ;
    wire \dron_frame_decoder_1.un1_sink_data_valid_5_i_0_cascade_ ;
    wire \dron_frame_decoder_1.stateZ0Z_5 ;
    wire \dron_frame_decoder_1.stateZ0Z_4 ;
    wire \dron_frame_decoder_1.WDT_RNIPI9R2Z0Z_15 ;
    wire \dron_frame_decoder_1.stateZ0Z_7 ;
    wire bfn_8_11_0_;
    wire \pid_alt.un9lto29_i_a2 ;
    wire \pid_alt.un9lto29_i_a2_0 ;
    wire \pid_alt.un9lto29_i_a2_1 ;
    wire \pid_alt.un9lto29_i_a2_2 ;
    wire \pid_alt.un9lto29_i_a2_3 ;
    wire \pid_alt.un9lto29_i_a2_4 ;
    wire \pid_alt.N_232_i ;
    wire \pid_alt.un9lto29_i_a2_5 ;
    wire \pid_alt.un9lto29_i_a2_6 ;
    wire bfn_8_12_0_;
    wire \dron_frame_decoder_1.stateZ0Z_0 ;
    wire \dron_frame_decoder_1.state_ns_i_i_a2_2_0_0 ;
    wire \pid_alt.pid_preregZ0Z_22 ;
    wire \pid_alt.pid_preregZ0Z_21 ;
    wire \pid_alt.pid_preregZ0Z_23 ;
    wire \pid_alt.pid_preregZ0Z_20 ;
    wire \pid_alt.source_pid10lt4_0 ;
    wire \pid_alt.un9lto29_i_a2_2_and ;
    wire \pid_alt.pid_preregZ0Z_28 ;
    wire \pid_alt.pid_preregZ0Z_15 ;
    wire \pid_alt.pid_preregZ0Z_29 ;
    wire \pid_alt.pid_preregZ0Z_14 ;
    wire \pid_alt.error_d_reg_prev_esr_RNICV511_0Z0Z_6 ;
    wire \pid_alt.error_d_reg_prev_esr_RNICV511_0Z0Z_6_cascade_ ;
    wire \pid_alt.error_d_reg_prev_esr_RNI171A6Z0Z_5 ;
    wire \pid_alt.error_d_reg_prev_esr_RNICUVC3Z0Z_4 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI9S511_0Z0Z_5 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI9S511_0Z0Z_5_cascade_ ;
    wire \pid_alt.error_d_reg_prev_esr_RNIOGSO6Z0Z_4 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIL8611Z0Z_9_cascade_ ;
    wire \pid_alt.error_d_reg_prev_esr_RNICI045Z0Z_9 ;
    wire \pid_alt.error_p_regZ0Z_10 ;
    wire \pid_alt.error_d_reg_prevZ0Z_10 ;
    wire \pid_alt.error_d_regZ0Z_10 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIG75T2Z0Z_8 ;
    wire \pid_alt.error_p_regZ0Z_9 ;
    wire \pid_alt.error_d_reg_prevZ0Z_9 ;
    wire \pid_alt.error_d_regZ0Z_9 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIL8611_0Z0Z_9 ;
    wire \pid_alt.error_d_reg_prev_esr_RNII5611Z0Z_8 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI7T3T2Z0Z_7 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIL8611_0Z0Z_9_cascade_ ;
    wire \pid_alt.error_d_reg_prev_esr_RNIN49Q5Z0Z_8 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIL81T2Z0Z_5 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIJR3Q5Z0Z_6 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIGGKM_0Z0Z_20 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI86IMZ0Z_19 ;
    wire \dron_frame_decoder_1.state_RNI3T3K1Z0Z_7 ;
    wire \pid_alt.error_d_reg_prevZ0Z_26 ;
    wire \pid_alt.error_d_regZ0Z_26 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIL8611Z0Z_9 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIDAHM_0Z0Z_10 ;
    wire \pid_alt.error_d_reg_prev_esr_RNISAR62Z0Z_9 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI27U12Z0Z_21 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIIIKMZ0Z_21 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIKKKM_0Z0Z_22 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIIIKMZ0Z_21_cascade_ ;
    wire \pid_alt.error_d_reg_prev_esr_RNI0AS34Z0Z_21 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIU2U12Z0Z_20 ;
    wire \pid_alt.error_d_reg_prevZ0Z_21 ;
    wire \pid_alt.error_d_regZ0Z_21 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIIIKM_0Z0Z_21 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIS5212Z0Z_19 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIGGKMZ0Z_20 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIIIKM_0Z0Z_21_cascade_ ;
    wire \pid_alt.error_d_reg_prev_esr_RNIQ8034Z0Z_20 ;
    wire \pid_alt.drone_altitude_i_0 ;
    wire \pid_alt.error_axbZ0Z_3 ;
    wire drone_altitude_i_10;
    wire drone_altitude_i_11;
    wire \pid_alt.error_axbZ0Z_1 ;
    wire \pid_alt.error_axbZ0Z_12 ;
    wire \pid_alt.error_axbZ0Z_13 ;
    wire \pid_alt.error_axbZ0Z_14 ;
    wire \pid_alt.error_axbZ0Z_2 ;
    wire alt_ki_0;
    wire drone_altitude_i_9;
    wire alt_command_0;
    wire \pid_alt.O_1_9 ;
    wire uart_input_pc_c;
    wire \Commands_frame_decoder.state_0_sqmuxa ;
    wire \Commands_frame_decoder.WDTZ0Z_0 ;
    wire bfn_9_5_0_;
    wire \Commands_frame_decoder.WDTZ0Z_1 ;
    wire \Commands_frame_decoder.un1_WDT_cry_0 ;
    wire \Commands_frame_decoder.WDTZ0Z_2 ;
    wire \Commands_frame_decoder.un1_WDT_cry_1 ;
    wire \Commands_frame_decoder.WDTZ0Z_3 ;
    wire \Commands_frame_decoder.un1_WDT_cry_2 ;
    wire \Commands_frame_decoder.WDTZ0Z_4 ;
    wire \Commands_frame_decoder.un1_WDT_cry_3 ;
    wire \Commands_frame_decoder.WDTZ0Z_5 ;
    wire \Commands_frame_decoder.un1_WDT_cry_4 ;
    wire \Commands_frame_decoder.WDTZ0Z_6 ;
    wire \Commands_frame_decoder.un1_WDT_cry_5 ;
    wire \Commands_frame_decoder.WDTZ0Z_7 ;
    wire \Commands_frame_decoder.un1_WDT_cry_6 ;
    wire \Commands_frame_decoder.un1_WDT_cry_7 ;
    wire \Commands_frame_decoder.WDTZ0Z_8 ;
    wire bfn_9_6_0_;
    wire \Commands_frame_decoder.WDTZ0Z_9 ;
    wire \Commands_frame_decoder.un1_WDT_cry_8 ;
    wire \Commands_frame_decoder.WDTZ0Z_10 ;
    wire \Commands_frame_decoder.un1_WDT_cry_9 ;
    wire \Commands_frame_decoder.un1_WDT_cry_10 ;
    wire \Commands_frame_decoder.un1_WDT_cry_11 ;
    wire \Commands_frame_decoder.un1_WDT_cry_12 ;
    wire \Commands_frame_decoder.un1_WDT_cry_13 ;
    wire \Commands_frame_decoder.un1_WDT_cry_14 ;
    wire \Commands_frame_decoder.N_327 ;
    wire \Commands_frame_decoder.stateZ0Z_2 ;
    wire \Commands_frame_decoder.stateZ0Z_11 ;
    wire \Commands_frame_decoder.stateZ0Z_7 ;
    wire \Commands_frame_decoder.WDT8lt14_0 ;
    wire \Commands_frame_decoder.N_358_cascade_ ;
    wire \Commands_frame_decoder.stateZ0Z_10 ;
    wire \Commands_frame_decoder.stateZ0Z_3 ;
    wire \Commands_frame_decoder.source_CH2data_1_sqmuxa ;
    wire \pid_alt.un9lto29_i_a2_3_and ;
    wire \pid_alt.source_pid_1_sqmuxa_0_a2_1_0 ;
    wire \pid_alt.un9lto29_i_a2_4_and ;
    wire \pid_alt.source_pid_1_sqmuxa_0_a2_0_5 ;
    wire \pid_alt.N_123_cascade_ ;
    wire \pid_alt.pid_preregZ0Z_12 ;
    wire \pid_alt.N_123 ;
    wire \pid_alt.N_106_cascade_ ;
    wire \pid_alt.source_pid_1_sqmuxa_0_a2_0 ;
    wire \pid_alt.N_100 ;
    wire \pid_alt.N_91_1_cascade_ ;
    wire \pid_alt.un1_reset_0_i_cascade_ ;
    wire \pid_alt.pid_preregZ0Z_26 ;
    wire \pid_alt.pid_preregZ0Z_25 ;
    wire \pid_alt.pid_preregZ0Z_27 ;
    wire \pid_alt.pid_preregZ0Z_24 ;
    wire \pid_alt.un9lto29_i_a2_5_and ;
    wire \pid_alt.pid_preregZ0Z_13 ;
    wire \pid_alt.N_124 ;
    wire \pid_alt.pid_preregZ0Z_8 ;
    wire \pid_alt.N_12_i ;
    wire \pid_alt.un9lto29_i_a2_0_and ;
    wire \pid_alt.N_96 ;
    wire \pid_alt.pid_preregZ0Z_5 ;
    wire \pid_alt.pid_preregZ0Z_4 ;
    wire \pid_alt.source_pid_1_sqmuxa_0_a2_0_4 ;
    wire \pid_alt.state_RNIFCSD1Z0Z_0 ;
    wire \Commands_frame_decoder.source_CH1data8 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI6P511Z0Z_4 ;
    wire \pid_alt.error_p_regZ0Z_4 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI0BT34Z0Z_25 ;
    wire \pid_alt.error_d_reg_prev_esr_RNISSKM_0Z0Z_26 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIQQKMZ0Z_25 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIINU12Z0Z_25 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIO2T34Z0Z_24 ;
    wire \pid_alt.error_d_reg_prevZ0Z_25 ;
    wire \pid_alt.error_d_regZ0Z_25 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIQQKM_0Z0Z_25 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIQQKM_0Z0Z_25_cascade_ ;
    wire \pid_alt.error_d_reg_prev_esr_RNIEJU12Z0Z_24 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIOOKM_0Z0Z_24_cascade_ ;
    wire \pid_alt.error_d_reg_prev_esr_RNIAFU12Z0Z_23 ;
    wire \pid_alt.error_d_reg_prevZ0Z_24 ;
    wire \pid_alt.error_d_regZ0Z_24 ;
    wire \pid_alt.error_p_regZ0Z_20 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIOOKMZ0Z_24 ;
    wire \pid_alt.error_p_regZ0Z_6 ;
    wire \pid_alt.error_d_reg_prevZ0Z_6 ;
    wire \pid_alt.error_d_regZ0Z_6 ;
    wire drone_altitude_0;
    wire drone_altitude_1;
    wire drone_altitude_2;
    wire drone_altitude_3;
    wire \dron_frame_decoder_1.N_392_0 ;
    wire \Commands_frame_decoder.source_offset3data_1_sqmuxa ;
    wire \Commands_frame_decoder.N_358 ;
    wire \dron_frame_decoder_1.drone_altitude_4 ;
    wire drone_altitude_i_4;
    wire \dron_frame_decoder_1.drone_altitude_5 ;
    wire drone_altitude_i_5;
    wire \dron_frame_decoder_1.drone_altitude_6 ;
    wire drone_altitude_i_6;
    wire \dron_frame_decoder_1.drone_altitude_7 ;
    wire drone_altitude_i_7;
    wire drone_altitude_i_8;
    wire uart_drone_data_2;
    wire \dron_frame_decoder_1.drone_altitude_10 ;
    wire uart_drone_data_4;
    wire drone_altitude_12;
    wire uart_drone_data_5;
    wire drone_altitude_13;
    wire uart_drone_data_6;
    wire drone_altitude_14;
    wire uart_drone_data_7;
    wire drone_altitude_15;
    wire uart_drone_data_0;
    wire \dron_frame_decoder_1.drone_altitude_8 ;
    wire uart_drone_data_1;
    wire \dron_frame_decoder_1.drone_altitude_9 ;
    wire \pid_alt.stateZ0Z_0 ;
    wire \pid_alt.state_0_0 ;
    wire \uart_pc_sync.aux_2__0_Z0Z_0 ;
    wire \uart_pc_sync.aux_0__0_Z0Z_0 ;
    wire \uart_pc_sync.aux_1__0_Z0Z_0 ;
    wire \Commands_frame_decoder.un1_state53_iZ0 ;
    wire \Commands_frame_decoder.WDTZ0Z_13 ;
    wire \Commands_frame_decoder.WDTZ0Z_12 ;
    wire \Commands_frame_decoder.WDTZ0Z_11 ;
    wire \Commands_frame_decoder.WDTZ0Z_15 ;
    wire \Commands_frame_decoder.state_0_sqmuxacf0_1_cascade_ ;
    wire \Commands_frame_decoder.WDTZ0Z_14 ;
    wire \Commands_frame_decoder.state_0_sqmuxacf0 ;
    wire \Commands_frame_decoder.preinitZ0 ;
    wire \Commands_frame_decoder.count_1_sqmuxa ;
    wire \Commands_frame_decoder.stateZ0Z_0 ;
    wire \Commands_frame_decoder.state_ns_0_a4_0_1_1 ;
    wire \Commands_frame_decoder.N_320_0 ;
    wire \Commands_frame_decoder.state_ns_i_a2_2_1Z0Z_0 ;
    wire \Commands_frame_decoder.state_ns_0_a4_0_0_2_cascade_ ;
    wire \Commands_frame_decoder.state_ns_0_a4_0_3_2 ;
    wire \Commands_frame_decoder.stateZ0Z_1 ;
    wire \Commands_frame_decoder.N_364 ;
    wire \Commands_frame_decoder.N_360_cascade_ ;
    wire \Commands_frame_decoder.N_359 ;
    wire \Commands_frame_decoder.state_ns_i_0_0 ;
    wire \Commands_frame_decoder.stateZ0Z_6 ;
    wire alt_kp_4;
    wire \Commands_frame_decoder.stateZ0Z_4 ;
    wire \Commands_frame_decoder.source_CH3data_1_sqmuxa ;
    wire \Commands_frame_decoder.source_CH3data_1_sqmuxa_cascade_ ;
    wire \Commands_frame_decoder.stateZ0Z_5 ;
    wire \Commands_frame_decoder.source_CH4data_1_sqmuxa ;
    wire \Commands_frame_decoder.source_CH4data_1_sqmuxa_cascade_ ;
    wire \uart_drone.data_AuxZ0Z_0 ;
    wire \uart_drone.data_AuxZ0Z_1 ;
    wire \uart_drone.data_AuxZ0Z_2 ;
    wire \uart_drone.data_AuxZ0Z_3 ;
    wire \uart_drone.data_AuxZ0Z_4 ;
    wire \uart_drone.data_AuxZ0Z_5 ;
    wire \uart_drone.data_AuxZ0Z_6 ;
    wire \uart_drone.data_AuxZ0Z_7 ;
    wire \Commands_frame_decoder.source_CH3data_1_sqmuxa_0 ;
    wire \pid_alt.pid_preregZ0Z_6 ;
    wire \pid_alt.pid_preregZ0Z_0 ;
    wire \pid_alt.pid_preregZ0Z_1 ;
    wire \pid_alt.pid_preregZ0Z_2 ;
    wire \pid_alt.N_91_1 ;
    wire \pid_alt.pid_preregZ0Z_3 ;
    wire \Commands_frame_decoder.state_ns_i_a2_1_1Z0Z_0 ;
    wire \pid_alt.error_p_regZ0Z_5 ;
    wire \pid_alt.error_d_reg_prevZ0Z_5 ;
    wire \pid_alt.error_d_regZ0Z_5 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI9S511Z0Z_5 ;
    wire \pid_alt.error_p_reg_esr_RNIFTRL5Z0Z_3 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIRFO19Z0Z_3 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI3M511Z0Z_3 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI6P511_0Z0Z_4 ;
    wire \pid_alt.error_d_reg_prev_esr_RNICISB3Z0Z_3 ;
    wire \pid_alt.error_d_reg_prevZ0Z_4 ;
    wire \Commands_frame_decoder.source_CH4data_1_sqmuxa_0 ;
    wire \Commands_frame_decoder.source_CH1data8lt7_0 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIF2611_0Z0Z_7 ;
    wire \pid_alt.error_d_reg_prev_esr_RNICV511Z0Z_6 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIUI2T2Z0Z_6 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIOOKM_0Z0Z_24 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIMMKMZ0Z_23 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI6BU12Z0Z_22 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIGQS34Z0Z_23 ;
    wire uart_drone_data_3;
    wire \dron_frame_decoder_1.drone_altitude_11 ;
    wire \dron_frame_decoder_1.N_384_0 ;
    wire \uart_pc_sync.aux_3__0_Z0Z_0 ;
    wire bfn_11_6_0_;
    wire \uart_pc.un4_timer_Count_1_cry_1 ;
    wire \uart_pc.un4_timer_Count_1_cry_2 ;
    wire \uart_pc.un4_timer_Count_1_cry_3 ;
    wire \uart_pc.timer_Count_RNO_0Z0Z_2 ;
    wire \uart_pc.timer_Count_RNO_0Z0Z_4 ;
    wire \uart_pc.timer_CountZ0Z_0 ;
    wire \uart_pc.timer_Count_RNO_0Z0Z_1_cascade_ ;
    wire \uart_pc.timer_CountZ1Z_1 ;
    wire \Commands_frame_decoder.state_ns_0_a4_0_0Z0Z_1 ;
    wire \Commands_frame_decoder.state_ns_i_a4_2_0_0_cascade_ ;
    wire \Commands_frame_decoder.stateZ0Z_12 ;
    wire \Commands_frame_decoder.N_330 ;
    wire \Commands_frame_decoder.state_ns_i_a4_2_0_0 ;
    wire \Commands_frame_decoder.countZ0Z_0 ;
    wire \Commands_frame_decoder.countZ0Z_1 ;
    wire \uart_drone.timer_Count_RNIES9Q1Z0Z_2 ;
    wire \uart_drone.timer_Count_RNIES9Q1Z0Z_2_cascade_ ;
    wire \uart_drone.data_rdyc_1_0 ;
    wire \uart_pc.data_rdyc_1 ;
    wire \uart_drone.data_Auxce_0_0_0 ;
    wire \uart_drone.data_Auxce_0_1 ;
    wire frame_decoder_OFF3data_7;
    wire frame_decoder_CH3data_7;
    wire \Commands_frame_decoder.source_CH2data_1_sqmuxa_0 ;
    wire \Commands_frame_decoder.source_offset3data_1_sqmuxa_0 ;
    wire bfn_11_13_0_;
    wire frame_decoder_OFF3data_1;
    wire frame_decoder_CH3data_1;
    wire \scaler_3.un3_source_data_0_cry_0 ;
    wire frame_decoder_CH3data_2;
    wire frame_decoder_OFF3data_2;
    wire \scaler_3.un3_source_data_0_cry_1 ;
    wire frame_decoder_CH3data_3;
    wire frame_decoder_OFF3data_3;
    wire \scaler_3.un3_source_data_0_cry_2 ;
    wire frame_decoder_CH3data_4;
    wire frame_decoder_OFF3data_4;
    wire \scaler_3.un3_source_data_0_cry_3 ;
    wire frame_decoder_CH3data_5;
    wire frame_decoder_OFF3data_5;
    wire \scaler_3.un3_source_data_0_cry_4 ;
    wire frame_decoder_CH3data_6;
    wire frame_decoder_OFF3data_6;
    wire \scaler_3.un3_source_data_0_cry_5 ;
    wire \scaler_3.un3_source_data_0_axb_7 ;
    wire \scaler_3.un3_source_data_0_cry_6 ;
    wire \scaler_3.un3_source_data_0_cry_7 ;
    wire \scaler_3.N_1239_i_l_ofxZ0 ;
    wire bfn_11_14_0_;
    wire \scaler_3.un3_source_data_0_cry_8 ;
    wire \pid_alt.pid_preregZ0Z_7 ;
    wire \pid_alt.pid_preregZ0Z_11 ;
    wire \pid_alt.pid_preregZ0Z_10 ;
    wire \pid_alt.source_pid_1_sqmuxa_0_a2_2_4 ;
    wire \Commands_frame_decoder.stateZ0Z_9 ;
    wire uart_pc_data_rdy;
    wire bfn_11_16_0_;
    wire frame_decoder_CH4data_1;
    wire frame_decoder_OFF4data_1;
    wire \scaler_4.un3_source_data_0_cry_0 ;
    wire frame_decoder_CH4data_2;
    wire frame_decoder_OFF4data_2;
    wire \scaler_4.un3_source_data_0_cry_1 ;
    wire frame_decoder_CH4data_3;
    wire frame_decoder_OFF4data_3;
    wire \scaler_4.un3_source_data_0_cry_2 ;
    wire frame_decoder_CH4data_4;
    wire frame_decoder_OFF4data_4;
    wire \scaler_4.un3_source_data_0_cry_3 ;
    wire frame_decoder_OFF4data_5;
    wire frame_decoder_CH4data_5;
    wire \scaler_4.un3_source_data_0_cry_4 ;
    wire frame_decoder_CH4data_6;
    wire frame_decoder_OFF4data_6;
    wire \scaler_4.un3_source_data_0_cry_5 ;
    wire \scaler_4.un3_source_data_0_cry_6 ;
    wire \scaler_4.un3_source_data_0_cry_7 ;
    wire bfn_11_17_0_;
    wire \scaler_4.un3_source_data_0_cry_8 ;
    wire \scaler_4.un3_source_data_0_axb_7 ;
    wire frame_decoder_CH4data_7;
    wire frame_decoder_OFF4data_7;
    wire \scaler_4.N_1251_i_l_ofxZ0 ;
    wire \Commands_frame_decoder.source_offset4data_1_sqmuxa ;
    wire \Commands_frame_decoder.source_offset4data_1_sqmuxa_0 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_16 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_15 ;
    wire \pid_alt.m7_e_4_cascade_ ;
    wire \pid_alt.N_238_cascade_ ;
    wire \pid_alt.error_i_acumm_preregZ0Z_18 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_19 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_14 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_17 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_20 ;
    wire \uart_pc.timer_CountZ1Z_2 ;
    wire \uart_pc.un1_state_2_0_a3_0 ;
    wire \uart_pc.N_126_li_cascade_ ;
    wire \uart_pc.timer_Count_0_sqmuxa ;
    wire \uart_pc.timer_Count_RNO_0Z0Z_3 ;
    wire \uart_pc.timer_Count_0_sqmuxa_cascade_ ;
    wire \uart_pc.N_143 ;
    wire \uart_pc.N_145_cascade_ ;
    wire \uart_drone.data_Auxce_0_0_4 ;
    wire \uart_drone.data_Auxce_0_3 ;
    wire \uart_drone.data_Auxce_0_5 ;
    wire uart_pc_data_0;
    wire \Commands_frame_decoder.source_offset2data_1_sqmuxa_0 ;
    wire bfn_12_11_0_;
    wire frame_decoder_CH2data_1;
    wire frame_decoder_OFF2data_1;
    wire \scaler_2.un3_source_data_0_cry_0 ;
    wire frame_decoder_CH2data_2;
    wire frame_decoder_OFF2data_2;
    wire \scaler_2.un3_source_data_0_cry_1 ;
    wire frame_decoder_CH2data_3;
    wire frame_decoder_OFF2data_3;
    wire \scaler_2.un3_source_data_0_cry_2 ;
    wire frame_decoder_CH2data_4;
    wire frame_decoder_OFF2data_4;
    wire \scaler_2.un3_source_data_0_cry_3 ;
    wire frame_decoder_CH2data_5;
    wire frame_decoder_OFF2data_5;
    wire \scaler_2.un3_source_data_0_cry_4 ;
    wire frame_decoder_CH2data_6;
    wire frame_decoder_OFF2data_6;
    wire \scaler_2.un3_source_data_0_cry_5 ;
    wire \scaler_2.un3_source_data_0_axb_7 ;
    wire \scaler_2.un3_source_data_0_cry_6 ;
    wire \scaler_2.un3_source_data_0_cry_7 ;
    wire bfn_12_12_0_;
    wire \scaler_2.un3_source_data_0_cry_8 ;
    wire frame_decoder_OFF2data_7;
    wire frame_decoder_CH2data_7;
    wire \scaler_2.N_1227_i_l_ofxZ0 ;
    wire \pid_alt.pid_preregZ0Z_30 ;
    wire \pid_alt.N_106 ;
    wire \pid_alt.pid_preregZ0Z_9 ;
    wire \pid_alt.N_96_i_1 ;
    wire \pid_alt.un1_reset_0_i ;
    wire \scaler_3.un2_source_data_0_cry_1_c_RNO_0 ;
    wire bfn_12_14_0_;
    wire \scaler_3.un2_source_data_0_cry_1 ;
    wire \scaler_3.un3_source_data_0_cry_1_c_RNI44VK ;
    wire \scaler_3.un2_source_data_0_cry_2 ;
    wire \scaler_3.un3_source_data_0_cry_2_c_RNI780L ;
    wire \scaler_3.un2_source_data_0_cry_3 ;
    wire \scaler_3.un3_source_data_0_cry_3_c_RNIAC1L ;
    wire \scaler_3.un2_source_data_0_cry_4 ;
    wire \scaler_3.un3_source_data_0_cry_4_c_RNIDG2L ;
    wire \scaler_3.un2_source_data_0_cry_5 ;
    wire \scaler_3.un3_source_data_0_cry_5_c_RNIGK3L ;
    wire \scaler_3.un2_source_data_0_cry_6 ;
    wire \scaler_3.un3_source_data_0_cry_6_c_RNILUAN ;
    wire \scaler_3.un2_source_data_0_cry_7 ;
    wire \scaler_3.un2_source_data_0_cry_8 ;
    wire \scaler_3.un3_source_data_0_cry_7_c_RNIM0CN ;
    wire \scaler_3.un3_source_data_0_cry_8_c_RNIRV25 ;
    wire bfn_12_15_0_;
    wire \scaler_3.un2_source_data_0_cry_9 ;
    wire \scaler_4.un2_source_data_0_cry_1_c_RNO_1 ;
    wire bfn_12_16_0_;
    wire \scaler_4.un2_source_data_0_cry_1 ;
    wire \scaler_4.un3_source_data_0_cry_1_c_RNI74CL ;
    wire \scaler_4.un2_source_data_0_cry_2 ;
    wire \scaler_4.un3_source_data_0_cry_2_c_RNIA8DL ;
    wire \scaler_4.un2_source_data_0_cry_3 ;
    wire \scaler_4.un3_source_data_0_cry_3_c_RNIDCEL ;
    wire \scaler_4.un2_source_data_0_cry_4 ;
    wire \scaler_4.un3_source_data_0_cry_4_c_RNIGGFL ;
    wire \scaler_4.un2_source_data_0_cry_5 ;
    wire \scaler_4.un3_source_data_0_cry_5_c_RNIJKGL ;
    wire \scaler_4.un2_source_data_0_cry_6 ;
    wire \scaler_4.un3_source_data_0_cry_6_c_RNIOUNN ;
    wire \scaler_4.un2_source_data_0_cry_7 ;
    wire \scaler_4.un2_source_data_0_cry_8 ;
    wire \scaler_4.un3_source_data_0_cry_7_c_RNIP0PN ;
    wire \scaler_4.un3_source_data_0_cry_8_c_RNIS918 ;
    wire bfn_12_17_0_;
    wire \scaler_4.un2_source_data_0_cry_9 ;
    wire \pid_alt.un1_reset_1_0_i_cascade_ ;
    wire \pid_alt.error_i_acumm7lto4 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_2 ;
    wire \pid_alt.m21_e_8 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_3 ;
    wire \pid_alt.m21_e_2 ;
    wire \pid_alt.m21_e_10_cascade_ ;
    wire \pid_alt.N_138 ;
    wire \pid_alt.m35_e_3 ;
    wire \pid_alt.N_62_mux_cascade_ ;
    wire \pid_alt.N_129 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_1 ;
    wire \pid_alt.m21_e_0_cascade_ ;
    wire \pid_alt.m21_e_9 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_8 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_9 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_10 ;
    wire \pid_alt.m35_e_2 ;
    wire \pid_alt.N_62_mux ;
    wire \pid_alt.error_i_acumm7lto5 ;
    wire \pid_alt.error_i_acumm7lto12 ;
    wire \pid_alt.N_9_0 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_7 ;
    wire \uart_pc.N_144_1 ;
    wire \reset_module_System.count_1_1_cascade_ ;
    wire \uart_pc.data_AuxZ1Z_0 ;
    wire \uart_pc.data_AuxZ1Z_1 ;
    wire \uart_pc.data_AuxZ1Z_2 ;
    wire \uart_pc.data_AuxZ0Z_4 ;
    wire \uart_pc.data_AuxZ0Z_5 ;
    wire \uart_pc.data_AuxZ0Z_6 ;
    wire \uart_pc.un1_state_2_0 ;
    wire \uart_pc.data_AuxZ0Z_7 ;
    wire \uart_pc.state_RNIEAGSZ0Z_4 ;
    wire \uart_pc.data_Auxce_0_3 ;
    wire \uart_pc.data_Auxce_0_0_2 ;
    wire \uart_pc.data_Auxce_0_5 ;
    wire frame_decoder_OFF2data_0;
    wire frame_decoder_CH2data_0;
    wire \scaler_3.un2_source_data_0 ;
    wire frame_decoder_OFF3data_0;
    wire frame_decoder_CH3data_0;
    wire \scaler_4.un2_source_data_0 ;
    wire \uart_pc.data_Auxce_0_0_0 ;
    wire \uart_pc.data_Auxce_0_1 ;
    wire \uart_pc.data_Auxce_0_0_4 ;
    wire scaler_2_data_4;
    wire scaler_2_data_5;
    wire scaler_3_data_4;
    wire scaler_3_data_5;
    wire scaler_4_data_5;
    wire bfn_13_13_0_;
    wire \ppm_encoder_1.un1_throttle_cry_0 ;
    wire \ppm_encoder_1.un1_throttle_cry_1 ;
    wire \ppm_encoder_1.un1_throttle_cry_2 ;
    wire \ppm_encoder_1.un1_throttle_cry_3 ;
    wire throttle_command_5;
    wire \ppm_encoder_1.un1_throttle_cry_4_THRU_CO ;
    wire \ppm_encoder_1.un1_throttle_cry_4 ;
    wire \ppm_encoder_1.un1_throttle_cry_5 ;
    wire \ppm_encoder_1.un1_throttle_cry_6 ;
    wire \ppm_encoder_1.un1_throttle_cry_7 ;
    wire bfn_13_14_0_;
    wire \ppm_encoder_1.un1_throttle_cry_8 ;
    wire \ppm_encoder_1.un1_throttle_cry_9 ;
    wire \ppm_encoder_1.un1_throttle_cry_10 ;
    wire \ppm_encoder_1.un1_throttle_cry_11 ;
    wire \ppm_encoder_1.un1_throttle_cry_12 ;
    wire \ppm_encoder_1.un1_throttle_cry_13 ;
    wire throttle_command_2;
    wire \ppm_encoder_1.un1_throttle_cry_1_THRU_CO ;
    wire \ppm_encoder_1.un1_throttle_cry_0_THRU_CO ;
    wire throttle_command_1;
    wire \dron_frame_decoder_1.stateZ0Z_6 ;
    wire uart_drone_data_rdy;
    wire debug_CH1_0A_c;
    wire frame_decoder_OFF4data_0;
    wire frame_decoder_CH4data_0;
    wire scaler_4_data_4;
    wire ppm_output_c;
    wire throttle_command_10;
    wire \ppm_encoder_1.un1_throttle_cry_9_THRU_CO ;
    wire \ppm_encoder_1.un1_throttle_cry_3_THRU_CO ;
    wire throttle_command_4;
    wire scaler_4_data_6;
    wire bfn_13_17_0_;
    wire scaler_4_data_7;
    wire \ppm_encoder_1.un1_rudder_cry_6_THRU_CO ;
    wire \ppm_encoder_1.un1_rudder_cry_6 ;
    wire \ppm_encoder_1.un1_rudder_cry_7 ;
    wire scaler_4_data_9;
    wire \ppm_encoder_1.un1_rudder_cry_8_THRU_CO ;
    wire \ppm_encoder_1.un1_rudder_cry_8 ;
    wire \ppm_encoder_1.un1_rudder_cry_9 ;
    wire \ppm_encoder_1.un1_rudder_cry_10 ;
    wire \ppm_encoder_1.un1_rudder_cry_11 ;
    wire \ppm_encoder_1.un1_rudder_cry_12 ;
    wire \ppm_encoder_1.un1_rudder_cry_13 ;
    wire scaler_4_data_14;
    wire bfn_13_18_0_;
    wire bfn_13_19_0_;
    wire \ppm_encoder_1.un1_elevator_cry_6 ;
    wire scaler_3_data_8;
    wire \ppm_encoder_1.un1_elevator_cry_7_THRU_CO ;
    wire \ppm_encoder_1.un1_elevator_cry_7 ;
    wire \ppm_encoder_1.un1_elevator_cry_8 ;
    wire \ppm_encoder_1.un1_elevator_cry_9 ;
    wire \ppm_encoder_1.un1_elevator_cry_10 ;
    wire \ppm_encoder_1.un1_elevator_cry_11 ;
    wire \ppm_encoder_1.un1_elevator_cry_12 ;
    wire \ppm_encoder_1.un1_elevator_cry_13 ;
    wire scaler_3_data_14;
    wire bfn_13_20_0_;
    wire \pid_alt.un1_pid_prereg_0 ;
    wire bfn_13_21_0_;
    wire \pid_alt.error_i_acummZ0Z_1 ;
    wire \pid_alt.error_i_acumm_esr_RNIQMD91Z0Z_1 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_0 ;
    wire \pid_alt.error_i_acummZ0Z_2 ;
    wire \pid_alt.error_i_acumm_esr_RNITQE91Z0Z_2 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_1 ;
    wire \pid_alt.error_i_acummZ0Z_3 ;
    wire \pid_alt.error_i_acumm_esr_RNI0VF91Z0Z_3 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_2 ;
    wire \pid_alt.error_i_acummZ0Z_4 ;
    wire \pid_alt.error_i_acumm_esr_RNI33H91Z0Z_4 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_3 ;
    wire \pid_alt.error_i_acummZ0Z_5 ;
    wire \pid_alt.error_i_reg_esr_RNIT8KA1Z0Z_5 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_4 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_5_c_RNI0DLQ ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_5 ;
    wire \pid_alt.error_i_acummZ0Z_7 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_6_c_RNI3HMQ ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_6 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_7 ;
    wire \pid_alt.error_i_acummZ0Z_8 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_7_c_RNI6LNQ ;
    wire bfn_13_22_0_;
    wire \pid_alt.error_i_acummZ0Z_9 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_8_c_RNI9POQ ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_8 ;
    wire \pid_alt.error_i_acummZ0Z_10 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_9_c_RNIQN3F ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_9 ;
    wire \pid_alt.error_i_reg_esr_RNI4NMPZ0Z_11 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_10 ;
    wire \pid_alt.error_i_acummZ0Z_12 ;
    wire \pid_alt.error_i_reg_esr_RNI7RNPZ0Z_12 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_11 ;
    wire \pid_alt.error_i_acumm_esr_RNIJ6LMZ0Z_13 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_12 ;
    wire \pid_alt.error_i_reg_esr_RNI15KJZ0Z_14 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_13 ;
    wire \pid_alt.error_i_reg_esr_RNI38LJZ0Z_15 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_14 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_15 ;
    wire \pid_alt.error_i_reg_esr_RNI5BMJZ0Z_16 ;
    wire bfn_13_23_0_;
    wire \pid_alt.error_i_reg_esr_RNI7ENJZ0Z_17 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_16 ;
    wire \pid_alt.error_i_reg_esr_RNI9HOJZ0Z_18 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_17 ;
    wire \pid_alt.error_i_reg_esr_RNIBKPJZ0Z_19 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_18 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_19_c_RNI4FRJ ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_19 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_20 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_20_c_RNISVKK ;
    wire debug_CH3_20A_c;
    wire debug_CH3_20A_c_0;
    wire \uart_pc.N_126_li ;
    wire \uart_pc.state_srsts_0_0_0_cascade_ ;
    wire \uart_drone.state_srsts_0_0_0 ;
    wire \uart_pc.stateZ0Z_0 ;
    wire \uart_drone.N_126_li_cascade_ ;
    wire debug_CH2_18A_c;
    wire \uart_pc.state_srsts_i_0_2_cascade_ ;
    wire \uart_pc.stateZ0Z_1 ;
    wire \uart_pc.stateZ0Z_2 ;
    wire \uart_pc.timer_Count_RNILR1B2Z0Z_2 ;
    wire \uart_pc.data_AuxZ0Z_3 ;
    wire \uart_pc.timer_Count_RNIMQ8T1Z0Z_2 ;
    wire \uart_drone.stateZ0Z_0 ;
    wire \uart_drone.data_rdyc_1 ;
    wire \uart_pc.timer_CountZ1Z_3 ;
    wire \uart_pc.stateZ0Z_4 ;
    wire \uart_pc.timer_CountZ0Z_4 ;
    wire \uart_drone.N_126_li ;
    wire \uart_drone.un1_state_2_0 ;
    wire debug_CH0_16A_c;
    wire \uart_drone.state_srsts_i_0_2_cascade_ ;
    wire \uart_drone.stateZ0Z_1 ;
    wire \uart_drone.state_RNIOU0NZ0Z_4 ;
    wire \uart_pc.CO0_cascade_ ;
    wire \Commands_frame_decoder.un1_sink_data_valid_2_0 ;
    wire \Commands_frame_decoder.un1_sink_data_valid_2_0_0 ;
    wire \uart_pc.N_152 ;
    wire \uart_pc.un1_state_4_0 ;
    wire \uart_pc.N_152_cascade_ ;
    wire \uart_pc.stateZ0Z_3 ;
    wire \uart_pc.un1_state_7_0 ;
    wire \uart_pc.bit_CountZ0Z_0 ;
    wire \uart_pc.bit_CountZ0Z_1 ;
    wire \uart_pc.bit_CountZ0Z_2 ;
    wire \uart_pc.data_Auxce_0_6 ;
    wire \ppm_encoder_1.un2_throttle_iv_1_7_cascade_ ;
    wire \ppm_encoder_1.N_299_cascade_ ;
    wire \ppm_encoder_1.aileronZ0Z_7 ;
    wire \ppm_encoder_1.un1_elevator_cry_6_THRU_CO ;
    wire scaler_3_data_7;
    wire \ppm_encoder_1.elevatorZ0Z_7 ;
    wire \ppm_encoder_1.un1_throttle_cry_6_THRU_CO ;
    wire throttle_command_7;
    wire \scaler_2.un2_source_data_0_cry_1_c_RNOZ0 ;
    wire bfn_14_13_0_;
    wire \scaler_2.un2_source_data_0 ;
    wire \scaler_2.un2_source_data_0_cry_1 ;
    wire \scaler_2.un3_source_data_0_cry_1_c_RNI14IK ;
    wire \scaler_2.un2_source_data_0_cry_2 ;
    wire \scaler_2.un3_source_data_0_cry_2_c_RNI48JK ;
    wire \scaler_2.un2_source_data_0_cry_3 ;
    wire \scaler_2.un3_source_data_0_cry_3_c_RNI7CKK ;
    wire \scaler_2.un2_source_data_0_cry_4 ;
    wire \scaler_2.un3_source_data_0_cry_4_c_RNIAGLK ;
    wire \scaler_2.un2_source_data_0_cry_5 ;
    wire \scaler_2.un3_source_data_0_cry_5_c_RNIDKMK ;
    wire \scaler_2.un2_source_data_0_cry_6 ;
    wire \scaler_2.un3_source_data_0_cry_6_c_RNIIUTM ;
    wire \scaler_2.un2_source_data_0_cry_7 ;
    wire \scaler_2.un2_source_data_0_cry_8 ;
    wire \scaler_2.un3_source_data_0_cry_7_c_RNIJ0VM ;
    wire \scaler_2.un3_source_data_0_cry_8_c_RNIQL42 ;
    wire bfn_14_14_0_;
    wire \scaler_2.un2_source_data_0_cry_9 ;
    wire debug_CH3_20A_c_0_g;
    wire \ppm_encoder_1.un2_throttle_iv_0_9_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_1_9 ;
    wire \ppm_encoder_1.N_301_cascade_ ;
    wire \ppm_encoder_1.aileronZ0Z_9 ;
    wire scaler_3_data_9;
    wire \ppm_encoder_1.un1_elevator_cry_8_THRU_CO ;
    wire \ppm_encoder_1.elevatorZ0Z_9 ;
    wire throttle_command_9;
    wire \ppm_encoder_1.un1_throttle_cry_8_THRU_CO ;
    wire \ppm_encoder_1.throttleZ0Z_9 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_12_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_1_12 ;
    wire \ppm_encoder_1.aileronZ0Z_12 ;
    wire scaler_3_data_12;
    wire \ppm_encoder_1.un1_elevator_cry_11_THRU_CO ;
    wire throttle_command_12;
    wire \ppm_encoder_1.un1_throttle_cry_11_THRU_CO ;
    wire \ppm_encoder_1.un1_rudder_cry_10_THRU_CO ;
    wire scaler_4_data_11;
    wire throttle_command_11;
    wire \ppm_encoder_1.un1_throttle_cry_10_THRU_CO ;
    wire scaler_3_data_11;
    wire \ppm_encoder_1.un1_elevator_cry_10_THRU_CO ;
    wire scaler_4_data_12;
    wire \ppm_encoder_1.un1_rudder_cry_11_THRU_CO ;
    wire \ppm_encoder_1.rudderZ0Z_12 ;
    wire \ppm_encoder_1.N_320_cascade_ ;
    wire \ppm_encoder_1.throttleZ0Z_10 ;
    wire scaler_3_data_10;
    wire \ppm_encoder_1.un1_elevator_cry_9_THRU_CO ;
    wire \ppm_encoder_1.elevatorZ0Z_10 ;
    wire scaler_4_data_10;
    wire \ppm_encoder_1.un1_rudder_cry_9_THRU_CO ;
    wire reset_system;
    wire \ppm_encoder_1.counter24_0_I_57_c_RNIGCOZ0Z83 ;
    wire \ppm_encoder_1.N_145 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_21 ;
    wire \pid_alt.error_i_acumm7lto13 ;
    wire \pid_alt.N_238 ;
    wire \pid_alt.error_i_acummZ0Z_13 ;
    wire \pid_alt.N_96_i_0 ;
    wire uart_pc_data_6;
    wire alt_ki_6;
    wire \pid_alt.error_i_acumm_preregZ0Z_6 ;
    wire \pid_alt.error_i_acummZ0Z_6 ;
    wire \pid_alt.N_96_i ;
    wire \pid_alt.error_i_acumm_preregZ0Z_11 ;
    wire \pid_alt.N_128 ;
    wire \pid_alt.error_i_acummZ0Z_11 ;
    wire \pid_alt.un1_reset_1_0_i ;
    wire \pid_alt.error_i_acummZ0Z_0 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_0 ;
    wire \pid_alt.state_0_g_0 ;
    wire \uart_drone.un1_state_2_0_a3_0 ;
    wire bfn_15_6_0_;
    wire \uart_drone.timer_CountZ1Z_2 ;
    wire \uart_drone.timer_Count_RNO_0_0_2 ;
    wire \uart_drone.un4_timer_Count_1_cry_1 ;
    wire \uart_drone.timer_Count_RNO_0_0_3 ;
    wire \uart_drone.un4_timer_Count_1_cry_2 ;
    wire \uart_drone.un4_timer_Count_1_cry_3 ;
    wire \uart_drone.timer_Count_RNO_0_0_4 ;
    wire \reset_module_System.reset6_13_cascade_ ;
    wire \reset_module_System.reset6_3 ;
    wire \uart_drone.timer_CountZ0Z_0 ;
    wire \uart_drone.timer_Count_RNO_0_0_1_cascade_ ;
    wire \uart_drone.timer_CountZ1Z_1 ;
    wire \uart_drone.N_143 ;
    wire \uart_drone.timer_Count_0_sqmuxa ;
    wire \reset_module_System.reset6_15 ;
    wire \reset_module_System.reset6_17 ;
    wire \reset_module_System.reset6_19 ;
    wire \uart_drone.stateZ0Z_2 ;
    wire \uart_drone.N_145_cascade_ ;
    wire \uart_drone.data_Auxce_0_0_2 ;
    wire \uart_drone.data_Auxce_0_6 ;
    wire \ppm_encoder_1.throttleZ0Z_12 ;
    wire \ppm_encoder_1.elevatorZ0Z_12 ;
    wire \ppm_encoder_1.N_304 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_ns_2 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_ns_2_cascade_ ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_1 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_d_4_cascade_ ;
    wire \ppm_encoder_1.N_227_cascade_ ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1Z0Z_0_cascade_ ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_d_4 ;
    wire \ppm_encoder_1.un2_throttle_iv_1_1_cascade_ ;
    wire \ppm_encoder_1.elevatorZ0Z_4 ;
    wire \ppm_encoder_1.N_296_cascade_ ;
    wire \ppm_encoder_1.aileronZ0Z_4 ;
    wire \ppm_encoder_1.init_pulses_0_sqmuxa_0_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_1_6_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_0_6 ;
    wire \ppm_encoder_1.N_298_cascade_ ;
    wire \ppm_encoder_1.aileronZ0Z_6 ;
    wire scaler_3_data_6;
    wire \ppm_encoder_1.elevatorZ0Z_6 ;
    wire \ppm_encoder_1.un1_throttle_cry_5_THRU_CO ;
    wire throttle_command_6;
    wire \ppm_encoder_1.throttleZ0Z_6 ;
    wire \ppm_encoder_1.un2_throttle_iv_1_8_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_0_8 ;
    wire \ppm_encoder_1.elevatorZ0Z_8 ;
    wire throttle_command_8;
    wire \ppm_encoder_1.un1_throttle_cry_7_THRU_CO ;
    wire \ppm_encoder_1.throttleZ0Z_8 ;
    wire \ppm_encoder_1.un1_rudder_cry_7_THRU_CO ;
    wire scaler_4_data_8;
    wire \ppm_encoder_1.un2_throttle_iv_0_13_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_1_13 ;
    wire scaler_3_data_13;
    wire \ppm_encoder_1.un1_elevator_cry_12_THRU_CO ;
    wire throttle_command_13;
    wire \ppm_encoder_1.un1_throttle_cry_12_THRU_CO ;
    wire \ppm_encoder_1.throttleZ0Z_13 ;
    wire \ppm_encoder_1.elevatorZ0Z_13 ;
    wire \ppm_encoder_1.N_305_cascade_ ;
    wire \ppm_encoder_1.aileronZ0Z_13 ;
    wire \ppm_encoder_1.throttleZ0Z_11 ;
    wire \ppm_encoder_1.N_303_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_0_11 ;
    wire \ppm_encoder_1.rudderZ0Z_11 ;
    wire \ppm_encoder_1.N_319_cascade_ ;
    wire \ppm_encoder_1.throttleZ0Z_1 ;
    wire \ppm_encoder_1.N_302 ;
    wire \ppm_encoder_1.aileronZ0Z_10 ;
    wire \ppm_encoder_1.N_145_17 ;
    wire \ppm_encoder_1.N_145_17_cascade_ ;
    wire \ppm_encoder_1.N_238 ;
    wire \ppm_encoder_1.un1_PPM_STATE_1_sqmuxa_i_a3_0_1 ;
    wire \ppm_encoder_1.un2_throttle_iv_1_10 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_10 ;
    wire \ppm_encoder_1.PPM_STATEZ0Z_1 ;
    wire \ppm_encoder_1.PPM_STATE_ns_0_a3_0_1_0 ;
    wire \ppm_encoder_1.PPM_STATE_ns_0_a3_0_17_4_0 ;
    wire \ppm_encoder_1.PPM_STATE_ns_0_a3_0_17_3_0 ;
    wire \ppm_encoder_1.elevatorZ0Z_11 ;
    wire \ppm_encoder_1.un2_throttle_iv_1_11 ;
    wire \ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_5_0 ;
    wire \pid_alt.O_0_5 ;
    wire \pid_alt.error_i_regZ0Z_1 ;
    wire \reset_module_System.countZ0Z_1 ;
    wire \reset_module_System.countZ0Z_0 ;
    wire bfn_16_7_0_;
    wire \reset_module_System.countZ0Z_2 ;
    wire \reset_module_System.count_1_2 ;
    wire \reset_module_System.count_1_cry_1 ;
    wire \reset_module_System.countZ0Z_3 ;
    wire \reset_module_System.count_1_cry_2 ;
    wire \reset_module_System.countZ0Z_4 ;
    wire \reset_module_System.count_1_cry_3 ;
    wire \reset_module_System.countZ0Z_5 ;
    wire \reset_module_System.count_1_cry_4 ;
    wire \reset_module_System.countZ0Z_6 ;
    wire \reset_module_System.count_1_cry_5 ;
    wire \reset_module_System.countZ0Z_7 ;
    wire \reset_module_System.count_1_cry_6 ;
    wire \reset_module_System.countZ0Z_8 ;
    wire \reset_module_System.count_1_cry_7 ;
    wire \reset_module_System.count_1_cry_8 ;
    wire \reset_module_System.countZ0Z_9 ;
    wire bfn_16_8_0_;
    wire \reset_module_System.count_1_cry_9 ;
    wire \reset_module_System.count_1_cry_10 ;
    wire \reset_module_System.countZ0Z_12 ;
    wire \reset_module_System.count_1_cry_11 ;
    wire \reset_module_System.count_1_cry_12 ;
    wire \reset_module_System.count_1_cry_13 ;
    wire \reset_module_System.count_1_cry_14 ;
    wire \reset_module_System.countZ0Z_16 ;
    wire \reset_module_System.count_1_cry_15 ;
    wire \reset_module_System.count_1_cry_16 ;
    wire bfn_16_9_0_;
    wire \reset_module_System.countZ0Z_18 ;
    wire \reset_module_System.count_1_cry_17 ;
    wire \reset_module_System.count_1_cry_18 ;
    wire \reset_module_System.countZ0Z_20 ;
    wire \reset_module_System.count_1_cry_19 ;
    wire \reset_module_System.count_1_cry_20 ;
    wire \reset_module_System.countZ0Z_19 ;
    wire \reset_module_System.countZ0Z_15 ;
    wire \reset_module_System.countZ0Z_21 ;
    wire \reset_module_System.countZ0Z_13 ;
    wire \reset_module_System.reset6_11 ;
    wire \ppm_encoder_1.N_297_cascade_ ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_159_d_cascade_ ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_3 ;
    wire \ppm_encoder_1.pulses2count_9_sn_N_10_mux_cascade_ ;
    wire \ppm_encoder_1.throttleZ0Z_4 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_4_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_1_4 ;
    wire \ppm_encoder_1.throttleZ0Z_7 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_7 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2 ;
    wire \ppm_encoder_1.init_pulses_3_sqmuxa_0 ;
    wire \ppm_encoder_1.throttleZ0Z_5 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_ns_3 ;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_3_cascade_ ;
    wire \ppm_encoder_1.init_pulsesZ0Z_3 ;
    wire \ppm_encoder_1.pulses2count_9_sn_N_10_mux ;
    wire \ppm_encoder_1.un1_throttle_cry_2_THRU_CO ;
    wire throttle_command_3;
    wire \ppm_encoder_1.throttleZ0Z_3 ;
    wire \ppm_encoder_1.aileronZ0Z_5 ;
    wire \ppm_encoder_1.elevatorZ0Z_5 ;
    wire \ppm_encoder_1.un2_throttle_iv_1_5_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_0_5 ;
    wire \ppm_encoder_1.init_pulses_2_sqmuxa_0 ;
    wire \ppm_encoder_1.init_pulses_1_sqmuxa_0 ;
    wire \ppm_encoder_1.un2_throttle_iv_1_14_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_0_14 ;
    wire \ppm_encoder_1.throttleZ0Z_14 ;
    wire \ppm_encoder_1.elevatorZ0Z_14 ;
    wire scaler_2_data_6;
    wire bfn_16_15_0_;
    wire scaler_2_data_7;
    wire \ppm_encoder_1.un1_aileron_cry_6_THRU_CO ;
    wire \ppm_encoder_1.un1_aileron_cry_6 ;
    wire scaler_2_data_8;
    wire \ppm_encoder_1.un1_aileron_cry_7_THRU_CO ;
    wire \ppm_encoder_1.un1_aileron_cry_7 ;
    wire scaler_2_data_9;
    wire \ppm_encoder_1.un1_aileron_cry_8_THRU_CO ;
    wire \ppm_encoder_1.un1_aileron_cry_8 ;
    wire scaler_2_data_10;
    wire \ppm_encoder_1.un1_aileron_cry_9_THRU_CO ;
    wire \ppm_encoder_1.un1_aileron_cry_9 ;
    wire \ppm_encoder_1.un1_aileron_cry_10 ;
    wire scaler_2_data_12;
    wire \ppm_encoder_1.un1_aileron_cry_11_THRU_CO ;
    wire \ppm_encoder_1.un1_aileron_cry_11 ;
    wire scaler_2_data_13;
    wire \ppm_encoder_1.un1_aileron_cry_12_THRU_CO ;
    wire \ppm_encoder_1.un1_aileron_cry_12 ;
    wire \ppm_encoder_1.un1_aileron_cry_13 ;
    wire scaler_2_data_14;
    wire bfn_16_16_0_;
    wire \ppm_encoder_1.rudderZ0Z_10 ;
    wire scaler_4_data_13;
    wire \ppm_encoder_1.un1_rudder_cry_12_THRU_CO ;
    wire \ppm_encoder_1.pid_altitude_dv_0 ;
    wire \ppm_encoder_1.rudderZ0Z_6 ;
    wire scaler_2_data_11;
    wire \ppm_encoder_1.un1_aileron_cry_10_THRU_CO ;
    wire \ppm_encoder_1.aileronZ0Z_11 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_4 ;
    wire \ppm_encoder_1.pulses2countZ0Z_4 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_5 ;
    wire \ppm_encoder_1.pulses2countZ0Z_5 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_0 ;
    wire \ppm_encoder_1.pulses2countZ0Z_0 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_1 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_1 ;
    wire \ppm_encoder_1.pulses2countZ0Z_1 ;
    wire \ppm_encoder_1.N_1330_i ;
    wire \ppm_encoder_1.counterZ0Z_0 ;
    wire bfn_16_19_0_;
    wire \ppm_encoder_1.counterZ0Z_1 ;
    wire \ppm_encoder_1.un1_counter_13_cry_0 ;
    wire \ppm_encoder_1.un1_counter_13_cry_1 ;
    wire \ppm_encoder_1.un1_counter_13_cry_2 ;
    wire \ppm_encoder_1.counterZ0Z_4 ;
    wire \ppm_encoder_1.un1_counter_13_cry_3 ;
    wire \ppm_encoder_1.counterZ0Z_5 ;
    wire \ppm_encoder_1.un1_counter_13_cry_4 ;
    wire \ppm_encoder_1.un1_counter_13_cry_5 ;
    wire \ppm_encoder_1.un1_counter_13_cry_6 ;
    wire \ppm_encoder_1.un1_counter_13_cry_7 ;
    wire bfn_16_20_0_;
    wire \ppm_encoder_1.un1_counter_13_cry_8 ;
    wire \ppm_encoder_1.un1_counter_13_cry_9 ;
    wire \ppm_encoder_1.un1_counter_13_cry_10 ;
    wire \ppm_encoder_1.un1_counter_13_cry_11 ;
    wire \ppm_encoder_1.un1_counter_13_cry_12 ;
    wire \ppm_encoder_1.un1_counter_13_cry_13 ;
    wire \ppm_encoder_1.un1_counter_13_cry_14 ;
    wire \ppm_encoder_1.un1_counter_13_cry_15 ;
    wire bfn_16_21_0_;
    wire \ppm_encoder_1.un1_counter_13_cry_16 ;
    wire \ppm_encoder_1.un1_counter_13_cry_17 ;
    wire \ppm_encoder_1.N_322_g ;
    wire uart_pc_data_2;
    wire alt_ki_2;
    wire \pid_alt.O_0_6 ;
    wire \pid_alt.error_i_regZ0Z_2 ;
    wire \uart_drone.N_144_1 ;
    wire \uart_drone.bit_CountZ0Z_2 ;
    wire \uart_drone.timer_CountZ0Z_4 ;
    wire \uart_drone.timer_CountZ1Z_3 ;
    wire \uart_drone.stateZ0Z_4 ;
    wire \uart_drone.un1_state_4_0_cascade_ ;
    wire \reset_module_System.countZ0Z_11 ;
    wire \reset_module_System.countZ0Z_14 ;
    wire \reset_module_System.countZ0Z_17 ;
    wire \reset_module_System.countZ0Z_10 ;
    wire \reset_module_System.reset6_14 ;
    wire \ppm_encoder_1.un1_init_pulses_10_0 ;
    wire \ppm_encoder_1.un1_init_pulses_11_0_cascade_ ;
    wire \ppm_encoder_1.un1_init_pulses_0_cascade_ ;
    wire pid_altitude_dv;
    wire throttle_command_0;
    wire \ppm_encoder_1.throttleZ0Z_0 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_0 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_0 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_4 ;
    wire \ppm_encoder_1.rudderZ0Z_4 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_4 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_5 ;
    wire \ppm_encoder_1.rudderZ0Z_5 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_5 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_1 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_11 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_12 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1Z0Z_0 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_2 ;
    wire \ppm_encoder_1.throttleZ0Z_2 ;
    wire \ppm_encoder_1.init_pulses_0_sqmuxa_0 ;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_2_cascade_ ;
    wire \ppm_encoder_1.init_pulsesZ0Z_6 ;
    wire \ppm_encoder_1.throttle_RNIN3352Z0Z_0 ;
    wire \ppm_encoder_1.un1_init_pulses_0 ;
    wire bfn_17_14_0_;
    wire \ppm_encoder_1.throttle_RNIALN65Z0Z_1 ;
    wire \ppm_encoder_1.un1_init_pulses_0_1 ;
    wire \ppm_encoder_1.un1_init_pulses_10_1 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_0 ;
    wire \ppm_encoder_1.throttle_RNI5V123Z0Z_2 ;
    wire \ppm_encoder_1.un1_init_pulses_0_2 ;
    wire \ppm_encoder_1.un1_init_pulses_10_2 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_1 ;
    wire \ppm_encoder_1.throttle_RNI82223Z0Z_3 ;
    wire \ppm_encoder_1.un1_init_pulses_0_3 ;
    wire \ppm_encoder_1.un1_init_pulses_10_3 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_2 ;
    wire \ppm_encoder_1.aileron_esr_RNIV9IN5Z0Z_4 ;
    wire \ppm_encoder_1.un1_init_pulses_0_4 ;
    wire \ppm_encoder_1.un1_init_pulses_10_4 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_3 ;
    wire \ppm_encoder_1.aileron_esr_RNI4FIN5Z0Z_5 ;
    wire \ppm_encoder_1.un1_init_pulses_0_5 ;
    wire \ppm_encoder_1.un1_init_pulses_10_5 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_4 ;
    wire \ppm_encoder_1.throttle_RNIEDI96Z0Z_6 ;
    wire \ppm_encoder_1.un1_init_pulses_0_6 ;
    wire \ppm_encoder_1.un1_init_pulses_10_6 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_5 ;
    wire \ppm_encoder_1.throttle_RNIJII96Z0Z_7 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_6 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_7 ;
    wire \ppm_encoder_1.throttle_RNIONI96Z0Z_8 ;
    wire bfn_17_15_0_;
    wire \ppm_encoder_1.throttle_RNITSI96Z0Z_9 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_8 ;
    wire \ppm_encoder_1.elevator_RNI5GRT5Z0Z_10 ;
    wire \ppm_encoder_1.un1_init_pulses_10_10 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_9 ;
    wire \ppm_encoder_1.elevator_RNIALRT5Z0Z_11 ;
    wire \ppm_encoder_1.un1_init_pulses_0_11 ;
    wire \ppm_encoder_1.un1_init_pulses_10_11 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_10 ;
    wire \ppm_encoder_1.elevator_RNIFQRT5Z0Z_12 ;
    wire \ppm_encoder_1.un1_init_pulses_0_12 ;
    wire \ppm_encoder_1.un1_init_pulses_10_12 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_11 ;
    wire \ppm_encoder_1.elevator_RNIKVRT5Z0Z_13 ;
    wire \ppm_encoder_1.un1_init_pulses_0_13 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_12 ;
    wire \ppm_encoder_1.aileron_esr_RNITH3L6Z0Z_14 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_13 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI7O1NZ0Z_2 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_14 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_15 ;
    wire bfn_17_16_0_;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_17 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_16 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_17 ;
    wire \ppm_encoder_1.rudderZ0Z_8 ;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_16 ;
    wire \ppm_encoder_1.aileronZ0Z_14 ;
    wire \ppm_encoder_1.N_306 ;
    wire \pid_alt.un9_error_filt_1_15 ;
    wire \pid_alt.un9_error_filt_2_0 ;
    wire \pid_alt.un9_error_filt_add_1_axbZ0Z_0 ;
    wire bfn_17_17_0_;
    wire \pid_alt.un9_error_filt_1_16 ;
    wire \pid_alt.un9_error_filt_2_1 ;
    wire \pid_alt.un9_error_filt_add_1_cry_1_sZ0 ;
    wire \pid_alt.un9_error_filt_add_1_cry_0 ;
    wire \pid_alt.un9_error_filt_1_17 ;
    wire \pid_alt.un9_error_filt_2_2 ;
    wire \pid_alt.un9_error_filt_add_1_cry_2_sZ0 ;
    wire \pid_alt.un9_error_filt_add_1_cry_1 ;
    wire \pid_alt.un9_error_filt_1_18 ;
    wire \pid_alt.un9_error_filt_2_3 ;
    wire \pid_alt.un9_error_filt_add_1_cry_3_sZ0 ;
    wire \pid_alt.un9_error_filt_add_1_cry_2 ;
    wire \pid_alt.un9_error_filt_2_4 ;
    wire \pid_alt.un9_error_filt_add_1_cry_4_sZ0 ;
    wire \pid_alt.un9_error_filt_add_1_cry_3 ;
    wire \pid_alt.un9_error_filt_2_5 ;
    wire \pid_alt.un9_error_filt_add_1_cry_5_sZ0 ;
    wire \pid_alt.un9_error_filt_add_1_cry_4 ;
    wire \pid_alt.un9_error_filt_2_6 ;
    wire \pid_alt.un9_error_filt_add_1_cry_6_sZ0 ;
    wire \pid_alt.un9_error_filt_add_1_cry_5 ;
    wire \pid_alt.un9_error_filt_2_7 ;
    wire \pid_alt.un9_error_filt_add_1_cry_7_sZ0 ;
    wire \pid_alt.un9_error_filt_add_1_cry_6 ;
    wire \pid_alt.un9_error_filt_add_1_cry_7 ;
    wire \pid_alt.un9_error_filt_2_8 ;
    wire \pid_alt.un9_error_filt_add_1_cry_8_sZ0 ;
    wire bfn_17_18_0_;
    wire \pid_alt.un9_error_filt_2_9 ;
    wire \pid_alt.un9_error_filt_add_1_cry_9_sZ0 ;
    wire \pid_alt.un9_error_filt_add_1_cry_8 ;
    wire \pid_alt.un9_error_filt_2_10 ;
    wire \pid_alt.un9_error_filt_add_1_cry_10_sZ0 ;
    wire \pid_alt.un9_error_filt_add_1_cry_9 ;
    wire \pid_alt.un9_error_filt_1_19 ;
    wire \pid_alt.un9_error_filt_2_11 ;
    wire \pid_alt.un9_error_filt_add_1_cry_10 ;
    wire \pid_alt.un9_error_filt_add_1_sZ0Z_11 ;
    wire \ppm_encoder_1.N_140_0 ;
    wire \ppm_encoder_1.un1_init_pulses_0_10 ;
    wire \ppm_encoder_1.rudderZ0Z_13 ;
    wire \ppm_encoder_1.CHOOSE_CHANNELZ0Z_0 ;
    wire \ppm_encoder_1.N_300 ;
    wire \ppm_encoder_1.aileronZ0Z_8 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_8_cascade_ ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_8 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_9 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_13 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_13 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_2 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_2 ;
    wire \ppm_encoder_1.counterZ0Z_3 ;
    wire \ppm_encoder_1.pulses2countZ0Z_2 ;
    wire \ppm_encoder_1.counterZ0Z_2 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_3 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_3 ;
    wire \ppm_encoder_1.pulses2countZ0Z_3 ;
    wire \ppm_encoder_1.pulses2countZ0Z_8 ;
    wire \ppm_encoder_1.counterZ0Z_9 ;
    wire \ppm_encoder_1.pulses2countZ0Z_9 ;
    wire \ppm_encoder_1.counterZ0Z_8 ;
    wire \ppm_encoder_1.counterZ0Z_14 ;
    wire \ppm_encoder_1.pulses2countZ0Z_15 ;
    wire \ppm_encoder_1.pulses2countZ0Z_16 ;
    wire \ppm_encoder_1.pulses2countZ0Z_17 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_159_d ;
    wire \ppm_encoder_1.counterZ0Z_15 ;
    wire \ppm_encoder_1.counterZ0Z_17 ;
    wire \ppm_encoder_1.counterZ0Z_16 ;
    wire \ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_4_0 ;
    wire \ppm_encoder_1.pulses2countZ0Z_18 ;
    wire \ppm_encoder_1.counterZ0Z_18 ;
    wire \pid_alt.O_0_4 ;
    wire \pid_alt.error_i_regZ0Z_0 ;
    wire \pid_alt.O_0_7 ;
    wire \pid_alt.error_i_regZ0Z_3 ;
    wire \uart_drone.CO0 ;
    wire \uart_drone.un1_state_7_0 ;
    wire \uart_drone.bit_CountZ0Z_1 ;
    wire \ppm_encoder_1.CHOOSE_CHANNELZ0Z_1 ;
    wire \ppm_encoder_1.CHOOSE_CHANNELZ0Z_3 ;
    wire \ppm_encoder_1.PPM_STATE_RNI2APU1_2Z0Z_1 ;
    wire \ppm_encoder_1.init_pulses_RNIAVNR2Z0Z_0 ;
    wire bfn_18_11_0_;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_1 ;
    wire \ppm_encoder_1.un1_init_pulses_11_1 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_0 ;
    wire \ppm_encoder_1.PPM_STATE_RNI2APU1_1Z0Z_1 ;
    wire \ppm_encoder_1.init_pulses_RNIC1OR2Z0Z_2 ;
    wire \ppm_encoder_1.un1_init_pulses_11_2 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_1 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_3 ;
    wire \ppm_encoder_1.un1_init_pulses_11_3 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_2 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_4 ;
    wire \ppm_encoder_1.un1_init_pulses_11_4 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_3 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_5 ;
    wire \ppm_encoder_1.un1_init_pulses_11_5 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_4 ;
    wire \ppm_encoder_1.PPM_STATE_RNI2APU1_0Z0Z_1 ;
    wire \ppm_encoder_1.init_pulses_RNIG5OR2Z0Z_6 ;
    wire \ppm_encoder_1.un1_init_pulses_11_6 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_5 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_6 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_7 ;
    wire bfn_18_12_0_;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_8 ;
    wire \ppm_encoder_1.un1_init_pulses_11_10 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_9 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_11 ;
    wire \ppm_encoder_1.un1_init_pulses_11_11 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_10 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_12 ;
    wire \ppm_encoder_1.un1_init_pulses_11_12 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_11 ;
    wire \ppm_encoder_1.init_pulses_RNIUPKO2Z0Z_13 ;
    wire \ppm_encoder_1.PPM_STATE_RNI2APU1Z0Z_1 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_12 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_13 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_14 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_15 ;
    wire bfn_18_13_0_;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_16 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_17 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1 ;
    wire \ppm_encoder_1.N_227 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1 ;
    wire \ppm_encoder_1.PPM_STATEZ0Z_0 ;
    wire \ppm_encoder_1.init_pulses_0_sqmuxa_1_0_cascade_ ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_8 ;
    wire \ppm_encoder_1.un1_init_pulses_11_7 ;
    wire \ppm_encoder_1.un1_init_pulses_10_7 ;
    wire \ppm_encoder_1.un1_init_pulses_0_7 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_7 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_7 ;
    wire \ppm_encoder_1.rudderZ0Z_7 ;
    wire \ppm_encoder_1.un1_init_pulses_11_8 ;
    wire \ppm_encoder_1.un1_init_pulses_10_8 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_8 ;
    wire \ppm_encoder_1.un1_init_pulses_0_8 ;
    wire \ppm_encoder_1.un1_init_pulses_10_9 ;
    wire \ppm_encoder_1.un1_init_pulses_11_9 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_9 ;
    wire \ppm_encoder_1.un1_init_pulses_0_9 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_9 ;
    wire \ppm_encoder_1.rudderZ0Z_9 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_9 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_17 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_10 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_10 ;
    wire \ppm_encoder_1.un1_init_pulses_11_14 ;
    wire \ppm_encoder_1.un1_init_pulses_10_14 ;
    wire \ppm_encoder_1.un1_init_pulses_0_14 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_14 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_14 ;
    wire \ppm_encoder_1.pulses2count_9_sn_N_7 ;
    wire \ppm_encoder_1.rudderZ0Z_14 ;
    wire \ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ;
    wire \ppm_encoder_1.un1_init_pulses_11_16 ;
    wire \ppm_encoder_1.un1_init_pulses_10_16 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_16 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_16 ;
    wire \ppm_encoder_1.un1_init_pulses_11_17 ;
    wire \ppm_encoder_1.un1_init_pulses_10_17 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_17 ;
    wire \ppm_encoder_1.init_pulses_RNI5ATG1Z0Z_15 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_15 ;
    wire \ppm_encoder_1.un1_init_pulses_11_15 ;
    wire \ppm_encoder_1.un1_init_pulses_10_15 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_15 ;
    wire \ppm_encoder_1.un1_init_pulses_0Z0Z_1 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_d_12 ;
    wire \ppm_encoder_1.PPM_STATE_59_d ;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_18 ;
    wire \ppm_encoder_1.un1_init_pulses_11_18 ;
    wire \ppm_encoder_1.un1_init_pulses_10_18 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_18 ;
    wire \ppm_encoder_1.init_pulses_0_sqmuxa_1 ;
    wire \ppm_encoder_1.un1_init_pulses_11_13 ;
    wire \ppm_encoder_1.un1_init_pulses_4_sqmuxa_0 ;
    wire \ppm_encoder_1.un1_init_pulses_10_13 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_13 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_14 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_14 ;
    wire \ppm_encoder_1.pulses2countZ0Z_14 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_10 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_10 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_7 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_7 ;
    wire \ppm_encoder_1.counterZ0Z_7 ;
    wire \ppm_encoder_1.pulses2countZ0Z_7 ;
    wire \ppm_encoder_1.counterZ0Z_6 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_6 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_6 ;
    wire \ppm_encoder_1.pulses2countZ0Z_6 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_11 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_11 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_12 ;
    wire \ppm_encoder_1.pulses2count_9_sn_N_11_mux ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_12 ;
    wire \ppm_encoder_1.N_1330_0 ;
    wire \ppm_encoder_1.counterZ0Z_13 ;
    wire \ppm_encoder_1.pulses2countZ0Z_12 ;
    wire \ppm_encoder_1.pulses2countZ0Z_13 ;
    wire \ppm_encoder_1.counterZ0Z_12 ;
    wire \ppm_encoder_1.counter24_0_I_1_c_RNOZ0 ;
    wire bfn_18_20_0_;
    wire \ppm_encoder_1.counter24_0_I_9_c_RNOZ0 ;
    wire \ppm_encoder_1.counter24_0_data_tmp_0 ;
    wire \ppm_encoder_1.counter24_0_I_15_c_RNOZ0 ;
    wire \ppm_encoder_1.counter24_0_data_tmp_1 ;
    wire \ppm_encoder_1.counter24_0_I_21_c_RNOZ0 ;
    wire \ppm_encoder_1.counter24_0_data_tmp_2 ;
    wire \ppm_encoder_1.counter24_0_I_27_c_RNOZ0 ;
    wire \ppm_encoder_1.counter24_0_data_tmp_3 ;
    wire \ppm_encoder_1.counter24_0_data_tmp_4 ;
    wire \ppm_encoder_1.counter24_0_I_39_c_RNOZ0 ;
    wire \ppm_encoder_1.counter24_0_data_tmp_5 ;
    wire \ppm_encoder_1.counter24_0_I_45_c_RNOZ0 ;
    wire \ppm_encoder_1.counter24_0_data_tmp_6 ;
    wire \ppm_encoder_1.counter24_0_data_tmp_7 ;
    wire \ppm_encoder_1.counter24_0_I_51_c_RNOZ0 ;
    wire bfn_18_21_0_;
    wire CONSTANT_ONE_NET;
    wire \ppm_encoder_1.counter24_0_I_57_c_RNOZ0 ;
    wire \ppm_encoder_1.counter24_0_data_tmp_8 ;
    wire \ppm_encoder_1.counter24_0_N_2 ;
    wire \ppm_encoder_1.counter24_0_N_2_THRU_CO ;
    wire \ppm_encoder_1.pulses2countZ0Z_10 ;
    wire \ppm_encoder_1.counterZ0Z_11 ;
    wire \ppm_encoder_1.pulses2countZ0Z_11 ;
    wire \ppm_encoder_1.counterZ0Z_10 ;
    wire \ppm_encoder_1.counter24_0_I_33_c_RNOZ0 ;
    wire \uart_drone.stateZ0Z_3 ;
    wire \uart_drone.un1_state_4_0 ;
    wire \uart_drone.N_152 ;
    wire \uart_drone.bit_CountZ0Z_0 ;
    wire \pid_alt.error_filt_21 ;
    wire \pid_alt.error_filt_prevZ0Z_21 ;
    wire uart_pc_data_5;
    wire alt_ki_5;
    wire reset_system_g;
    wire GB_BUFFER_reset_system_g_THRU_CO;
    wire uart_pc_data_3;
    wire alt_ki_3;
    wire \pid_alt.O_0_8 ;
    wire \pid_alt.error_i_regZ0Z_4 ;
    wire \pid_alt.O_0_9 ;
    wire \pid_alt.error_i_regZ0Z_5 ;
    wire \pid_alt.O_0_12 ;
    wire \pid_alt.error_i_regZ0Z_8 ;
    wire uart_pc_data_4;
    wire alt_ki_4;
    wire uart_pc_data_1;
    wire alt_ki_1;
    wire \pid_alt.error_filt_19 ;
    wire \pid_alt.error_filt_prevZ0Z_19 ;
    wire uart_pc_data_7;
    wire alt_ki_7;
    wire \Commands_frame_decoder.state_RNIQRI31Z0Z_10 ;
    wire \pid_alt.O_0_14 ;
    wire \pid_alt.error_i_regZ0Z_10 ;
    wire \pid_alt.O_15 ;
    wire \pid_alt.error_i_regZ0Z_11 ;
    wire \pid_alt.O_16 ;
    wire \pid_alt.error_i_regZ0Z_12 ;
    wire \pid_alt.O_17 ;
    wire \pid_alt.error_i_regZ0Z_13 ;
    wire \pid_alt.error_filt_17 ;
    wire \pid_alt.error_filt_prevZ0Z_17 ;
    wire \pid_alt.error_filt_18 ;
    wire \pid_alt.error_filt_prevZ0Z_18 ;
    wire \pid_alt.error_filt_22 ;
    wire \pid_alt.error_filt_prevZ0Z_22 ;
    wire \pid_alt.error_filt_20 ;
    wire \pid_alt.error_filt_prevZ0Z_20 ;
    wire \pid_alt.error_filt_8 ;
    wire \pid_alt.error_filt_prevZ0Z_8 ;
    wire \pid_alt.O_8 ;
    wire \pid_alt.error_d_regZ0Z_4 ;
    wire \pid_alt.error_filt_1 ;
    wire \pid_alt.error_filt_prevZ0Z_1 ;
    wire \pid_alt.error_filt_2 ;
    wire \pid_alt.error_filt_prevZ0Z_2 ;
    wire \pid_alt.error_filt_10 ;
    wire \pid_alt.error_filt_prevZ0Z_10 ;
    wire \pid_alt.error_filt_11 ;
    wire \pid_alt.error_filt_prevZ0Z_11 ;
    wire \pid_alt.error_filt_12 ;
    wire \pid_alt.error_filt_prevZ0Z_12 ;
    wire \pid_alt.error_filt_13 ;
    wire \pid_alt.error_filt_prevZ0Z_13 ;
    wire \pid_alt.error_filt_15 ;
    wire \pid_alt.error_filt_prevZ0Z_15 ;
    wire \pid_alt.error_filt_16 ;
    wire \pid_alt.error_filt_prevZ0Z_16 ;
    wire \pid_alt.error_filt_4 ;
    wire \pid_alt.error_filt_prevZ0Z_4 ;
    wire \pid_alt.error_filt_5 ;
    wire \pid_alt.error_filt_prevZ0Z_5 ;
    wire \pid_alt.error_filt_6 ;
    wire \pid_alt.error_filt_prevZ0Z_6 ;
    wire \pid_alt.error_filt_7 ;
    wire \pid_alt.error_filt_prevZ0Z_7 ;
    wire \pid_alt.error_filt_9 ;
    wire \pid_alt.error_filt_prevZ0Z_9 ;
    wire \pid_alt.error_filt_3 ;
    wire \pid_alt.error_filt_prevZ0Z_3 ;
    wire \pid_alt.error_filt_14 ;
    wire \pid_alt.error_filt_prevZ0Z_14 ;
    wire \pid_alt.O_0_11 ;
    wire \pid_alt.error_i_regZ0Z_7 ;
    wire \pid_alt.O_0_10 ;
    wire \pid_alt.error_i_regZ0Z_6 ;
    wire \pid_alt.O_19 ;
    wire \pid_alt.error_i_regZ0Z_15 ;
    wire \pid_alt.O_0_13 ;
    wire \pid_alt.error_i_regZ0Z_9 ;
    wire \pid_alt.O_18 ;
    wire \pid_alt.error_i_regZ0Z_14 ;
    wire \pid_alt.O_24 ;
    wire \pid_alt.error_i_regZ0Z_20 ;
    wire \pid_alt.O_21 ;
    wire \pid_alt.error_i_regZ0Z_17 ;
    wire \pid_alt.O_22 ;
    wire \pid_alt.error_i_regZ0Z_18 ;
    wire \pid_alt.O_20 ;
    wire \pid_alt.error_i_regZ0Z_16 ;
    wire \pid_alt.O_23 ;
    wire \pid_alt.error_i_regZ0Z_19 ;
    wire _gnd_net_;
    wire clk_system_c_g;
    wire \pid_alt.N_410_0_g ;
    wire N_411_g;

    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .A_REG=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .NEG_TRIGGER=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .MODE_8x8=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .D_REG=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .C_REG=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .B_SIGNED=1'b1;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .B_REG=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .A_SIGNED=1'b1;
    SB_MAC16 \pid_alt.un2_error_1_mulonly_0_24_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__43117),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__43116),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_0,dangling_wire_1,dangling_wire_2,dangling_wire_3,dangling_wire_4,dangling_wire_5,dangling_wire_6,dangling_wire_7,dangling_wire_8,dangling_wire_9,dangling_wire_10,dangling_wire_11,dangling_wire_12,dangling_wire_13,dangling_wire_14,dangling_wire_15}),
            .ADDSUBBOT(),
            .A({N__22139,N__22196,N__22243,N__21569,N__21616,N__21672,N__21716,N__21770,N__21830,N__21889,N__21953,N__21329,N__21379,N__21435,N__21485,N__24458}),
            .C({dangling_wire_16,dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21,dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27,dangling_wire_28,dangling_wire_29,dangling_wire_30,dangling_wire_31}),
            .B({dangling_wire_32,dangling_wire_33,dangling_wire_34,dangling_wire_35,dangling_wire_36,dangling_wire_37,dangling_wire_38,dangling_wire_39,N__18534,N__19032,N__19020,N__25506,N__18561,N__18777,N__18546,N__19047}),
            .OHOLDTOP(),
            .O({dangling_wire_40,dangling_wire_41,dangling_wire_42,dangling_wire_43,dangling_wire_44,dangling_wire_45,dangling_wire_46,\pid_alt.O_0_24 ,\pid_alt.O_0_23 ,\pid_alt.O_0_22 ,\pid_alt.O_0_21 ,\pid_alt.O_0_20 ,\pid_alt.O_0_19 ,\pid_alt.O_0_18 ,\pid_alt.O_0_17 ,\pid_alt.O_0_16 ,\pid_alt.O_0_15 ,\pid_alt.O_1_14 ,\pid_alt.O_1_13 ,\pid_alt.O_1_12 ,\pid_alt.O_1_11 ,\pid_alt.O_1_10 ,\pid_alt.O_1_9 ,\pid_alt.O_1_8 ,\pid_alt.O_1_7 ,\pid_alt.O_1_6 ,\pid_alt.O_1_5 ,\pid_alt.O_1_4 ,dangling_wire_47,dangling_wire_48,dangling_wire_49,dangling_wire_50}));
    defparam \pid_alt.un9_error_filt_1_mulonly_0_19_0 .A_REG=1'b0;
    defparam \pid_alt.un9_error_filt_1_mulonly_0_19_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pid_alt.un9_error_filt_1_mulonly_0_19_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pid_alt.un9_error_filt_1_mulonly_0_19_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pid_alt.un9_error_filt_1_mulonly_0_19_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pid_alt.un9_error_filt_1_mulonly_0_19_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pid_alt.un9_error_filt_1_mulonly_0_19_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pid_alt.un9_error_filt_1_mulonly_0_19_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pid_alt.un9_error_filt_1_mulonly_0_19_0 .NEG_TRIGGER=1'b0;
    defparam \pid_alt.un9_error_filt_1_mulonly_0_19_0 .MODE_8x8=1'b0;
    defparam \pid_alt.un9_error_filt_1_mulonly_0_19_0 .D_REG=1'b0;
    defparam \pid_alt.un9_error_filt_1_mulonly_0_19_0 .C_REG=1'b0;
    defparam \pid_alt.un9_error_filt_1_mulonly_0_19_0 .B_SIGNED=1'b1;
    defparam \pid_alt.un9_error_filt_1_mulonly_0_19_0 .B_REG=1'b0;
    defparam \pid_alt.un9_error_filt_1_mulonly_0_19_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pid_alt.un9_error_filt_1_mulonly_0_19_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pid_alt.un9_error_filt_1_mulonly_0_19_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pid_alt.un9_error_filt_1_mulonly_0_19_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pid_alt.un9_error_filt_1_mulonly_0_19_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pid_alt.un9_error_filt_1_mulonly_0_19_0 .A_SIGNED=1'b1;
    SB_MAC16 \pid_alt.un9_error_filt_1_mulonly_0_19_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__43130),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__43085),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_51,dangling_wire_52,dangling_wire_53,dangling_wire_54,dangling_wire_55,dangling_wire_56,dangling_wire_57,dangling_wire_58,dangling_wire_59,dangling_wire_60,dangling_wire_61,dangling_wire_62,dangling_wire_63,dangling_wire_64,dangling_wire_65,dangling_wire_66}),
            .ADDSUBBOT(),
            .A({dangling_wire_67,N__46254,N__45996,N__46032,N__46071,N__46113,N__46320,N__45534,N__46365,N__46398,N__45837,N__45870,N__46287,N__46149,N__45429,N__17958}),
            .C({dangling_wire_68,dangling_wire_69,dangling_wire_70,dangling_wire_71,dangling_wire_72,dangling_wire_73,dangling_wire_74,dangling_wire_75,dangling_wire_76,dangling_wire_77,dangling_wire_78,dangling_wire_79,dangling_wire_80,dangling_wire_81,dangling_wire_82,dangling_wire_83}),
            .B({dangling_wire_84,dangling_wire_85,dangling_wire_86,dangling_wire_87,dangling_wire_88,dangling_wire_89,dangling_wire_90,dangling_wire_91,dangling_wire_92,dangling_wire_93,dangling_wire_94,dangling_wire_95,dangling_wire_96,N__43087,N__43129,N__43086}),
            .OHOLDTOP(),
            .O({dangling_wire_97,dangling_wire_98,dangling_wire_99,dangling_wire_100,dangling_wire_101,dangling_wire_102,dangling_wire_103,dangling_wire_104,dangling_wire_105,dangling_wire_106,dangling_wire_107,dangling_wire_108,\pid_alt.un9_error_filt_1_19 ,\pid_alt.un9_error_filt_1_18 ,\pid_alt.un9_error_filt_1_17 ,\pid_alt.un9_error_filt_1_16 ,\pid_alt.un9_error_filt_1_15 ,\pid_alt.O_3_14 ,\pid_alt.O_3_13 ,\pid_alt.O_3_12 ,\pid_alt.O_3_11 ,\pid_alt.O_3_10 ,\pid_alt.O_3_9 ,\pid_alt.O_3_8 ,\pid_alt.O_3_7 ,\pid_alt.O_3_6 ,\pid_alt.error_filt ,dangling_wire_109,dangling_wire_110,dangling_wire_111,dangling_wire_112,dangling_wire_113}));
    defparam \pid_alt.un2_error_mulonly_0_21_0 .A_REG=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_21_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_21_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pid_alt.un2_error_mulonly_0_21_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_21_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pid_alt.un2_error_mulonly_0_21_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pid_alt.un2_error_mulonly_0_21_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_21_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_21_0 .NEG_TRIGGER=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_21_0 .MODE_8x8=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_21_0 .D_REG=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_21_0 .C_REG=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_21_0 .B_SIGNED=1'b1;
    defparam \pid_alt.un2_error_mulonly_0_21_0 .B_REG=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_21_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_21_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pid_alt.un2_error_mulonly_0_21_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_21_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pid_alt.un2_error_mulonly_0_21_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pid_alt.un2_error_mulonly_0_21_0 .A_SIGNED=1'b1;
    SB_MAC16 \pid_alt.un2_error_mulonly_0_21_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__43053),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__43051),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_114,dangling_wire_115,dangling_wire_116,dangling_wire_117,dangling_wire_118,dangling_wire_119,dangling_wire_120,dangling_wire_121,dangling_wire_122,dangling_wire_123,dangling_wire_124,dangling_wire_125,dangling_wire_126,dangling_wire_127,dangling_wire_128,dangling_wire_129}),
            .ADDSUBBOT(),
            .A({N__22132,N__22189,N__22247,N__21562,N__21620,N__21664,N__21709,N__21763,N__21820,N__21890,N__21946,N__21322,N__21383,N__21430,N__21472,N__24451}),
            .C({dangling_wire_130,dangling_wire_131,dangling_wire_132,dangling_wire_133,dangling_wire_134,dangling_wire_135,dangling_wire_136,dangling_wire_137,dangling_wire_138,dangling_wire_139,dangling_wire_140,dangling_wire_141,dangling_wire_142,dangling_wire_143,dangling_wire_144,dangling_wire_145}),
            .B({dangling_wire_146,dangling_wire_147,dangling_wire_148,dangling_wire_149,dangling_wire_150,dangling_wire_151,dangling_wire_152,dangling_wire_153,dangling_wire_154,dangling_wire_155,dangling_wire_156,N__43055,N__43052,dangling_wire_157,dangling_wire_158,N__43054}),
            .OHOLDTOP(),
            .O({dangling_wire_159,dangling_wire_160,dangling_wire_161,dangling_wire_162,dangling_wire_163,dangling_wire_164,dangling_wire_165,dangling_wire_166,dangling_wire_167,dangling_wire_168,\pid_alt.O_1_21 ,\pid_alt.O_1_20 ,\pid_alt.O_1_19 ,\pid_alt.O_1_18 ,\pid_alt.O_1_17 ,\pid_alt.O_1_16 ,\pid_alt.O_1_15 ,\pid_alt.O_2_14 ,\pid_alt.O_2_13 ,\pid_alt.O_2_12 ,\pid_alt.O_2_11 ,\pid_alt.O_2_10 ,\pid_alt.O_2_9 ,\pid_alt.O_2_8 ,\pid_alt.O_2_7 ,\pid_alt.O_2_6 ,\pid_alt.O_2_5 ,dangling_wire_169,dangling_wire_170,dangling_wire_171,dangling_wire_172,dangling_wire_173}));
    defparam \pid_alt.un1_error_d_reg_1_mulonly_0_24_0 .A_REG=1'b0;
    defparam \pid_alt.un1_error_d_reg_1_mulonly_0_24_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pid_alt.un1_error_d_reg_1_mulonly_0_24_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pid_alt.un1_error_d_reg_1_mulonly_0_24_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pid_alt.un1_error_d_reg_1_mulonly_0_24_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pid_alt.un1_error_d_reg_1_mulonly_0_24_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pid_alt.un1_error_d_reg_1_mulonly_0_24_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pid_alt.un1_error_d_reg_1_mulonly_0_24_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pid_alt.un1_error_d_reg_1_mulonly_0_24_0 .NEG_TRIGGER=1'b0;
    defparam \pid_alt.un1_error_d_reg_1_mulonly_0_24_0 .MODE_8x8=1'b0;
    defparam \pid_alt.un1_error_d_reg_1_mulonly_0_24_0 .D_REG=1'b0;
    defparam \pid_alt.un1_error_d_reg_1_mulonly_0_24_0 .C_REG=1'b0;
    defparam \pid_alt.un1_error_d_reg_1_mulonly_0_24_0 .B_SIGNED=1'b1;
    defparam \pid_alt.un1_error_d_reg_1_mulonly_0_24_0 .B_REG=1'b0;
    defparam \pid_alt.un1_error_d_reg_1_mulonly_0_24_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pid_alt.un1_error_d_reg_1_mulonly_0_24_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pid_alt.un1_error_d_reg_1_mulonly_0_24_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pid_alt.un1_error_d_reg_1_mulonly_0_24_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pid_alt.un1_error_d_reg_1_mulonly_0_24_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pid_alt.un1_error_d_reg_1_mulonly_0_24_0 .A_SIGNED=1'b1;
    SB_MAC16 \pid_alt.un1_error_d_reg_1_mulonly_0_24_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__43122),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__43110),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_174,dangling_wire_175,dangling_wire_176,dangling_wire_177,dangling_wire_178,dangling_wire_179,dangling_wire_180,dangling_wire_181,dangling_wire_182,dangling_wire_183,dangling_wire_184,dangling_wire_185,dangling_wire_186,dangling_wire_187,dangling_wire_188,dangling_wire_189}),
            .ADDSUBBOT(),
            .A({dangling_wire_190,N__46277,N__46019,N__46055,N__46094,N__46136,N__46343,N__45557,N__46388,N__46421,N__45860,N__45893,N__46310,N__46172,N__45452,N__17883}),
            .C({dangling_wire_191,dangling_wire_192,dangling_wire_193,dangling_wire_194,dangling_wire_195,dangling_wire_196,dangling_wire_197,dangling_wire_198,dangling_wire_199,dangling_wire_200,dangling_wire_201,dangling_wire_202,dangling_wire_203,dangling_wire_204,dangling_wire_205,dangling_wire_206}),
            .B({dangling_wire_207,dangling_wire_208,dangling_wire_209,dangling_wire_210,dangling_wire_211,dangling_wire_212,dangling_wire_213,dangling_wire_214,N__18392,N__18752,N__18731,N__18992,N__18416,N__18440,N__18368,N__18341}),
            .OHOLDTOP(),
            .O({dangling_wire_215,dangling_wire_216,dangling_wire_217,dangling_wire_218,dangling_wire_219,dangling_wire_220,dangling_wire_221,\pid_alt.un1_error_d_reg_1_24 ,\pid_alt.un1_error_d_reg_1_23 ,\pid_alt.un1_error_d_reg_1_22 ,\pid_alt.un1_error_d_reg_1_21 ,\pid_alt.un1_error_d_reg_1_20 ,\pid_alt.un1_error_d_reg_1_19 ,\pid_alt.un1_error_d_reg_1_18 ,\pid_alt.un1_error_d_reg_1_17 ,\pid_alt.un1_error_d_reg_1_16 ,\pid_alt.un1_error_d_reg_1_15 ,\pid_alt.O_14 ,\pid_alt.O_13 ,\pid_alt.O_12 ,\pid_alt.O_11 ,\pid_alt.O_10 ,\pid_alt.O_9 ,\pid_alt.O_8 ,\pid_alt.O_7 ,\pid_alt.O_6 ,\pid_alt.O_5 ,\pid_alt.O_4 ,dangling_wire_222,dangling_wire_223,dangling_wire_224,dangling_wire_225}));
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .A_REG=1'b0;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .NEG_TRIGGER=1'b0;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .MODE_8x8=1'b0;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .D_REG=1'b0;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .C_REG=1'b0;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .B_SIGNED=1'b1;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .B_REG=1'b0;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .A_SIGNED=1'b1;
    SB_MAC16 \pid_alt.un2_error_2_mulonly_0_24_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__43131),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__43138),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_226,dangling_wire_227,dangling_wire_228,dangling_wire_229,dangling_wire_230,dangling_wire_231,dangling_wire_232,dangling_wire_233,dangling_wire_234,dangling_wire_235,dangling_wire_236,dangling_wire_237,dangling_wire_238,dangling_wire_239,dangling_wire_240,dangling_wire_241}),
            .ADDSUBBOT(),
            .A({N__22149,N__22206,N__22248,N__21579,N__21627,N__21668,N__21726,N__21780,N__21837,N__21891,N__21963,N__21339,N__21390,N__21434,N__21486,N__24462}),
            .C({dangling_wire_242,dangling_wire_243,dangling_wire_244,dangling_wire_245,dangling_wire_246,dangling_wire_247,dangling_wire_248,dangling_wire_249,dangling_wire_250,dangling_wire_251,dangling_wire_252,dangling_wire_253,dangling_wire_254,dangling_wire_255,dangling_wire_256,dangling_wire_257}),
            .B({dangling_wire_258,dangling_wire_259,dangling_wire_260,dangling_wire_261,dangling_wire_262,dangling_wire_263,dangling_wire_264,dangling_wire_265,N__44877,N__33300,N__44154,N__45237,N__43230,N__36750,N__45078,N__23391}),
            .OHOLDTOP(),
            .O({dangling_wire_266,dangling_wire_267,dangling_wire_268,dangling_wire_269,dangling_wire_270,dangling_wire_271,dangling_wire_272,\pid_alt.O_24 ,\pid_alt.O_23 ,\pid_alt.O_22 ,\pid_alt.O_21 ,\pid_alt.O_20 ,\pid_alt.O_19 ,\pid_alt.O_18 ,\pid_alt.O_17 ,\pid_alt.O_16 ,\pid_alt.O_15 ,\pid_alt.O_0_14 ,\pid_alt.O_0_13 ,\pid_alt.O_0_12 ,\pid_alt.O_0_11 ,\pid_alt.O_0_10 ,\pid_alt.O_0_9 ,\pid_alt.O_0_8 ,\pid_alt.O_0_7 ,\pid_alt.O_0_6 ,\pid_alt.O_0_5 ,\pid_alt.O_0_4 ,dangling_wire_273,dangling_wire_274,dangling_wire_275,dangling_wire_276}));
    defparam \pid_alt.un1_error_d_reg_2_mulonly_0_16_0 .A_REG=1'b0;
    defparam \pid_alt.un1_error_d_reg_2_mulonly_0_16_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pid_alt.un1_error_d_reg_2_mulonly_0_16_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pid_alt.un1_error_d_reg_2_mulonly_0_16_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pid_alt.un1_error_d_reg_2_mulonly_0_16_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pid_alt.un1_error_d_reg_2_mulonly_0_16_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pid_alt.un1_error_d_reg_2_mulonly_0_16_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pid_alt.un1_error_d_reg_2_mulonly_0_16_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pid_alt.un1_error_d_reg_2_mulonly_0_16_0 .NEG_TRIGGER=1'b0;
    defparam \pid_alt.un1_error_d_reg_2_mulonly_0_16_0 .MODE_8x8=1'b0;
    defparam \pid_alt.un1_error_d_reg_2_mulonly_0_16_0 .D_REG=1'b0;
    defparam \pid_alt.un1_error_d_reg_2_mulonly_0_16_0 .C_REG=1'b0;
    defparam \pid_alt.un1_error_d_reg_2_mulonly_0_16_0 .B_SIGNED=1'b1;
    defparam \pid_alt.un1_error_d_reg_2_mulonly_0_16_0 .B_REG=1'b0;
    defparam \pid_alt.un1_error_d_reg_2_mulonly_0_16_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pid_alt.un1_error_d_reg_2_mulonly_0_16_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pid_alt.un1_error_d_reg_2_mulonly_0_16_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pid_alt.un1_error_d_reg_2_mulonly_0_16_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pid_alt.un1_error_d_reg_2_mulonly_0_16_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pid_alt.un1_error_d_reg_2_mulonly_0_16_0 .A_SIGNED=1'b1;
    SB_MAC16 \pid_alt.un1_error_d_reg_2_mulonly_0_16_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__43140),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__43139),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_277,dangling_wire_278,dangling_wire_279,dangling_wire_280,dangling_wire_281,dangling_wire_282,dangling_wire_283,dangling_wire_284,dangling_wire_285,dangling_wire_286,dangling_wire_287,dangling_wire_288,dangling_wire_289,dangling_wire_290,dangling_wire_291,dangling_wire_292}),
            .ADDSUBBOT(),
            .A({N__45692,N__45698,N__45694,N__45695,N__45693,N__45696,N__45691,N__45697,N__45690,N__44330,N__45596,N__45050,N__45734,N__45785,N__45935,N__45983}),
            .C({dangling_wire_293,dangling_wire_294,dangling_wire_295,dangling_wire_296,dangling_wire_297,dangling_wire_298,dangling_wire_299,dangling_wire_300,dangling_wire_301,dangling_wire_302,dangling_wire_303,dangling_wire_304,dangling_wire_305,dangling_wire_306,dangling_wire_307,dangling_wire_308}),
            .B({dangling_wire_309,dangling_wire_310,dangling_wire_311,dangling_wire_312,dangling_wire_313,dangling_wire_314,dangling_wire_315,dangling_wire_316,N__18393,N__18753,N__18732,N__18996,N__18417,N__18441,N__18369,N__18345}),
            .OHOLDTOP(),
            .O({dangling_wire_317,dangling_wire_318,dangling_wire_319,dangling_wire_320,dangling_wire_321,dangling_wire_322,dangling_wire_323,dangling_wire_324,dangling_wire_325,dangling_wire_326,dangling_wire_327,dangling_wire_328,dangling_wire_329,dangling_wire_330,dangling_wire_331,\pid_alt.un1_error_d_reg_2_16 ,\pid_alt.un1_error_d_reg_2_15 ,\pid_alt.un1_error_d_reg_2_14 ,\pid_alt.un1_error_d_reg_2_13 ,\pid_alt.un1_error_d_reg_2_12 ,\pid_alt.un1_error_d_reg_2_11 ,\pid_alt.un1_error_d_reg_2_10 ,\pid_alt.un1_error_d_reg_2_9 ,\pid_alt.un1_error_d_reg_2_8 ,\pid_alt.un1_error_d_reg_2_7 ,\pid_alt.un1_error_d_reg_2_6 ,\pid_alt.un1_error_d_reg_2_5 ,\pid_alt.un1_error_d_reg_2_4 ,\pid_alt.un1_error_d_reg_2_3 ,\pid_alt.un1_error_d_reg_2_2 ,\pid_alt.un1_error_d_reg_2_1 ,\pid_alt.un1_error_d_reg_2_0 }));
    defparam \pid_alt.un9_error_filt_2_mulonly_0_11_0 .A_REG=1'b0;
    defparam \pid_alt.un9_error_filt_2_mulonly_0_11_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pid_alt.un9_error_filt_2_mulonly_0_11_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pid_alt.un9_error_filt_2_mulonly_0_11_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pid_alt.un9_error_filt_2_mulonly_0_11_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pid_alt.un9_error_filt_2_mulonly_0_11_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pid_alt.un9_error_filt_2_mulonly_0_11_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pid_alt.un9_error_filt_2_mulonly_0_11_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pid_alt.un9_error_filt_2_mulonly_0_11_0 .NEG_TRIGGER=1'b0;
    defparam \pid_alt.un9_error_filt_2_mulonly_0_11_0 .MODE_8x8=1'b0;
    defparam \pid_alt.un9_error_filt_2_mulonly_0_11_0 .D_REG=1'b0;
    defparam \pid_alt.un9_error_filt_2_mulonly_0_11_0 .C_REG=1'b0;
    defparam \pid_alt.un9_error_filt_2_mulonly_0_11_0 .B_SIGNED=1'b1;
    defparam \pid_alt.un9_error_filt_2_mulonly_0_11_0 .B_REG=1'b0;
    defparam \pid_alt.un9_error_filt_2_mulonly_0_11_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pid_alt.un9_error_filt_2_mulonly_0_11_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pid_alt.un9_error_filt_2_mulonly_0_11_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pid_alt.un9_error_filt_2_mulonly_0_11_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pid_alt.un9_error_filt_2_mulonly_0_11_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pid_alt.un9_error_filt_2_mulonly_0_11_0 .A_SIGNED=1'b1;
    SB_MAC16 \pid_alt.un9_error_filt_2_mulonly_0_11_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__43128),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__43124),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_332,dangling_wire_333,dangling_wire_334,dangling_wire_335,dangling_wire_336,dangling_wire_337,dangling_wire_338,dangling_wire_339,dangling_wire_340,dangling_wire_341,dangling_wire_342,dangling_wire_343,dangling_wire_344,dangling_wire_345,dangling_wire_346,dangling_wire_347}),
            .ADDSUBBOT(),
            .A({N__45632,N__45635,N__45631,N__45636,N__45630,N__45633,N__45629,N__45634,N__45628,N__44307,N__45567,N__45027,N__45711,N__45762,N__45906,N__45954}),
            .C({dangling_wire_348,dangling_wire_349,dangling_wire_350,dangling_wire_351,dangling_wire_352,dangling_wire_353,dangling_wire_354,dangling_wire_355,dangling_wire_356,dangling_wire_357,dangling_wire_358,dangling_wire_359,dangling_wire_360,dangling_wire_361,dangling_wire_362,dangling_wire_363}),
            .B({dangling_wire_364,dangling_wire_365,dangling_wire_366,dangling_wire_367,dangling_wire_368,dangling_wire_369,dangling_wire_370,dangling_wire_371,dangling_wire_372,dangling_wire_373,dangling_wire_374,dangling_wire_375,dangling_wire_376,N__43127,N__43125,N__43126}),
            .OHOLDTOP(),
            .O({dangling_wire_377,dangling_wire_378,dangling_wire_379,dangling_wire_380,dangling_wire_381,dangling_wire_382,dangling_wire_383,dangling_wire_384,dangling_wire_385,dangling_wire_386,dangling_wire_387,dangling_wire_388,dangling_wire_389,dangling_wire_390,dangling_wire_391,dangling_wire_392,dangling_wire_393,dangling_wire_394,dangling_wire_395,dangling_wire_396,\pid_alt.un9_error_filt_2_11 ,\pid_alt.un9_error_filt_2_10 ,\pid_alt.un9_error_filt_2_9 ,\pid_alt.un9_error_filt_2_8 ,\pid_alt.un9_error_filt_2_7 ,\pid_alt.un9_error_filt_2_6 ,\pid_alt.un9_error_filt_2_5 ,\pid_alt.un9_error_filt_2_4 ,\pid_alt.un9_error_filt_2_3 ,\pid_alt.un9_error_filt_2_2 ,\pid_alt.un9_error_filt_2_1 ,\pid_alt.un9_error_filt_2_0 }));
    PRE_IO_GBUF clk_system_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__47734),
            .GLOBALBUFFEROUTPUT(clk_system_c_g));
    defparam clk_system_ibuf_gb_io_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD clk_system_ibuf_gb_io_iopad (
            .OE(N__47736),
            .DIN(N__47735),
            .DOUT(N__47734),
            .PACKAGEPIN(clk_system));
    defparam clk_system_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam clk_system_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO clk_system_ibuf_gb_io_preio (
            .PADOEN(N__47736),
            .PADOUT(N__47735),
            .PADIN(N__47734),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam uart_input_drone_ibuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD uart_input_drone_ibuf_iopad (
            .OE(N__47725),
            .DIN(N__47724),
            .DOUT(N__47723),
            .PACKAGEPIN(uart_input_drone));
    defparam uart_input_drone_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam uart_input_drone_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO uart_input_drone_ibuf_preio (
            .PADOEN(N__47725),
            .PADOUT(N__47724),
            .PADIN(N__47723),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(uart_input_drone_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam uart_input_pc_ibuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD uart_input_pc_ibuf_iopad (
            .OE(N__47716),
            .DIN(N__47715),
            .DOUT(N__47714),
            .PACKAGEPIN(uart_input_pc));
    defparam uart_input_pc_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam uart_input_pc_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO uart_input_pc_ibuf_preio (
            .PADOEN(N__47716),
            .PADOUT(N__47715),
            .PADIN(N__47714),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(uart_input_pc_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam debug_CH2_18A_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD debug_CH2_18A_obuf_iopad (
            .OE(N__47707),
            .DIN(N__47706),
            .DOUT(N__47705),
            .PACKAGEPIN(debug_CH2_18A));
    defparam debug_CH2_18A_obuf_preio.NEG_TRIGGER=1'b0;
    defparam debug_CH2_18A_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_CH2_18A_obuf_preio (
            .PADOEN(N__47707),
            .PADOUT(N__47706),
            .PADIN(N__47705),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__31229),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam debug_CH0_16A_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD debug_CH0_16A_obuf_iopad (
            .OE(N__47698),
            .DIN(N__47697),
            .DOUT(N__47696),
            .PACKAGEPIN(debug_CH0_16A));
    defparam debug_CH0_16A_obuf_preio.NEG_TRIGGER=1'b0;
    defparam debug_CH0_16A_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_CH0_16A_obuf_preio (
            .PADOEN(N__47698),
            .PADOUT(N__47697),
            .PADIN(N__47696),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__31404),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam debug_CH1_0A_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD debug_CH1_0A_obuf_iopad (
            .OE(N__47689),
            .DIN(N__47688),
            .DOUT(N__47687),
            .PACKAGEPIN(debug_CH1_0A));
    defparam debug_CH1_0A_obuf_preio.NEG_TRIGGER=1'b0;
    defparam debug_CH1_0A_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_CH1_0A_obuf_preio (
            .PADOEN(N__47689),
            .PADOUT(N__47688),
            .PADIN(N__47687),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__29600),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam debug_CH5_31B_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD debug_CH5_31B_obuf_iopad (
            .OE(N__47680),
            .DIN(N__47679),
            .DOUT(N__47678),
            .PACKAGEPIN(debug_CH5_31B));
    defparam debug_CH5_31B_obuf_preio.NEG_TRIGGER=1'b0;
    defparam debug_CH5_31B_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_CH5_31B_obuf_preio (
            .PADOEN(N__47680),
            .PADOUT(N__47679),
            .PADIN(N__47678),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam debug_CH4_2A_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD debug_CH4_2A_obuf_iopad (
            .OE(N__47671),
            .DIN(N__47670),
            .DOUT(N__47669),
            .PACKAGEPIN(debug_CH4_2A));
    defparam debug_CH4_2A_obuf_preio.NEG_TRIGGER=1'b0;
    defparam debug_CH4_2A_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_CH4_2A_obuf_preio (
            .PADOEN(N__47671),
            .PADOUT(N__47670),
            .PADIN(N__47669),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ppm_output_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD ppm_output_obuf_iopad (
            .OE(N__47662),
            .DIN(N__47661),
            .DOUT(N__47660),
            .PACKAGEPIN(ppm_output));
    defparam ppm_output_obuf_preio.NEG_TRIGGER=1'b0;
    defparam ppm_output_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO ppm_output_obuf_preio (
            .PADOEN(N__47662),
            .PADOUT(N__47661),
            .PADIN(N__47660),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__29457),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam debug_CH3_20A_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD debug_CH3_20A_obuf_iopad (
            .OE(N__47653),
            .DIN(N__47652),
            .DOUT(N__47651),
            .PACKAGEPIN(debug_CH3_20A));
    defparam debug_CH3_20A_obuf_preio.NEG_TRIGGER=1'b0;
    defparam debug_CH3_20A_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_CH3_20A_obuf_preio (
            .PADOEN(N__47653),
            .PADOUT(N__47652),
            .PADIN(N__47651),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__30578),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam debug_CH6_5B_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD debug_CH6_5B_obuf_iopad (
            .OE(N__47644),
            .DIN(N__47643),
            .DOUT(N__47642),
            .PACKAGEPIN(debug_CH6_5B));
    defparam debug_CH6_5B_obuf_preio.NEG_TRIGGER=1'b0;
    defparam debug_CH6_5B_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_CH6_5B_obuf_preio (
            .PADOEN(N__47644),
            .PADOUT(N__47643),
            .PADIN(N__47642),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__11503 (
            .O(N__47625),
            .I(N__47622));
    LocalMux I__11502 (
            .O(N__47622),
            .I(N__47619));
    Odrv4 I__11501 (
            .O(N__47619),
            .I(\pid_alt.O_0_13 ));
    InMux I__11500 (
            .O(N__47616),
            .I(N__47613));
    LocalMux I__11499 (
            .O(N__47613),
            .I(N__47610));
    Span12Mux_h I__11498 (
            .O(N__47610),
            .I(N__47607));
    Odrv12 I__11497 (
            .O(N__47607),
            .I(\pid_alt.error_i_regZ0Z_9 ));
    InMux I__11496 (
            .O(N__47604),
            .I(N__47601));
    LocalMux I__11495 (
            .O(N__47601),
            .I(N__47598));
    Odrv4 I__11494 (
            .O(N__47598),
            .I(\pid_alt.O_18 ));
    InMux I__11493 (
            .O(N__47595),
            .I(N__47592));
    LocalMux I__11492 (
            .O(N__47592),
            .I(N__47589));
    Odrv12 I__11491 (
            .O(N__47589),
            .I(\pid_alt.error_i_regZ0Z_14 ));
    InMux I__11490 (
            .O(N__47586),
            .I(N__47583));
    LocalMux I__11489 (
            .O(N__47583),
            .I(N__47580));
    Odrv4 I__11488 (
            .O(N__47580),
            .I(\pid_alt.O_24 ));
    InMux I__11487 (
            .O(N__47577),
            .I(N__47571));
    InMux I__11486 (
            .O(N__47576),
            .I(N__47571));
    LocalMux I__11485 (
            .O(N__47571),
            .I(N__47568));
    Span12Mux_h I__11484 (
            .O(N__47568),
            .I(N__47565));
    Odrv12 I__11483 (
            .O(N__47565),
            .I(\pid_alt.error_i_regZ0Z_20 ));
    InMux I__11482 (
            .O(N__47562),
            .I(N__47559));
    LocalMux I__11481 (
            .O(N__47559),
            .I(N__47556));
    Odrv4 I__11480 (
            .O(N__47556),
            .I(\pid_alt.O_21 ));
    InMux I__11479 (
            .O(N__47553),
            .I(N__47550));
    LocalMux I__11478 (
            .O(N__47550),
            .I(N__47547));
    Span12Mux_h I__11477 (
            .O(N__47547),
            .I(N__47544));
    Odrv12 I__11476 (
            .O(N__47544),
            .I(\pid_alt.error_i_regZ0Z_17 ));
    InMux I__11475 (
            .O(N__47541),
            .I(N__47538));
    LocalMux I__11474 (
            .O(N__47538),
            .I(N__47535));
    Odrv4 I__11473 (
            .O(N__47535),
            .I(\pid_alt.O_22 ));
    InMux I__11472 (
            .O(N__47532),
            .I(N__47529));
    LocalMux I__11471 (
            .O(N__47529),
            .I(N__47526));
    Span12Mux_h I__11470 (
            .O(N__47526),
            .I(N__47523));
    Odrv12 I__11469 (
            .O(N__47523),
            .I(\pid_alt.error_i_regZ0Z_18 ));
    InMux I__11468 (
            .O(N__47520),
            .I(N__47517));
    LocalMux I__11467 (
            .O(N__47517),
            .I(N__47514));
    Odrv4 I__11466 (
            .O(N__47514),
            .I(\pid_alt.O_20 ));
    InMux I__11465 (
            .O(N__47511),
            .I(N__47508));
    LocalMux I__11464 (
            .O(N__47508),
            .I(N__47505));
    Odrv12 I__11463 (
            .O(N__47505),
            .I(\pid_alt.error_i_regZ0Z_16 ));
    InMux I__11462 (
            .O(N__47502),
            .I(N__47499));
    LocalMux I__11461 (
            .O(N__47499),
            .I(\pid_alt.O_23 ));
    InMux I__11460 (
            .O(N__47496),
            .I(N__47493));
    LocalMux I__11459 (
            .O(N__47493),
            .I(N__47490));
    Span4Mux_h I__11458 (
            .O(N__47490),
            .I(N__47487));
    Span4Mux_h I__11457 (
            .O(N__47487),
            .I(N__47484));
    Span4Mux_h I__11456 (
            .O(N__47484),
            .I(N__47481));
    Odrv4 I__11455 (
            .O(N__47481),
            .I(\pid_alt.error_i_regZ0Z_19 ));
    ClkMux I__11454 (
            .O(N__47478),
            .I(N__46830));
    ClkMux I__11453 (
            .O(N__47477),
            .I(N__46830));
    ClkMux I__11452 (
            .O(N__47476),
            .I(N__46830));
    ClkMux I__11451 (
            .O(N__47475),
            .I(N__46830));
    ClkMux I__11450 (
            .O(N__47474),
            .I(N__46830));
    ClkMux I__11449 (
            .O(N__47473),
            .I(N__46830));
    ClkMux I__11448 (
            .O(N__47472),
            .I(N__46830));
    ClkMux I__11447 (
            .O(N__47471),
            .I(N__46830));
    ClkMux I__11446 (
            .O(N__47470),
            .I(N__46830));
    ClkMux I__11445 (
            .O(N__47469),
            .I(N__46830));
    ClkMux I__11444 (
            .O(N__47468),
            .I(N__46830));
    ClkMux I__11443 (
            .O(N__47467),
            .I(N__46830));
    ClkMux I__11442 (
            .O(N__47466),
            .I(N__46830));
    ClkMux I__11441 (
            .O(N__47465),
            .I(N__46830));
    ClkMux I__11440 (
            .O(N__47464),
            .I(N__46830));
    ClkMux I__11439 (
            .O(N__47463),
            .I(N__46830));
    ClkMux I__11438 (
            .O(N__47462),
            .I(N__46830));
    ClkMux I__11437 (
            .O(N__47461),
            .I(N__46830));
    ClkMux I__11436 (
            .O(N__47460),
            .I(N__46830));
    ClkMux I__11435 (
            .O(N__47459),
            .I(N__46830));
    ClkMux I__11434 (
            .O(N__47458),
            .I(N__46830));
    ClkMux I__11433 (
            .O(N__47457),
            .I(N__46830));
    ClkMux I__11432 (
            .O(N__47456),
            .I(N__46830));
    ClkMux I__11431 (
            .O(N__47455),
            .I(N__46830));
    ClkMux I__11430 (
            .O(N__47454),
            .I(N__46830));
    ClkMux I__11429 (
            .O(N__47453),
            .I(N__46830));
    ClkMux I__11428 (
            .O(N__47452),
            .I(N__46830));
    ClkMux I__11427 (
            .O(N__47451),
            .I(N__46830));
    ClkMux I__11426 (
            .O(N__47450),
            .I(N__46830));
    ClkMux I__11425 (
            .O(N__47449),
            .I(N__46830));
    ClkMux I__11424 (
            .O(N__47448),
            .I(N__46830));
    ClkMux I__11423 (
            .O(N__47447),
            .I(N__46830));
    ClkMux I__11422 (
            .O(N__47446),
            .I(N__46830));
    ClkMux I__11421 (
            .O(N__47445),
            .I(N__46830));
    ClkMux I__11420 (
            .O(N__47444),
            .I(N__46830));
    ClkMux I__11419 (
            .O(N__47443),
            .I(N__46830));
    ClkMux I__11418 (
            .O(N__47442),
            .I(N__46830));
    ClkMux I__11417 (
            .O(N__47441),
            .I(N__46830));
    ClkMux I__11416 (
            .O(N__47440),
            .I(N__46830));
    ClkMux I__11415 (
            .O(N__47439),
            .I(N__46830));
    ClkMux I__11414 (
            .O(N__47438),
            .I(N__46830));
    ClkMux I__11413 (
            .O(N__47437),
            .I(N__46830));
    ClkMux I__11412 (
            .O(N__47436),
            .I(N__46830));
    ClkMux I__11411 (
            .O(N__47435),
            .I(N__46830));
    ClkMux I__11410 (
            .O(N__47434),
            .I(N__46830));
    ClkMux I__11409 (
            .O(N__47433),
            .I(N__46830));
    ClkMux I__11408 (
            .O(N__47432),
            .I(N__46830));
    ClkMux I__11407 (
            .O(N__47431),
            .I(N__46830));
    ClkMux I__11406 (
            .O(N__47430),
            .I(N__46830));
    ClkMux I__11405 (
            .O(N__47429),
            .I(N__46830));
    ClkMux I__11404 (
            .O(N__47428),
            .I(N__46830));
    ClkMux I__11403 (
            .O(N__47427),
            .I(N__46830));
    ClkMux I__11402 (
            .O(N__47426),
            .I(N__46830));
    ClkMux I__11401 (
            .O(N__47425),
            .I(N__46830));
    ClkMux I__11400 (
            .O(N__47424),
            .I(N__46830));
    ClkMux I__11399 (
            .O(N__47423),
            .I(N__46830));
    ClkMux I__11398 (
            .O(N__47422),
            .I(N__46830));
    ClkMux I__11397 (
            .O(N__47421),
            .I(N__46830));
    ClkMux I__11396 (
            .O(N__47420),
            .I(N__46830));
    ClkMux I__11395 (
            .O(N__47419),
            .I(N__46830));
    ClkMux I__11394 (
            .O(N__47418),
            .I(N__46830));
    ClkMux I__11393 (
            .O(N__47417),
            .I(N__46830));
    ClkMux I__11392 (
            .O(N__47416),
            .I(N__46830));
    ClkMux I__11391 (
            .O(N__47415),
            .I(N__46830));
    ClkMux I__11390 (
            .O(N__47414),
            .I(N__46830));
    ClkMux I__11389 (
            .O(N__47413),
            .I(N__46830));
    ClkMux I__11388 (
            .O(N__47412),
            .I(N__46830));
    ClkMux I__11387 (
            .O(N__47411),
            .I(N__46830));
    ClkMux I__11386 (
            .O(N__47410),
            .I(N__46830));
    ClkMux I__11385 (
            .O(N__47409),
            .I(N__46830));
    ClkMux I__11384 (
            .O(N__47408),
            .I(N__46830));
    ClkMux I__11383 (
            .O(N__47407),
            .I(N__46830));
    ClkMux I__11382 (
            .O(N__47406),
            .I(N__46830));
    ClkMux I__11381 (
            .O(N__47405),
            .I(N__46830));
    ClkMux I__11380 (
            .O(N__47404),
            .I(N__46830));
    ClkMux I__11379 (
            .O(N__47403),
            .I(N__46830));
    ClkMux I__11378 (
            .O(N__47402),
            .I(N__46830));
    ClkMux I__11377 (
            .O(N__47401),
            .I(N__46830));
    ClkMux I__11376 (
            .O(N__47400),
            .I(N__46830));
    ClkMux I__11375 (
            .O(N__47399),
            .I(N__46830));
    ClkMux I__11374 (
            .O(N__47398),
            .I(N__46830));
    ClkMux I__11373 (
            .O(N__47397),
            .I(N__46830));
    ClkMux I__11372 (
            .O(N__47396),
            .I(N__46830));
    ClkMux I__11371 (
            .O(N__47395),
            .I(N__46830));
    ClkMux I__11370 (
            .O(N__47394),
            .I(N__46830));
    ClkMux I__11369 (
            .O(N__47393),
            .I(N__46830));
    ClkMux I__11368 (
            .O(N__47392),
            .I(N__46830));
    ClkMux I__11367 (
            .O(N__47391),
            .I(N__46830));
    ClkMux I__11366 (
            .O(N__47390),
            .I(N__46830));
    ClkMux I__11365 (
            .O(N__47389),
            .I(N__46830));
    ClkMux I__11364 (
            .O(N__47388),
            .I(N__46830));
    ClkMux I__11363 (
            .O(N__47387),
            .I(N__46830));
    ClkMux I__11362 (
            .O(N__47386),
            .I(N__46830));
    ClkMux I__11361 (
            .O(N__47385),
            .I(N__46830));
    ClkMux I__11360 (
            .O(N__47384),
            .I(N__46830));
    ClkMux I__11359 (
            .O(N__47383),
            .I(N__46830));
    ClkMux I__11358 (
            .O(N__47382),
            .I(N__46830));
    ClkMux I__11357 (
            .O(N__47381),
            .I(N__46830));
    ClkMux I__11356 (
            .O(N__47380),
            .I(N__46830));
    ClkMux I__11355 (
            .O(N__47379),
            .I(N__46830));
    ClkMux I__11354 (
            .O(N__47378),
            .I(N__46830));
    ClkMux I__11353 (
            .O(N__47377),
            .I(N__46830));
    ClkMux I__11352 (
            .O(N__47376),
            .I(N__46830));
    ClkMux I__11351 (
            .O(N__47375),
            .I(N__46830));
    ClkMux I__11350 (
            .O(N__47374),
            .I(N__46830));
    ClkMux I__11349 (
            .O(N__47373),
            .I(N__46830));
    ClkMux I__11348 (
            .O(N__47372),
            .I(N__46830));
    ClkMux I__11347 (
            .O(N__47371),
            .I(N__46830));
    ClkMux I__11346 (
            .O(N__47370),
            .I(N__46830));
    ClkMux I__11345 (
            .O(N__47369),
            .I(N__46830));
    ClkMux I__11344 (
            .O(N__47368),
            .I(N__46830));
    ClkMux I__11343 (
            .O(N__47367),
            .I(N__46830));
    ClkMux I__11342 (
            .O(N__47366),
            .I(N__46830));
    ClkMux I__11341 (
            .O(N__47365),
            .I(N__46830));
    ClkMux I__11340 (
            .O(N__47364),
            .I(N__46830));
    ClkMux I__11339 (
            .O(N__47363),
            .I(N__46830));
    ClkMux I__11338 (
            .O(N__47362),
            .I(N__46830));
    ClkMux I__11337 (
            .O(N__47361),
            .I(N__46830));
    ClkMux I__11336 (
            .O(N__47360),
            .I(N__46830));
    ClkMux I__11335 (
            .O(N__47359),
            .I(N__46830));
    ClkMux I__11334 (
            .O(N__47358),
            .I(N__46830));
    ClkMux I__11333 (
            .O(N__47357),
            .I(N__46830));
    ClkMux I__11332 (
            .O(N__47356),
            .I(N__46830));
    ClkMux I__11331 (
            .O(N__47355),
            .I(N__46830));
    ClkMux I__11330 (
            .O(N__47354),
            .I(N__46830));
    ClkMux I__11329 (
            .O(N__47353),
            .I(N__46830));
    ClkMux I__11328 (
            .O(N__47352),
            .I(N__46830));
    ClkMux I__11327 (
            .O(N__47351),
            .I(N__46830));
    ClkMux I__11326 (
            .O(N__47350),
            .I(N__46830));
    ClkMux I__11325 (
            .O(N__47349),
            .I(N__46830));
    ClkMux I__11324 (
            .O(N__47348),
            .I(N__46830));
    ClkMux I__11323 (
            .O(N__47347),
            .I(N__46830));
    ClkMux I__11322 (
            .O(N__47346),
            .I(N__46830));
    ClkMux I__11321 (
            .O(N__47345),
            .I(N__46830));
    ClkMux I__11320 (
            .O(N__47344),
            .I(N__46830));
    ClkMux I__11319 (
            .O(N__47343),
            .I(N__46830));
    ClkMux I__11318 (
            .O(N__47342),
            .I(N__46830));
    ClkMux I__11317 (
            .O(N__47341),
            .I(N__46830));
    ClkMux I__11316 (
            .O(N__47340),
            .I(N__46830));
    ClkMux I__11315 (
            .O(N__47339),
            .I(N__46830));
    ClkMux I__11314 (
            .O(N__47338),
            .I(N__46830));
    ClkMux I__11313 (
            .O(N__47337),
            .I(N__46830));
    ClkMux I__11312 (
            .O(N__47336),
            .I(N__46830));
    ClkMux I__11311 (
            .O(N__47335),
            .I(N__46830));
    ClkMux I__11310 (
            .O(N__47334),
            .I(N__46830));
    ClkMux I__11309 (
            .O(N__47333),
            .I(N__46830));
    ClkMux I__11308 (
            .O(N__47332),
            .I(N__46830));
    ClkMux I__11307 (
            .O(N__47331),
            .I(N__46830));
    ClkMux I__11306 (
            .O(N__47330),
            .I(N__46830));
    ClkMux I__11305 (
            .O(N__47329),
            .I(N__46830));
    ClkMux I__11304 (
            .O(N__47328),
            .I(N__46830));
    ClkMux I__11303 (
            .O(N__47327),
            .I(N__46830));
    ClkMux I__11302 (
            .O(N__47326),
            .I(N__46830));
    ClkMux I__11301 (
            .O(N__47325),
            .I(N__46830));
    ClkMux I__11300 (
            .O(N__47324),
            .I(N__46830));
    ClkMux I__11299 (
            .O(N__47323),
            .I(N__46830));
    ClkMux I__11298 (
            .O(N__47322),
            .I(N__46830));
    ClkMux I__11297 (
            .O(N__47321),
            .I(N__46830));
    ClkMux I__11296 (
            .O(N__47320),
            .I(N__46830));
    ClkMux I__11295 (
            .O(N__47319),
            .I(N__46830));
    ClkMux I__11294 (
            .O(N__47318),
            .I(N__46830));
    ClkMux I__11293 (
            .O(N__47317),
            .I(N__46830));
    ClkMux I__11292 (
            .O(N__47316),
            .I(N__46830));
    ClkMux I__11291 (
            .O(N__47315),
            .I(N__46830));
    ClkMux I__11290 (
            .O(N__47314),
            .I(N__46830));
    ClkMux I__11289 (
            .O(N__47313),
            .I(N__46830));
    ClkMux I__11288 (
            .O(N__47312),
            .I(N__46830));
    ClkMux I__11287 (
            .O(N__47311),
            .I(N__46830));
    ClkMux I__11286 (
            .O(N__47310),
            .I(N__46830));
    ClkMux I__11285 (
            .O(N__47309),
            .I(N__46830));
    ClkMux I__11284 (
            .O(N__47308),
            .I(N__46830));
    ClkMux I__11283 (
            .O(N__47307),
            .I(N__46830));
    ClkMux I__11282 (
            .O(N__47306),
            .I(N__46830));
    ClkMux I__11281 (
            .O(N__47305),
            .I(N__46830));
    ClkMux I__11280 (
            .O(N__47304),
            .I(N__46830));
    ClkMux I__11279 (
            .O(N__47303),
            .I(N__46830));
    ClkMux I__11278 (
            .O(N__47302),
            .I(N__46830));
    ClkMux I__11277 (
            .O(N__47301),
            .I(N__46830));
    ClkMux I__11276 (
            .O(N__47300),
            .I(N__46830));
    ClkMux I__11275 (
            .O(N__47299),
            .I(N__46830));
    ClkMux I__11274 (
            .O(N__47298),
            .I(N__46830));
    ClkMux I__11273 (
            .O(N__47297),
            .I(N__46830));
    ClkMux I__11272 (
            .O(N__47296),
            .I(N__46830));
    ClkMux I__11271 (
            .O(N__47295),
            .I(N__46830));
    ClkMux I__11270 (
            .O(N__47294),
            .I(N__46830));
    ClkMux I__11269 (
            .O(N__47293),
            .I(N__46830));
    ClkMux I__11268 (
            .O(N__47292),
            .I(N__46830));
    ClkMux I__11267 (
            .O(N__47291),
            .I(N__46830));
    ClkMux I__11266 (
            .O(N__47290),
            .I(N__46830));
    ClkMux I__11265 (
            .O(N__47289),
            .I(N__46830));
    ClkMux I__11264 (
            .O(N__47288),
            .I(N__46830));
    ClkMux I__11263 (
            .O(N__47287),
            .I(N__46830));
    ClkMux I__11262 (
            .O(N__47286),
            .I(N__46830));
    ClkMux I__11261 (
            .O(N__47285),
            .I(N__46830));
    ClkMux I__11260 (
            .O(N__47284),
            .I(N__46830));
    ClkMux I__11259 (
            .O(N__47283),
            .I(N__46830));
    ClkMux I__11258 (
            .O(N__47282),
            .I(N__46830));
    ClkMux I__11257 (
            .O(N__47281),
            .I(N__46830));
    ClkMux I__11256 (
            .O(N__47280),
            .I(N__46830));
    ClkMux I__11255 (
            .O(N__47279),
            .I(N__46830));
    ClkMux I__11254 (
            .O(N__47278),
            .I(N__46830));
    ClkMux I__11253 (
            .O(N__47277),
            .I(N__46830));
    ClkMux I__11252 (
            .O(N__47276),
            .I(N__46830));
    ClkMux I__11251 (
            .O(N__47275),
            .I(N__46830));
    ClkMux I__11250 (
            .O(N__47274),
            .I(N__46830));
    ClkMux I__11249 (
            .O(N__47273),
            .I(N__46830));
    ClkMux I__11248 (
            .O(N__47272),
            .I(N__46830));
    ClkMux I__11247 (
            .O(N__47271),
            .I(N__46830));
    ClkMux I__11246 (
            .O(N__47270),
            .I(N__46830));
    ClkMux I__11245 (
            .O(N__47269),
            .I(N__46830));
    ClkMux I__11244 (
            .O(N__47268),
            .I(N__46830));
    ClkMux I__11243 (
            .O(N__47267),
            .I(N__46830));
    ClkMux I__11242 (
            .O(N__47266),
            .I(N__46830));
    ClkMux I__11241 (
            .O(N__47265),
            .I(N__46830));
    ClkMux I__11240 (
            .O(N__47264),
            .I(N__46830));
    ClkMux I__11239 (
            .O(N__47263),
            .I(N__46830));
    GlobalMux I__11238 (
            .O(N__46830),
            .I(N__46827));
    gio2CtrlBuf I__11237 (
            .O(N__46827),
            .I(clk_system_c_g));
    CEMux I__11236 (
            .O(N__46824),
            .I(N__46695));
    CEMux I__11235 (
            .O(N__46823),
            .I(N__46695));
    CEMux I__11234 (
            .O(N__46822),
            .I(N__46695));
    CEMux I__11233 (
            .O(N__46821),
            .I(N__46695));
    CEMux I__11232 (
            .O(N__46820),
            .I(N__46695));
    CEMux I__11231 (
            .O(N__46819),
            .I(N__46695));
    CEMux I__11230 (
            .O(N__46818),
            .I(N__46695));
    CEMux I__11229 (
            .O(N__46817),
            .I(N__46695));
    CEMux I__11228 (
            .O(N__46816),
            .I(N__46695));
    CEMux I__11227 (
            .O(N__46815),
            .I(N__46695));
    CEMux I__11226 (
            .O(N__46814),
            .I(N__46695));
    CEMux I__11225 (
            .O(N__46813),
            .I(N__46695));
    CEMux I__11224 (
            .O(N__46812),
            .I(N__46695));
    CEMux I__11223 (
            .O(N__46811),
            .I(N__46695));
    CEMux I__11222 (
            .O(N__46810),
            .I(N__46695));
    CEMux I__11221 (
            .O(N__46809),
            .I(N__46695));
    CEMux I__11220 (
            .O(N__46808),
            .I(N__46695));
    CEMux I__11219 (
            .O(N__46807),
            .I(N__46695));
    CEMux I__11218 (
            .O(N__46806),
            .I(N__46695));
    CEMux I__11217 (
            .O(N__46805),
            .I(N__46695));
    CEMux I__11216 (
            .O(N__46804),
            .I(N__46695));
    CEMux I__11215 (
            .O(N__46803),
            .I(N__46695));
    CEMux I__11214 (
            .O(N__46802),
            .I(N__46695));
    CEMux I__11213 (
            .O(N__46801),
            .I(N__46695));
    CEMux I__11212 (
            .O(N__46800),
            .I(N__46695));
    CEMux I__11211 (
            .O(N__46799),
            .I(N__46695));
    CEMux I__11210 (
            .O(N__46798),
            .I(N__46695));
    CEMux I__11209 (
            .O(N__46797),
            .I(N__46695));
    CEMux I__11208 (
            .O(N__46796),
            .I(N__46695));
    CEMux I__11207 (
            .O(N__46795),
            .I(N__46695));
    CEMux I__11206 (
            .O(N__46794),
            .I(N__46695));
    CEMux I__11205 (
            .O(N__46793),
            .I(N__46695));
    CEMux I__11204 (
            .O(N__46792),
            .I(N__46695));
    CEMux I__11203 (
            .O(N__46791),
            .I(N__46695));
    CEMux I__11202 (
            .O(N__46790),
            .I(N__46695));
    CEMux I__11201 (
            .O(N__46789),
            .I(N__46695));
    CEMux I__11200 (
            .O(N__46788),
            .I(N__46695));
    CEMux I__11199 (
            .O(N__46787),
            .I(N__46695));
    CEMux I__11198 (
            .O(N__46786),
            .I(N__46695));
    CEMux I__11197 (
            .O(N__46785),
            .I(N__46695));
    CEMux I__11196 (
            .O(N__46784),
            .I(N__46695));
    CEMux I__11195 (
            .O(N__46783),
            .I(N__46695));
    CEMux I__11194 (
            .O(N__46782),
            .I(N__46695));
    GlobalMux I__11193 (
            .O(N__46695),
            .I(N__46692));
    gio2CtrlBuf I__11192 (
            .O(N__46692),
            .I(\pid_alt.N_410_0_g ));
    InMux I__11191 (
            .O(N__46689),
            .I(N__46671));
    InMux I__11190 (
            .O(N__46688),
            .I(N__46668));
    InMux I__11189 (
            .O(N__46687),
            .I(N__46663));
    InMux I__11188 (
            .O(N__46686),
            .I(N__46663));
    InMux I__11187 (
            .O(N__46685),
            .I(N__46658));
    InMux I__11186 (
            .O(N__46684),
            .I(N__46658));
    InMux I__11185 (
            .O(N__46683),
            .I(N__46655));
    InMux I__11184 (
            .O(N__46682),
            .I(N__46652));
    InMux I__11183 (
            .O(N__46681),
            .I(N__46649));
    InMux I__11182 (
            .O(N__46680),
            .I(N__46646));
    InMux I__11181 (
            .O(N__46679),
            .I(N__46643));
    InMux I__11180 (
            .O(N__46678),
            .I(N__46640));
    InMux I__11179 (
            .O(N__46677),
            .I(N__46635));
    InMux I__11178 (
            .O(N__46676),
            .I(N__46635));
    InMux I__11177 (
            .O(N__46675),
            .I(N__46632));
    InMux I__11176 (
            .O(N__46674),
            .I(N__46629));
    LocalMux I__11175 (
            .O(N__46671),
            .I(N__46582));
    LocalMux I__11174 (
            .O(N__46668),
            .I(N__46579));
    LocalMux I__11173 (
            .O(N__46663),
            .I(N__46576));
    LocalMux I__11172 (
            .O(N__46658),
            .I(N__46573));
    LocalMux I__11171 (
            .O(N__46655),
            .I(N__46570));
    LocalMux I__11170 (
            .O(N__46652),
            .I(N__46567));
    LocalMux I__11169 (
            .O(N__46649),
            .I(N__46564));
    LocalMux I__11168 (
            .O(N__46646),
            .I(N__46561));
    LocalMux I__11167 (
            .O(N__46643),
            .I(N__46558));
    LocalMux I__11166 (
            .O(N__46640),
            .I(N__46555));
    LocalMux I__11165 (
            .O(N__46635),
            .I(N__46552));
    LocalMux I__11164 (
            .O(N__46632),
            .I(N__46549));
    LocalMux I__11163 (
            .O(N__46629),
            .I(N__46546));
    SRMux I__11162 (
            .O(N__46628),
            .I(N__46431));
    SRMux I__11161 (
            .O(N__46627),
            .I(N__46431));
    SRMux I__11160 (
            .O(N__46626),
            .I(N__46431));
    SRMux I__11159 (
            .O(N__46625),
            .I(N__46431));
    SRMux I__11158 (
            .O(N__46624),
            .I(N__46431));
    SRMux I__11157 (
            .O(N__46623),
            .I(N__46431));
    SRMux I__11156 (
            .O(N__46622),
            .I(N__46431));
    SRMux I__11155 (
            .O(N__46621),
            .I(N__46431));
    SRMux I__11154 (
            .O(N__46620),
            .I(N__46431));
    SRMux I__11153 (
            .O(N__46619),
            .I(N__46431));
    SRMux I__11152 (
            .O(N__46618),
            .I(N__46431));
    SRMux I__11151 (
            .O(N__46617),
            .I(N__46431));
    SRMux I__11150 (
            .O(N__46616),
            .I(N__46431));
    SRMux I__11149 (
            .O(N__46615),
            .I(N__46431));
    SRMux I__11148 (
            .O(N__46614),
            .I(N__46431));
    SRMux I__11147 (
            .O(N__46613),
            .I(N__46431));
    SRMux I__11146 (
            .O(N__46612),
            .I(N__46431));
    SRMux I__11145 (
            .O(N__46611),
            .I(N__46431));
    SRMux I__11144 (
            .O(N__46610),
            .I(N__46431));
    SRMux I__11143 (
            .O(N__46609),
            .I(N__46431));
    SRMux I__11142 (
            .O(N__46608),
            .I(N__46431));
    SRMux I__11141 (
            .O(N__46607),
            .I(N__46431));
    SRMux I__11140 (
            .O(N__46606),
            .I(N__46431));
    SRMux I__11139 (
            .O(N__46605),
            .I(N__46431));
    SRMux I__11138 (
            .O(N__46604),
            .I(N__46431));
    SRMux I__11137 (
            .O(N__46603),
            .I(N__46431));
    SRMux I__11136 (
            .O(N__46602),
            .I(N__46431));
    SRMux I__11135 (
            .O(N__46601),
            .I(N__46431));
    SRMux I__11134 (
            .O(N__46600),
            .I(N__46431));
    SRMux I__11133 (
            .O(N__46599),
            .I(N__46431));
    SRMux I__11132 (
            .O(N__46598),
            .I(N__46431));
    SRMux I__11131 (
            .O(N__46597),
            .I(N__46431));
    SRMux I__11130 (
            .O(N__46596),
            .I(N__46431));
    SRMux I__11129 (
            .O(N__46595),
            .I(N__46431));
    SRMux I__11128 (
            .O(N__46594),
            .I(N__46431));
    SRMux I__11127 (
            .O(N__46593),
            .I(N__46431));
    SRMux I__11126 (
            .O(N__46592),
            .I(N__46431));
    SRMux I__11125 (
            .O(N__46591),
            .I(N__46431));
    SRMux I__11124 (
            .O(N__46590),
            .I(N__46431));
    SRMux I__11123 (
            .O(N__46589),
            .I(N__46431));
    SRMux I__11122 (
            .O(N__46588),
            .I(N__46431));
    SRMux I__11121 (
            .O(N__46587),
            .I(N__46431));
    SRMux I__11120 (
            .O(N__46586),
            .I(N__46431));
    SRMux I__11119 (
            .O(N__46585),
            .I(N__46431));
    Glb2LocalMux I__11118 (
            .O(N__46582),
            .I(N__46431));
    Glb2LocalMux I__11117 (
            .O(N__46579),
            .I(N__46431));
    Glb2LocalMux I__11116 (
            .O(N__46576),
            .I(N__46431));
    Glb2LocalMux I__11115 (
            .O(N__46573),
            .I(N__46431));
    Glb2LocalMux I__11114 (
            .O(N__46570),
            .I(N__46431));
    Glb2LocalMux I__11113 (
            .O(N__46567),
            .I(N__46431));
    Glb2LocalMux I__11112 (
            .O(N__46564),
            .I(N__46431));
    Glb2LocalMux I__11111 (
            .O(N__46561),
            .I(N__46431));
    Glb2LocalMux I__11110 (
            .O(N__46558),
            .I(N__46431));
    Glb2LocalMux I__11109 (
            .O(N__46555),
            .I(N__46431));
    Glb2LocalMux I__11108 (
            .O(N__46552),
            .I(N__46431));
    Glb2LocalMux I__11107 (
            .O(N__46549),
            .I(N__46431));
    Glb2LocalMux I__11106 (
            .O(N__46546),
            .I(N__46431));
    GlobalMux I__11105 (
            .O(N__46431),
            .I(N__46428));
    gio2CtrlBuf I__11104 (
            .O(N__46428),
            .I(N_411_g));
    InMux I__11103 (
            .O(N__46425),
            .I(N__46422));
    LocalMux I__11102 (
            .O(N__46422),
            .I(N__46418));
    InMux I__11101 (
            .O(N__46421),
            .I(N__46415));
    Span12Mux_s2_h I__11100 (
            .O(N__46418),
            .I(N__46412));
    LocalMux I__11099 (
            .O(N__46415),
            .I(N__46409));
    Span12Mux_h I__11098 (
            .O(N__46412),
            .I(N__46406));
    Span4Mux_v I__11097 (
            .O(N__46409),
            .I(N__46403));
    Odrv12 I__11096 (
            .O(N__46406),
            .I(\pid_alt.error_filt_6 ));
    Odrv4 I__11095 (
            .O(N__46403),
            .I(\pid_alt.error_filt_6 ));
    InMux I__11094 (
            .O(N__46398),
            .I(N__46395));
    LocalMux I__11093 (
            .O(N__46395),
            .I(\pid_alt.error_filt_prevZ0Z_6 ));
    InMux I__11092 (
            .O(N__46392),
            .I(N__46389));
    LocalMux I__11091 (
            .O(N__46389),
            .I(N__46385));
    InMux I__11090 (
            .O(N__46388),
            .I(N__46382));
    Span12Mux_s3_h I__11089 (
            .O(N__46385),
            .I(N__46379));
    LocalMux I__11088 (
            .O(N__46382),
            .I(N__46376));
    Span12Mux_h I__11087 (
            .O(N__46379),
            .I(N__46373));
    Span4Mux_v I__11086 (
            .O(N__46376),
            .I(N__46370));
    Odrv12 I__11085 (
            .O(N__46373),
            .I(\pid_alt.error_filt_7 ));
    Odrv4 I__11084 (
            .O(N__46370),
            .I(\pid_alt.error_filt_7 ));
    InMux I__11083 (
            .O(N__46365),
            .I(N__46362));
    LocalMux I__11082 (
            .O(N__46362),
            .I(\pid_alt.error_filt_prevZ0Z_7 ));
    InMux I__11081 (
            .O(N__46359),
            .I(N__46356));
    LocalMux I__11080 (
            .O(N__46356),
            .I(N__46353));
    Span4Mux_v I__11079 (
            .O(N__46353),
            .I(N__46350));
    Span4Mux_h I__11078 (
            .O(N__46350),
            .I(N__46347));
    Span4Mux_h I__11077 (
            .O(N__46347),
            .I(N__46344));
    Span4Mux_h I__11076 (
            .O(N__46344),
            .I(N__46340));
    InMux I__11075 (
            .O(N__46343),
            .I(N__46337));
    Span4Mux_h I__11074 (
            .O(N__46340),
            .I(N__46334));
    LocalMux I__11073 (
            .O(N__46337),
            .I(N__46331));
    Span4Mux_h I__11072 (
            .O(N__46334),
            .I(N__46328));
    Span4Mux_v I__11071 (
            .O(N__46331),
            .I(N__46325));
    Odrv4 I__11070 (
            .O(N__46328),
            .I(\pid_alt.error_filt_9 ));
    Odrv4 I__11069 (
            .O(N__46325),
            .I(\pid_alt.error_filt_9 ));
    InMux I__11068 (
            .O(N__46320),
            .I(N__46317));
    LocalMux I__11067 (
            .O(N__46317),
            .I(\pid_alt.error_filt_prevZ0Z_9 ));
    InMux I__11066 (
            .O(N__46314),
            .I(N__46311));
    LocalMux I__11065 (
            .O(N__46311),
            .I(N__46307));
    InMux I__11064 (
            .O(N__46310),
            .I(N__46304));
    Span12Mux_s7_h I__11063 (
            .O(N__46307),
            .I(N__46301));
    LocalMux I__11062 (
            .O(N__46304),
            .I(N__46298));
    Span12Mux_h I__11061 (
            .O(N__46301),
            .I(N__46295));
    Span4Mux_s1_h I__11060 (
            .O(N__46298),
            .I(N__46292));
    Odrv12 I__11059 (
            .O(N__46295),
            .I(\pid_alt.error_filt_3 ));
    Odrv4 I__11058 (
            .O(N__46292),
            .I(\pid_alt.error_filt_3 ));
    InMux I__11057 (
            .O(N__46287),
            .I(N__46284));
    LocalMux I__11056 (
            .O(N__46284),
            .I(\pid_alt.error_filt_prevZ0Z_3 ));
    InMux I__11055 (
            .O(N__46281),
            .I(N__46278));
    LocalMux I__11054 (
            .O(N__46278),
            .I(N__46274));
    InMux I__11053 (
            .O(N__46277),
            .I(N__46271));
    Span12Mux_s2_h I__11052 (
            .O(N__46274),
            .I(N__46268));
    LocalMux I__11051 (
            .O(N__46271),
            .I(N__46265));
    Span12Mux_h I__11050 (
            .O(N__46268),
            .I(N__46262));
    Span4Mux_v I__11049 (
            .O(N__46265),
            .I(N__46259));
    Odrv12 I__11048 (
            .O(N__46262),
            .I(\pid_alt.error_filt_14 ));
    Odrv4 I__11047 (
            .O(N__46259),
            .I(\pid_alt.error_filt_14 ));
    InMux I__11046 (
            .O(N__46254),
            .I(N__46251));
    LocalMux I__11045 (
            .O(N__46251),
            .I(\pid_alt.error_filt_prevZ0Z_14 ));
    InMux I__11044 (
            .O(N__46248),
            .I(N__46245));
    LocalMux I__11043 (
            .O(N__46245),
            .I(N__46242));
    Odrv4 I__11042 (
            .O(N__46242),
            .I(\pid_alt.O_0_11 ));
    CascadeMux I__11041 (
            .O(N__46239),
            .I(N__46236));
    InMux I__11040 (
            .O(N__46236),
            .I(N__46233));
    LocalMux I__11039 (
            .O(N__46233),
            .I(N__46230));
    Span12Mux_h I__11038 (
            .O(N__46230),
            .I(N__46227));
    Odrv12 I__11037 (
            .O(N__46227),
            .I(\pid_alt.error_i_regZ0Z_7 ));
    InMux I__11036 (
            .O(N__46224),
            .I(N__46221));
    LocalMux I__11035 (
            .O(N__46221),
            .I(N__46218));
    Odrv4 I__11034 (
            .O(N__46218),
            .I(\pid_alt.O_0_10 ));
    InMux I__11033 (
            .O(N__46215),
            .I(N__46212));
    LocalMux I__11032 (
            .O(N__46212),
            .I(N__46209));
    Span12Mux_h I__11031 (
            .O(N__46209),
            .I(N__46206));
    Odrv12 I__11030 (
            .O(N__46206),
            .I(\pid_alt.error_i_regZ0Z_6 ));
    InMux I__11029 (
            .O(N__46203),
            .I(N__46200));
    LocalMux I__11028 (
            .O(N__46200),
            .I(N__46197));
    Odrv4 I__11027 (
            .O(N__46197),
            .I(\pid_alt.O_19 ));
    InMux I__11026 (
            .O(N__46194),
            .I(N__46191));
    LocalMux I__11025 (
            .O(N__46191),
            .I(N__46188));
    Span4Mux_h I__11024 (
            .O(N__46188),
            .I(N__46185));
    Span4Mux_h I__11023 (
            .O(N__46185),
            .I(N__46182));
    Span4Mux_h I__11022 (
            .O(N__46182),
            .I(N__46179));
    Odrv4 I__11021 (
            .O(N__46179),
            .I(\pid_alt.error_i_regZ0Z_15 ));
    InMux I__11020 (
            .O(N__46176),
            .I(N__46173));
    LocalMux I__11019 (
            .O(N__46173),
            .I(N__46169));
    InMux I__11018 (
            .O(N__46172),
            .I(N__46166));
    Span12Mux_h I__11017 (
            .O(N__46169),
            .I(N__46163));
    LocalMux I__11016 (
            .O(N__46166),
            .I(N__46160));
    Span12Mux_h I__11015 (
            .O(N__46163),
            .I(N__46157));
    Span4Mux_s1_h I__11014 (
            .O(N__46160),
            .I(N__46154));
    Odrv12 I__11013 (
            .O(N__46157),
            .I(\pid_alt.error_filt_2 ));
    Odrv4 I__11012 (
            .O(N__46154),
            .I(\pid_alt.error_filt_2 ));
    InMux I__11011 (
            .O(N__46149),
            .I(N__46146));
    LocalMux I__11010 (
            .O(N__46146),
            .I(N__46143));
    Odrv4 I__11009 (
            .O(N__46143),
            .I(\pid_alt.error_filt_prevZ0Z_2 ));
    InMux I__11008 (
            .O(N__46140),
            .I(N__46137));
    LocalMux I__11007 (
            .O(N__46137),
            .I(N__46133));
    InMux I__11006 (
            .O(N__46136),
            .I(N__46130));
    Span12Mux_h I__11005 (
            .O(N__46133),
            .I(N__46127));
    LocalMux I__11004 (
            .O(N__46130),
            .I(N__46124));
    Span12Mux_h I__11003 (
            .O(N__46127),
            .I(N__46121));
    Span4Mux_v I__11002 (
            .O(N__46124),
            .I(N__46118));
    Odrv12 I__11001 (
            .O(N__46121),
            .I(\pid_alt.error_filt_10 ));
    Odrv4 I__11000 (
            .O(N__46118),
            .I(\pid_alt.error_filt_10 ));
    InMux I__10999 (
            .O(N__46113),
            .I(N__46110));
    LocalMux I__10998 (
            .O(N__46110),
            .I(N__46107));
    Odrv4 I__10997 (
            .O(N__46107),
            .I(\pid_alt.error_filt_prevZ0Z_10 ));
    InMux I__10996 (
            .O(N__46104),
            .I(N__46101));
    LocalMux I__10995 (
            .O(N__46101),
            .I(N__46098));
    Span4Mux_v I__10994 (
            .O(N__46098),
            .I(N__46095));
    Span4Mux_h I__10993 (
            .O(N__46095),
            .I(N__46091));
    InMux I__10992 (
            .O(N__46094),
            .I(N__46088));
    Sp12to4 I__10991 (
            .O(N__46091),
            .I(N__46085));
    LocalMux I__10990 (
            .O(N__46088),
            .I(N__46082));
    Span12Mux_h I__10989 (
            .O(N__46085),
            .I(N__46079));
    Span4Mux_v I__10988 (
            .O(N__46082),
            .I(N__46076));
    Odrv12 I__10987 (
            .O(N__46079),
            .I(\pid_alt.error_filt_11 ));
    Odrv4 I__10986 (
            .O(N__46076),
            .I(\pid_alt.error_filt_11 ));
    InMux I__10985 (
            .O(N__46071),
            .I(N__46068));
    LocalMux I__10984 (
            .O(N__46068),
            .I(N__46065));
    Odrv4 I__10983 (
            .O(N__46065),
            .I(\pid_alt.error_filt_prevZ0Z_11 ));
    InMux I__10982 (
            .O(N__46062),
            .I(N__46059));
    LocalMux I__10981 (
            .O(N__46059),
            .I(N__46056));
    Span4Mux_v I__10980 (
            .O(N__46056),
            .I(N__46052));
    InMux I__10979 (
            .O(N__46055),
            .I(N__46049));
    Sp12to4 I__10978 (
            .O(N__46052),
            .I(N__46046));
    LocalMux I__10977 (
            .O(N__46049),
            .I(N__46043));
    Span12Mux_h I__10976 (
            .O(N__46046),
            .I(N__46040));
    Span4Mux_v I__10975 (
            .O(N__46043),
            .I(N__46037));
    Odrv12 I__10974 (
            .O(N__46040),
            .I(\pid_alt.error_filt_12 ));
    Odrv4 I__10973 (
            .O(N__46037),
            .I(\pid_alt.error_filt_12 ));
    InMux I__10972 (
            .O(N__46032),
            .I(N__46029));
    LocalMux I__10971 (
            .O(N__46029),
            .I(N__46026));
    Odrv4 I__10970 (
            .O(N__46026),
            .I(\pid_alt.error_filt_prevZ0Z_12 ));
    InMux I__10969 (
            .O(N__46023),
            .I(N__46020));
    LocalMux I__10968 (
            .O(N__46020),
            .I(N__46016));
    InMux I__10967 (
            .O(N__46019),
            .I(N__46013));
    Span12Mux_v I__10966 (
            .O(N__46016),
            .I(N__46010));
    LocalMux I__10965 (
            .O(N__46013),
            .I(N__46007));
    Span12Mux_h I__10964 (
            .O(N__46010),
            .I(N__46004));
    Span4Mux_v I__10963 (
            .O(N__46007),
            .I(N__46001));
    Odrv12 I__10962 (
            .O(N__46004),
            .I(\pid_alt.error_filt_13 ));
    Odrv4 I__10961 (
            .O(N__46001),
            .I(\pid_alt.error_filt_13 ));
    InMux I__10960 (
            .O(N__45996),
            .I(N__45993));
    LocalMux I__10959 (
            .O(N__45993),
            .I(N__45990));
    Odrv4 I__10958 (
            .O(N__45990),
            .I(\pid_alt.error_filt_prevZ0Z_13 ));
    InMux I__10957 (
            .O(N__45987),
            .I(N__45984));
    LocalMux I__10956 (
            .O(N__45984),
            .I(N__45980));
    InMux I__10955 (
            .O(N__45983),
            .I(N__45977));
    Span4Mux_v I__10954 (
            .O(N__45980),
            .I(N__45974));
    LocalMux I__10953 (
            .O(N__45977),
            .I(N__45971));
    Sp12to4 I__10952 (
            .O(N__45974),
            .I(N__45968));
    Span4Mux_v I__10951 (
            .O(N__45971),
            .I(N__45965));
    Span12Mux_h I__10950 (
            .O(N__45968),
            .I(N__45962));
    Span4Mux_v I__10949 (
            .O(N__45965),
            .I(N__45959));
    Odrv12 I__10948 (
            .O(N__45962),
            .I(\pid_alt.error_filt_15 ));
    Odrv4 I__10947 (
            .O(N__45959),
            .I(\pid_alt.error_filt_15 ));
    InMux I__10946 (
            .O(N__45954),
            .I(N__45951));
    LocalMux I__10945 (
            .O(N__45951),
            .I(N__45948));
    Span4Mux_s0_h I__10944 (
            .O(N__45948),
            .I(N__45945));
    Odrv4 I__10943 (
            .O(N__45945),
            .I(\pid_alt.error_filt_prevZ0Z_15 ));
    InMux I__10942 (
            .O(N__45942),
            .I(N__45939));
    LocalMux I__10941 (
            .O(N__45939),
            .I(N__45936));
    Span4Mux_v I__10940 (
            .O(N__45936),
            .I(N__45932));
    InMux I__10939 (
            .O(N__45935),
            .I(N__45929));
    Sp12to4 I__10938 (
            .O(N__45932),
            .I(N__45926));
    LocalMux I__10937 (
            .O(N__45929),
            .I(N__45923));
    Span12Mux_s4_h I__10936 (
            .O(N__45926),
            .I(N__45920));
    Span4Mux_v I__10935 (
            .O(N__45923),
            .I(N__45917));
    Span12Mux_h I__10934 (
            .O(N__45920),
            .I(N__45914));
    Span4Mux_v I__10933 (
            .O(N__45917),
            .I(N__45911));
    Odrv12 I__10932 (
            .O(N__45914),
            .I(\pid_alt.error_filt_16 ));
    Odrv4 I__10931 (
            .O(N__45911),
            .I(\pid_alt.error_filt_16 ));
    InMux I__10930 (
            .O(N__45906),
            .I(N__45903));
    LocalMux I__10929 (
            .O(N__45903),
            .I(N__45900));
    Span4Mux_s0_h I__10928 (
            .O(N__45900),
            .I(N__45897));
    Odrv4 I__10927 (
            .O(N__45897),
            .I(\pid_alt.error_filt_prevZ0Z_16 ));
    InMux I__10926 (
            .O(N__45894),
            .I(N__45890));
    InMux I__10925 (
            .O(N__45893),
            .I(N__45887));
    LocalMux I__10924 (
            .O(N__45890),
            .I(N__45884));
    LocalMux I__10923 (
            .O(N__45887),
            .I(N__45881));
    Span12Mux_h I__10922 (
            .O(N__45884),
            .I(N__45878));
    Span4Mux_s2_h I__10921 (
            .O(N__45881),
            .I(N__45875));
    Odrv12 I__10920 (
            .O(N__45878),
            .I(\pid_alt.error_filt_4 ));
    Odrv4 I__10919 (
            .O(N__45875),
            .I(\pid_alt.error_filt_4 ));
    InMux I__10918 (
            .O(N__45870),
            .I(N__45867));
    LocalMux I__10917 (
            .O(N__45867),
            .I(\pid_alt.error_filt_prevZ0Z_4 ));
    InMux I__10916 (
            .O(N__45864),
            .I(N__45861));
    LocalMux I__10915 (
            .O(N__45861),
            .I(N__45857));
    InMux I__10914 (
            .O(N__45860),
            .I(N__45854));
    Span12Mux_s1_h I__10913 (
            .O(N__45857),
            .I(N__45851));
    LocalMux I__10912 (
            .O(N__45854),
            .I(N__45848));
    Span12Mux_h I__10911 (
            .O(N__45851),
            .I(N__45845));
    Span4Mux_s1_h I__10910 (
            .O(N__45848),
            .I(N__45842));
    Odrv12 I__10909 (
            .O(N__45845),
            .I(\pid_alt.error_filt_5 ));
    Odrv4 I__10908 (
            .O(N__45842),
            .I(\pid_alt.error_filt_5 ));
    InMux I__10907 (
            .O(N__45837),
            .I(N__45834));
    LocalMux I__10906 (
            .O(N__45834),
            .I(\pid_alt.error_filt_prevZ0Z_5 ));
    InMux I__10905 (
            .O(N__45831),
            .I(N__45828));
    LocalMux I__10904 (
            .O(N__45828),
            .I(N__45825));
    Span4Mux_h I__10903 (
            .O(N__45825),
            .I(N__45822));
    Odrv4 I__10902 (
            .O(N__45822),
            .I(\pid_alt.O_17 ));
    CascadeMux I__10901 (
            .O(N__45819),
            .I(N__45816));
    InMux I__10900 (
            .O(N__45816),
            .I(N__45813));
    LocalMux I__10899 (
            .O(N__45813),
            .I(N__45810));
    Span4Mux_h I__10898 (
            .O(N__45810),
            .I(N__45807));
    Span4Mux_h I__10897 (
            .O(N__45807),
            .I(N__45804));
    Span4Mux_h I__10896 (
            .O(N__45804),
            .I(N__45801));
    Odrv4 I__10895 (
            .O(N__45801),
            .I(\pid_alt.error_i_regZ0Z_13 ));
    InMux I__10894 (
            .O(N__45798),
            .I(N__45795));
    LocalMux I__10893 (
            .O(N__45795),
            .I(N__45792));
    Span4Mux_s3_h I__10892 (
            .O(N__45792),
            .I(N__45789));
    Span4Mux_v I__10891 (
            .O(N__45789),
            .I(N__45786));
    Span4Mux_v I__10890 (
            .O(N__45786),
            .I(N__45782));
    InMux I__10889 (
            .O(N__45785),
            .I(N__45779));
    Sp12to4 I__10888 (
            .O(N__45782),
            .I(N__45776));
    LocalMux I__10887 (
            .O(N__45779),
            .I(N__45773));
    Span12Mux_h I__10886 (
            .O(N__45776),
            .I(N__45770));
    Span12Mux_s1_h I__10885 (
            .O(N__45773),
            .I(N__45767));
    Odrv12 I__10884 (
            .O(N__45770),
            .I(\pid_alt.error_filt_17 ));
    Odrv12 I__10883 (
            .O(N__45767),
            .I(\pid_alt.error_filt_17 ));
    InMux I__10882 (
            .O(N__45762),
            .I(N__45759));
    LocalMux I__10881 (
            .O(N__45759),
            .I(N__45756));
    Span4Mux_s1_h I__10880 (
            .O(N__45756),
            .I(N__45753));
    Odrv4 I__10879 (
            .O(N__45753),
            .I(\pid_alt.error_filt_prevZ0Z_17 ));
    InMux I__10878 (
            .O(N__45750),
            .I(N__45747));
    LocalMux I__10877 (
            .O(N__45747),
            .I(N__45744));
    Span4Mux_h I__10876 (
            .O(N__45744),
            .I(N__45741));
    Span4Mux_h I__10875 (
            .O(N__45741),
            .I(N__45738));
    Span4Mux_h I__10874 (
            .O(N__45738),
            .I(N__45735));
    Span4Mux_h I__10873 (
            .O(N__45735),
            .I(N__45731));
    InMux I__10872 (
            .O(N__45734),
            .I(N__45728));
    Span4Mux_h I__10871 (
            .O(N__45731),
            .I(N__45725));
    LocalMux I__10870 (
            .O(N__45728),
            .I(N__45722));
    Span4Mux_h I__10869 (
            .O(N__45725),
            .I(N__45717));
    Span4Mux_v I__10868 (
            .O(N__45722),
            .I(N__45717));
    Span4Mux_v I__10867 (
            .O(N__45717),
            .I(N__45714));
    Odrv4 I__10866 (
            .O(N__45714),
            .I(\pid_alt.error_filt_18 ));
    InMux I__10865 (
            .O(N__45711),
            .I(N__45708));
    LocalMux I__10864 (
            .O(N__45708),
            .I(N__45705));
    Odrv4 I__10863 (
            .O(N__45705),
            .I(\pid_alt.error_filt_prevZ0Z_18 ));
    InMux I__10862 (
            .O(N__45702),
            .I(N__45699));
    LocalMux I__10861 (
            .O(N__45699),
            .I(N__45687));
    InMux I__10860 (
            .O(N__45698),
            .I(N__45678));
    InMux I__10859 (
            .O(N__45697),
            .I(N__45678));
    InMux I__10858 (
            .O(N__45696),
            .I(N__45678));
    InMux I__10857 (
            .O(N__45695),
            .I(N__45678));
    InMux I__10856 (
            .O(N__45694),
            .I(N__45667));
    InMux I__10855 (
            .O(N__45693),
            .I(N__45667));
    InMux I__10854 (
            .O(N__45692),
            .I(N__45667));
    InMux I__10853 (
            .O(N__45691),
            .I(N__45667));
    InMux I__10852 (
            .O(N__45690),
            .I(N__45667));
    Span4Mux_s2_h I__10851 (
            .O(N__45687),
            .I(N__45664));
    LocalMux I__10850 (
            .O(N__45678),
            .I(N__45659));
    LocalMux I__10849 (
            .O(N__45667),
            .I(N__45659));
    Sp12to4 I__10848 (
            .O(N__45664),
            .I(N__45656));
    Span4Mux_s1_h I__10847 (
            .O(N__45659),
            .I(N__45653));
    Span12Mux_v I__10846 (
            .O(N__45656),
            .I(N__45650));
    Span4Mux_v I__10845 (
            .O(N__45653),
            .I(N__45647));
    Span12Mux_h I__10844 (
            .O(N__45650),
            .I(N__45644));
    Span4Mux_v I__10843 (
            .O(N__45647),
            .I(N__45641));
    Odrv12 I__10842 (
            .O(N__45644),
            .I(\pid_alt.error_filt_22 ));
    Odrv4 I__10841 (
            .O(N__45641),
            .I(\pid_alt.error_filt_22 ));
    InMux I__10840 (
            .O(N__45636),
            .I(N__45619));
    InMux I__10839 (
            .O(N__45635),
            .I(N__45619));
    InMux I__10838 (
            .O(N__45634),
            .I(N__45619));
    InMux I__10837 (
            .O(N__45633),
            .I(N__45619));
    InMux I__10836 (
            .O(N__45632),
            .I(N__45608));
    InMux I__10835 (
            .O(N__45631),
            .I(N__45608));
    InMux I__10834 (
            .O(N__45630),
            .I(N__45608));
    InMux I__10833 (
            .O(N__45629),
            .I(N__45608));
    InMux I__10832 (
            .O(N__45628),
            .I(N__45608));
    LocalMux I__10831 (
            .O(N__45619),
            .I(N__45603));
    LocalMux I__10830 (
            .O(N__45608),
            .I(N__45603));
    Odrv4 I__10829 (
            .O(N__45603),
            .I(\pid_alt.error_filt_prevZ0Z_22 ));
    InMux I__10828 (
            .O(N__45600),
            .I(N__45597));
    LocalMux I__10827 (
            .O(N__45597),
            .I(N__45593));
    InMux I__10826 (
            .O(N__45596),
            .I(N__45590));
    Sp12to4 I__10825 (
            .O(N__45593),
            .I(N__45587));
    LocalMux I__10824 (
            .O(N__45590),
            .I(N__45584));
    Span12Mux_v I__10823 (
            .O(N__45587),
            .I(N__45581));
    Span4Mux_v I__10822 (
            .O(N__45584),
            .I(N__45578));
    Span12Mux_h I__10821 (
            .O(N__45581),
            .I(N__45575));
    Span4Mux_v I__10820 (
            .O(N__45578),
            .I(N__45572));
    Odrv12 I__10819 (
            .O(N__45575),
            .I(\pid_alt.error_filt_20 ));
    Odrv4 I__10818 (
            .O(N__45572),
            .I(\pid_alt.error_filt_20 ));
    InMux I__10817 (
            .O(N__45567),
            .I(N__45564));
    LocalMux I__10816 (
            .O(N__45564),
            .I(\pid_alt.error_filt_prevZ0Z_20 ));
    InMux I__10815 (
            .O(N__45561),
            .I(N__45558));
    LocalMux I__10814 (
            .O(N__45558),
            .I(N__45554));
    InMux I__10813 (
            .O(N__45557),
            .I(N__45551));
    Span12Mux_h I__10812 (
            .O(N__45554),
            .I(N__45548));
    LocalMux I__10811 (
            .O(N__45551),
            .I(N__45545));
    Span12Mux_h I__10810 (
            .O(N__45548),
            .I(N__45542));
    Span4Mux_v I__10809 (
            .O(N__45545),
            .I(N__45539));
    Odrv12 I__10808 (
            .O(N__45542),
            .I(\pid_alt.error_filt_8 ));
    Odrv4 I__10807 (
            .O(N__45539),
            .I(\pid_alt.error_filt_8 ));
    InMux I__10806 (
            .O(N__45534),
            .I(N__45531));
    LocalMux I__10805 (
            .O(N__45531),
            .I(N__45528));
    Span4Mux_v I__10804 (
            .O(N__45528),
            .I(N__45525));
    Odrv4 I__10803 (
            .O(N__45525),
            .I(\pid_alt.error_filt_prevZ0Z_8 ));
    InMux I__10802 (
            .O(N__45522),
            .I(N__45519));
    LocalMux I__10801 (
            .O(N__45519),
            .I(N__45516));
    Span4Mux_v I__10800 (
            .O(N__45516),
            .I(N__45513));
    Span4Mux_h I__10799 (
            .O(N__45513),
            .I(N__45510));
    Span4Mux_h I__10798 (
            .O(N__45510),
            .I(N__45507));
    Span4Mux_h I__10797 (
            .O(N__45507),
            .I(N__45504));
    Span4Mux_h I__10796 (
            .O(N__45504),
            .I(N__45501));
    Span4Mux_h I__10795 (
            .O(N__45501),
            .I(N__45498));
    Odrv4 I__10794 (
            .O(N__45498),
            .I(\pid_alt.O_8 ));
    InMux I__10793 (
            .O(N__45495),
            .I(N__45490));
    InMux I__10792 (
            .O(N__45494),
            .I(N__45485));
    InMux I__10791 (
            .O(N__45493),
            .I(N__45485));
    LocalMux I__10790 (
            .O(N__45490),
            .I(N__45482));
    LocalMux I__10789 (
            .O(N__45485),
            .I(N__45479));
    Span4Mux_v I__10788 (
            .O(N__45482),
            .I(N__45476));
    Span4Mux_v I__10787 (
            .O(N__45479),
            .I(N__45473));
    Sp12to4 I__10786 (
            .O(N__45476),
            .I(N__45468));
    Sp12to4 I__10785 (
            .O(N__45473),
            .I(N__45468));
    Span12Mux_h I__10784 (
            .O(N__45468),
            .I(N__45465));
    Odrv12 I__10783 (
            .O(N__45465),
            .I(\pid_alt.error_d_regZ0Z_4 ));
    InMux I__10782 (
            .O(N__45462),
            .I(N__45459));
    LocalMux I__10781 (
            .O(N__45459),
            .I(N__45456));
    Span4Mux_v I__10780 (
            .O(N__45456),
            .I(N__45453));
    Span4Mux_h I__10779 (
            .O(N__45453),
            .I(N__45449));
    InMux I__10778 (
            .O(N__45452),
            .I(N__45446));
    Sp12to4 I__10777 (
            .O(N__45449),
            .I(N__45443));
    LocalMux I__10776 (
            .O(N__45446),
            .I(N__45440));
    Span12Mux_h I__10775 (
            .O(N__45443),
            .I(N__45437));
    Span4Mux_s1_h I__10774 (
            .O(N__45440),
            .I(N__45434));
    Odrv12 I__10773 (
            .O(N__45437),
            .I(\pid_alt.error_filt_1 ));
    Odrv4 I__10772 (
            .O(N__45434),
            .I(\pid_alt.error_filt_1 ));
    InMux I__10771 (
            .O(N__45429),
            .I(N__45426));
    LocalMux I__10770 (
            .O(N__45426),
            .I(N__45423));
    Odrv4 I__10769 (
            .O(N__45423),
            .I(\pid_alt.error_filt_prevZ0Z_1 ));
    InMux I__10768 (
            .O(N__45420),
            .I(N__45417));
    LocalMux I__10767 (
            .O(N__45417),
            .I(N__45414));
    Span4Mux_h I__10766 (
            .O(N__45414),
            .I(N__45411));
    Odrv4 I__10765 (
            .O(N__45411),
            .I(\pid_alt.O_0_9 ));
    InMux I__10764 (
            .O(N__45408),
            .I(N__45405));
    LocalMux I__10763 (
            .O(N__45405),
            .I(N__45402));
    Span12Mux_h I__10762 (
            .O(N__45402),
            .I(N__45399));
    Odrv12 I__10761 (
            .O(N__45399),
            .I(\pid_alt.error_i_regZ0Z_5 ));
    InMux I__10760 (
            .O(N__45396),
            .I(N__45393));
    LocalMux I__10759 (
            .O(N__45393),
            .I(N__45390));
    Span4Mux_v I__10758 (
            .O(N__45390),
            .I(N__45387));
    Odrv4 I__10757 (
            .O(N__45387),
            .I(\pid_alt.O_0_12 ));
    CascadeMux I__10756 (
            .O(N__45384),
            .I(N__45381));
    InMux I__10755 (
            .O(N__45381),
            .I(N__45378));
    LocalMux I__10754 (
            .O(N__45378),
            .I(N__45375));
    Span4Mux_h I__10753 (
            .O(N__45375),
            .I(N__45372));
    Span4Mux_h I__10752 (
            .O(N__45372),
            .I(N__45369));
    Odrv4 I__10751 (
            .O(N__45369),
            .I(\pid_alt.error_i_regZ0Z_8 ));
    InMux I__10750 (
            .O(N__45366),
            .I(N__45363));
    LocalMux I__10749 (
            .O(N__45363),
            .I(N__45359));
    InMux I__10748 (
            .O(N__45362),
            .I(N__45355));
    Span4Mux_h I__10747 (
            .O(N__45359),
            .I(N__45352));
    InMux I__10746 (
            .O(N__45358),
            .I(N__45347));
    LocalMux I__10745 (
            .O(N__45355),
            .I(N__45344));
    Span4Mux_h I__10744 (
            .O(N__45352),
            .I(N__45341));
    CascadeMux I__10743 (
            .O(N__45351),
            .I(N__45338));
    InMux I__10742 (
            .O(N__45350),
            .I(N__45335));
    LocalMux I__10741 (
            .O(N__45347),
            .I(N__45332));
    Span4Mux_v I__10740 (
            .O(N__45344),
            .I(N__45327));
    Span4Mux_h I__10739 (
            .O(N__45341),
            .I(N__45324));
    InMux I__10738 (
            .O(N__45338),
            .I(N__45321));
    LocalMux I__10737 (
            .O(N__45335),
            .I(N__45318));
    Span4Mux_v I__10736 (
            .O(N__45332),
            .I(N__45315));
    InMux I__10735 (
            .O(N__45331),
            .I(N__45310));
    InMux I__10734 (
            .O(N__45330),
            .I(N__45307));
    Span4Mux_h I__10733 (
            .O(N__45327),
            .I(N__45302));
    Span4Mux_v I__10732 (
            .O(N__45324),
            .I(N__45302));
    LocalMux I__10731 (
            .O(N__45321),
            .I(N__45299));
    Span4Mux_v I__10730 (
            .O(N__45318),
            .I(N__45293));
    Span4Mux_v I__10729 (
            .O(N__45315),
            .I(N__45290));
    InMux I__10728 (
            .O(N__45314),
            .I(N__45287));
    InMux I__10727 (
            .O(N__45313),
            .I(N__45284));
    LocalMux I__10726 (
            .O(N__45310),
            .I(N__45275));
    LocalMux I__10725 (
            .O(N__45307),
            .I(N__45275));
    Span4Mux_v I__10724 (
            .O(N__45302),
            .I(N__45275));
    Span4Mux_h I__10723 (
            .O(N__45299),
            .I(N__45275));
    InMux I__10722 (
            .O(N__45298),
            .I(N__45271));
    InMux I__10721 (
            .O(N__45297),
            .I(N__45268));
    InMux I__10720 (
            .O(N__45296),
            .I(N__45265));
    Span4Mux_h I__10719 (
            .O(N__45293),
            .I(N__45260));
    Span4Mux_v I__10718 (
            .O(N__45290),
            .I(N__45260));
    LocalMux I__10717 (
            .O(N__45287),
            .I(N__45253));
    LocalMux I__10716 (
            .O(N__45284),
            .I(N__45253));
    Span4Mux_v I__10715 (
            .O(N__45275),
            .I(N__45253));
    InMux I__10714 (
            .O(N__45274),
            .I(N__45250));
    LocalMux I__10713 (
            .O(N__45271),
            .I(uart_pc_data_4));
    LocalMux I__10712 (
            .O(N__45268),
            .I(uart_pc_data_4));
    LocalMux I__10711 (
            .O(N__45265),
            .I(uart_pc_data_4));
    Odrv4 I__10710 (
            .O(N__45260),
            .I(uart_pc_data_4));
    Odrv4 I__10709 (
            .O(N__45253),
            .I(uart_pc_data_4));
    LocalMux I__10708 (
            .O(N__45250),
            .I(uart_pc_data_4));
    InMux I__10707 (
            .O(N__45237),
            .I(N__45234));
    LocalMux I__10706 (
            .O(N__45234),
            .I(N__45231));
    Span4Mux_s3_h I__10705 (
            .O(N__45231),
            .I(N__45228));
    Odrv4 I__10704 (
            .O(N__45228),
            .I(alt_ki_4));
    InMux I__10703 (
            .O(N__45225),
            .I(N__45221));
    InMux I__10702 (
            .O(N__45224),
            .I(N__45218));
    LocalMux I__10701 (
            .O(N__45221),
            .I(N__45215));
    LocalMux I__10700 (
            .O(N__45218),
            .I(N__45208));
    Span4Mux_h I__10699 (
            .O(N__45215),
            .I(N__45205));
    InMux I__10698 (
            .O(N__45214),
            .I(N__45201));
    InMux I__10697 (
            .O(N__45213),
            .I(N__45197));
    InMux I__10696 (
            .O(N__45212),
            .I(N__45194));
    InMux I__10695 (
            .O(N__45211),
            .I(N__45191));
    Span4Mux_h I__10694 (
            .O(N__45208),
            .I(N__45187));
    Span4Mux_h I__10693 (
            .O(N__45205),
            .I(N__45183));
    InMux I__10692 (
            .O(N__45204),
            .I(N__45180));
    LocalMux I__10691 (
            .O(N__45201),
            .I(N__45177));
    InMux I__10690 (
            .O(N__45200),
            .I(N__45173));
    LocalMux I__10689 (
            .O(N__45197),
            .I(N__45168));
    LocalMux I__10688 (
            .O(N__45194),
            .I(N__45168));
    LocalMux I__10687 (
            .O(N__45191),
            .I(N__45165));
    InMux I__10686 (
            .O(N__45190),
            .I(N__45162));
    Sp12to4 I__10685 (
            .O(N__45187),
            .I(N__45158));
    InMux I__10684 (
            .O(N__45186),
            .I(N__45155));
    Span4Mux_v I__10683 (
            .O(N__45183),
            .I(N__45150));
    LocalMux I__10682 (
            .O(N__45180),
            .I(N__45150));
    Span4Mux_h I__10681 (
            .O(N__45177),
            .I(N__45147));
    InMux I__10680 (
            .O(N__45176),
            .I(N__45144));
    LocalMux I__10679 (
            .O(N__45173),
            .I(N__45141));
    Span4Mux_v I__10678 (
            .O(N__45168),
            .I(N__45134));
    Span4Mux_h I__10677 (
            .O(N__45165),
            .I(N__45134));
    LocalMux I__10676 (
            .O(N__45162),
            .I(N__45134));
    InMux I__10675 (
            .O(N__45161),
            .I(N__45131));
    Span12Mux_v I__10674 (
            .O(N__45158),
            .I(N__45127));
    LocalMux I__10673 (
            .O(N__45155),
            .I(N__45124));
    Span4Mux_h I__10672 (
            .O(N__45150),
            .I(N__45121));
    Span4Mux_v I__10671 (
            .O(N__45147),
            .I(N__45118));
    LocalMux I__10670 (
            .O(N__45144),
            .I(N__45115));
    Span12Mux_h I__10669 (
            .O(N__45141),
            .I(N__45112));
    Span4Mux_v I__10668 (
            .O(N__45134),
            .I(N__45109));
    LocalMux I__10667 (
            .O(N__45131),
            .I(N__45106));
    InMux I__10666 (
            .O(N__45130),
            .I(N__45103));
    Span12Mux_h I__10665 (
            .O(N__45127),
            .I(N__45096));
    Span12Mux_h I__10664 (
            .O(N__45124),
            .I(N__45096));
    Sp12to4 I__10663 (
            .O(N__45121),
            .I(N__45096));
    Span4Mux_v I__10662 (
            .O(N__45118),
            .I(N__45091));
    Span4Mux_h I__10661 (
            .O(N__45115),
            .I(N__45091));
    Odrv12 I__10660 (
            .O(N__45112),
            .I(uart_pc_data_1));
    Odrv4 I__10659 (
            .O(N__45109),
            .I(uart_pc_data_1));
    Odrv4 I__10658 (
            .O(N__45106),
            .I(uart_pc_data_1));
    LocalMux I__10657 (
            .O(N__45103),
            .I(uart_pc_data_1));
    Odrv12 I__10656 (
            .O(N__45096),
            .I(uart_pc_data_1));
    Odrv4 I__10655 (
            .O(N__45091),
            .I(uart_pc_data_1));
    InMux I__10654 (
            .O(N__45078),
            .I(N__45075));
    LocalMux I__10653 (
            .O(N__45075),
            .I(N__45072));
    Span4Mux_v I__10652 (
            .O(N__45072),
            .I(N__45069));
    Odrv4 I__10651 (
            .O(N__45069),
            .I(alt_ki_1));
    InMux I__10650 (
            .O(N__45066),
            .I(N__45063));
    LocalMux I__10649 (
            .O(N__45063),
            .I(N__45060));
    Span4Mux_h I__10648 (
            .O(N__45060),
            .I(N__45057));
    Span4Mux_h I__10647 (
            .O(N__45057),
            .I(N__45054));
    Span4Mux_h I__10646 (
            .O(N__45054),
            .I(N__45051));
    Span4Mux_h I__10645 (
            .O(N__45051),
            .I(N__45047));
    InMux I__10644 (
            .O(N__45050),
            .I(N__45044));
    Span4Mux_h I__10643 (
            .O(N__45047),
            .I(N__45041));
    LocalMux I__10642 (
            .O(N__45044),
            .I(N__45038));
    Span4Mux_h I__10641 (
            .O(N__45041),
            .I(N__45033));
    Span4Mux_v I__10640 (
            .O(N__45038),
            .I(N__45033));
    Span4Mux_v I__10639 (
            .O(N__45033),
            .I(N__45030));
    Odrv4 I__10638 (
            .O(N__45030),
            .I(\pid_alt.error_filt_19 ));
    InMux I__10637 (
            .O(N__45027),
            .I(N__45024));
    LocalMux I__10636 (
            .O(N__45024),
            .I(N__45021));
    Span4Mux_s2_h I__10635 (
            .O(N__45021),
            .I(N__45018));
    Odrv4 I__10634 (
            .O(N__45018),
            .I(\pid_alt.error_filt_prevZ0Z_19 ));
    InMux I__10633 (
            .O(N__45015),
            .I(N__45009));
    InMux I__10632 (
            .O(N__45014),
            .I(N__45006));
    InMux I__10631 (
            .O(N__45013),
            .I(N__45002));
    InMux I__10630 (
            .O(N__45012),
            .I(N__44998));
    LocalMux I__10629 (
            .O(N__45009),
            .I(N__44995));
    LocalMux I__10628 (
            .O(N__45006),
            .I(N__44992));
    InMux I__10627 (
            .O(N__45005),
            .I(N__44989));
    LocalMux I__10626 (
            .O(N__45002),
            .I(N__44985));
    InMux I__10625 (
            .O(N__45001),
            .I(N__44979));
    LocalMux I__10624 (
            .O(N__44998),
            .I(N__44976));
    Span4Mux_v I__10623 (
            .O(N__44995),
            .I(N__44973));
    Span4Mux_h I__10622 (
            .O(N__44992),
            .I(N__44970));
    LocalMux I__10621 (
            .O(N__44989),
            .I(N__44967));
    InMux I__10620 (
            .O(N__44988),
            .I(N__44964));
    Span4Mux_v I__10619 (
            .O(N__44985),
            .I(N__44961));
    InMux I__10618 (
            .O(N__44984),
            .I(N__44958));
    InMux I__10617 (
            .O(N__44983),
            .I(N__44955));
    InMux I__10616 (
            .O(N__44982),
            .I(N__44950));
    LocalMux I__10615 (
            .O(N__44979),
            .I(N__44947));
    Sp12to4 I__10614 (
            .O(N__44976),
            .I(N__44941));
    Sp12to4 I__10613 (
            .O(N__44973),
            .I(N__44941));
    Sp12to4 I__10612 (
            .O(N__44970),
            .I(N__44934));
    Sp12to4 I__10611 (
            .O(N__44967),
            .I(N__44934));
    LocalMux I__10610 (
            .O(N__44964),
            .I(N__44934));
    Sp12to4 I__10609 (
            .O(N__44961),
            .I(N__44931));
    LocalMux I__10608 (
            .O(N__44958),
            .I(N__44926));
    LocalMux I__10607 (
            .O(N__44955),
            .I(N__44926));
    InMux I__10606 (
            .O(N__44954),
            .I(N__44923));
    InMux I__10605 (
            .O(N__44953),
            .I(N__44920));
    LocalMux I__10604 (
            .O(N__44950),
            .I(N__44915));
    Span4Mux_h I__10603 (
            .O(N__44947),
            .I(N__44915));
    InMux I__10602 (
            .O(N__44946),
            .I(N__44911));
    Span12Mux_v I__10601 (
            .O(N__44941),
            .I(N__44908));
    Span12Mux_v I__10600 (
            .O(N__44934),
            .I(N__44903));
    Span12Mux_v I__10599 (
            .O(N__44931),
            .I(N__44903));
    Span4Mux_v I__10598 (
            .O(N__44926),
            .I(N__44898));
    LocalMux I__10597 (
            .O(N__44923),
            .I(N__44898));
    LocalMux I__10596 (
            .O(N__44920),
            .I(N__44893));
    Span4Mux_v I__10595 (
            .O(N__44915),
            .I(N__44893));
    InMux I__10594 (
            .O(N__44914),
            .I(N__44890));
    LocalMux I__10593 (
            .O(N__44911),
            .I(uart_pc_data_7));
    Odrv12 I__10592 (
            .O(N__44908),
            .I(uart_pc_data_7));
    Odrv12 I__10591 (
            .O(N__44903),
            .I(uart_pc_data_7));
    Odrv4 I__10590 (
            .O(N__44898),
            .I(uart_pc_data_7));
    Odrv4 I__10589 (
            .O(N__44893),
            .I(uart_pc_data_7));
    LocalMux I__10588 (
            .O(N__44890),
            .I(uart_pc_data_7));
    InMux I__10587 (
            .O(N__44877),
            .I(N__44874));
    LocalMux I__10586 (
            .O(N__44874),
            .I(N__44871));
    Span4Mux_v I__10585 (
            .O(N__44871),
            .I(N__44868));
    Odrv4 I__10584 (
            .O(N__44868),
            .I(alt_ki_7));
    CEMux I__10583 (
            .O(N__44865),
            .I(N__44861));
    CEMux I__10582 (
            .O(N__44864),
            .I(N__44857));
    LocalMux I__10581 (
            .O(N__44861),
            .I(N__44853));
    CEMux I__10580 (
            .O(N__44860),
            .I(N__44850));
    LocalMux I__10579 (
            .O(N__44857),
            .I(N__44846));
    CEMux I__10578 (
            .O(N__44856),
            .I(N__44843));
    Span4Mux_v I__10577 (
            .O(N__44853),
            .I(N__44838));
    LocalMux I__10576 (
            .O(N__44850),
            .I(N__44838));
    CEMux I__10575 (
            .O(N__44849),
            .I(N__44835));
    Span4Mux_v I__10574 (
            .O(N__44846),
            .I(N__44832));
    LocalMux I__10573 (
            .O(N__44843),
            .I(N__44829));
    Span4Mux_h I__10572 (
            .O(N__44838),
            .I(N__44825));
    LocalMux I__10571 (
            .O(N__44835),
            .I(N__44822));
    Span4Mux_h I__10570 (
            .O(N__44832),
            .I(N__44816));
    Span4Mux_h I__10569 (
            .O(N__44829),
            .I(N__44816));
    CEMux I__10568 (
            .O(N__44828),
            .I(N__44813));
    Span4Mux_h I__10567 (
            .O(N__44825),
            .I(N__44808));
    Span4Mux_v I__10566 (
            .O(N__44822),
            .I(N__44808));
    CEMux I__10565 (
            .O(N__44821),
            .I(N__44805));
    Span4Mux_h I__10564 (
            .O(N__44816),
            .I(N__44800));
    LocalMux I__10563 (
            .O(N__44813),
            .I(N__44800));
    Span4Mux_h I__10562 (
            .O(N__44808),
            .I(N__44795));
    LocalMux I__10561 (
            .O(N__44805),
            .I(N__44795));
    Span4Mux_v I__10560 (
            .O(N__44800),
            .I(N__44792));
    Span4Mux_h I__10559 (
            .O(N__44795),
            .I(N__44789));
    Sp12to4 I__10558 (
            .O(N__44792),
            .I(N__44786));
    Span4Mux_v I__10557 (
            .O(N__44789),
            .I(N__44783));
    Span12Mux_h I__10556 (
            .O(N__44786),
            .I(N__44780));
    Span4Mux_v I__10555 (
            .O(N__44783),
            .I(N__44777));
    Odrv12 I__10554 (
            .O(N__44780),
            .I(\Commands_frame_decoder.state_RNIQRI31Z0Z_10 ));
    Odrv4 I__10553 (
            .O(N__44777),
            .I(\Commands_frame_decoder.state_RNIQRI31Z0Z_10 ));
    InMux I__10552 (
            .O(N__44772),
            .I(N__44769));
    LocalMux I__10551 (
            .O(N__44769),
            .I(N__44766));
    Span4Mux_h I__10550 (
            .O(N__44766),
            .I(N__44763));
    Odrv4 I__10549 (
            .O(N__44763),
            .I(\pid_alt.O_0_14 ));
    CascadeMux I__10548 (
            .O(N__44760),
            .I(N__44757));
    InMux I__10547 (
            .O(N__44757),
            .I(N__44754));
    LocalMux I__10546 (
            .O(N__44754),
            .I(N__44751));
    Span4Mux_v I__10545 (
            .O(N__44751),
            .I(N__44748));
    Span4Mux_h I__10544 (
            .O(N__44748),
            .I(N__44745));
    Span4Mux_h I__10543 (
            .O(N__44745),
            .I(N__44742));
    Odrv4 I__10542 (
            .O(N__44742),
            .I(\pid_alt.error_i_regZ0Z_10 ));
    InMux I__10541 (
            .O(N__44739),
            .I(N__44736));
    LocalMux I__10540 (
            .O(N__44736),
            .I(N__44733));
    Span4Mux_h I__10539 (
            .O(N__44733),
            .I(N__44730));
    Odrv4 I__10538 (
            .O(N__44730),
            .I(\pid_alt.O_15 ));
    CascadeMux I__10537 (
            .O(N__44727),
            .I(N__44724));
    InMux I__10536 (
            .O(N__44724),
            .I(N__44721));
    LocalMux I__10535 (
            .O(N__44721),
            .I(N__44718));
    Span4Mux_v I__10534 (
            .O(N__44718),
            .I(N__44715));
    Span4Mux_h I__10533 (
            .O(N__44715),
            .I(N__44712));
    Span4Mux_h I__10532 (
            .O(N__44712),
            .I(N__44709));
    Odrv4 I__10531 (
            .O(N__44709),
            .I(\pid_alt.error_i_regZ0Z_11 ));
    InMux I__10530 (
            .O(N__44706),
            .I(N__44703));
    LocalMux I__10529 (
            .O(N__44703),
            .I(N__44700));
    Span4Mux_h I__10528 (
            .O(N__44700),
            .I(N__44697));
    Odrv4 I__10527 (
            .O(N__44697),
            .I(\pid_alt.O_16 ));
    CascadeMux I__10526 (
            .O(N__44694),
            .I(N__44691));
    InMux I__10525 (
            .O(N__44691),
            .I(N__44688));
    LocalMux I__10524 (
            .O(N__44688),
            .I(N__44685));
    Span4Mux_v I__10523 (
            .O(N__44685),
            .I(N__44682));
    Span4Mux_h I__10522 (
            .O(N__44682),
            .I(N__44679));
    Span4Mux_h I__10521 (
            .O(N__44679),
            .I(N__44676));
    Odrv4 I__10520 (
            .O(N__44676),
            .I(\pid_alt.error_i_regZ0Z_12 ));
    InMux I__10519 (
            .O(N__44673),
            .I(\ppm_encoder_1.counter24_0_N_2 ));
    InMux I__10518 (
            .O(N__44670),
            .I(N__44667));
    LocalMux I__10517 (
            .O(N__44667),
            .I(N__44662));
    InMux I__10516 (
            .O(N__44666),
            .I(N__44656));
    InMux I__10515 (
            .O(N__44665),
            .I(N__44656));
    Span4Mux_h I__10514 (
            .O(N__44662),
            .I(N__44653));
    InMux I__10513 (
            .O(N__44661),
            .I(N__44650));
    LocalMux I__10512 (
            .O(N__44656),
            .I(N__44647));
    Span4Mux_v I__10511 (
            .O(N__44653),
            .I(N__44642));
    LocalMux I__10510 (
            .O(N__44650),
            .I(N__44642));
    Span4Mux_v I__10509 (
            .O(N__44647),
            .I(N__44639));
    Odrv4 I__10508 (
            .O(N__44642),
            .I(\ppm_encoder_1.counter24_0_N_2_THRU_CO ));
    Odrv4 I__10507 (
            .O(N__44639),
            .I(\ppm_encoder_1.counter24_0_N_2_THRU_CO ));
    InMux I__10506 (
            .O(N__44634),
            .I(N__44631));
    LocalMux I__10505 (
            .O(N__44631),
            .I(N__44628));
    Odrv4 I__10504 (
            .O(N__44628),
            .I(\ppm_encoder_1.pulses2countZ0Z_10 ));
    InMux I__10503 (
            .O(N__44625),
            .I(N__44622));
    LocalMux I__10502 (
            .O(N__44622),
            .I(N__44617));
    InMux I__10501 (
            .O(N__44621),
            .I(N__44614));
    InMux I__10500 (
            .O(N__44620),
            .I(N__44611));
    Span4Mux_h I__10499 (
            .O(N__44617),
            .I(N__44608));
    LocalMux I__10498 (
            .O(N__44614),
            .I(\ppm_encoder_1.counterZ0Z_11 ));
    LocalMux I__10497 (
            .O(N__44611),
            .I(\ppm_encoder_1.counterZ0Z_11 ));
    Odrv4 I__10496 (
            .O(N__44608),
            .I(\ppm_encoder_1.counterZ0Z_11 ));
    CascadeMux I__10495 (
            .O(N__44601),
            .I(N__44598));
    InMux I__10494 (
            .O(N__44598),
            .I(N__44595));
    LocalMux I__10493 (
            .O(N__44595),
            .I(N__44592));
    Odrv4 I__10492 (
            .O(N__44592),
            .I(\ppm_encoder_1.pulses2countZ0Z_11 ));
    InMux I__10491 (
            .O(N__44589),
            .I(N__44586));
    LocalMux I__10490 (
            .O(N__44586),
            .I(N__44581));
    InMux I__10489 (
            .O(N__44585),
            .I(N__44578));
    InMux I__10488 (
            .O(N__44584),
            .I(N__44575));
    Span4Mux_h I__10487 (
            .O(N__44581),
            .I(N__44572));
    LocalMux I__10486 (
            .O(N__44578),
            .I(\ppm_encoder_1.counterZ0Z_10 ));
    LocalMux I__10485 (
            .O(N__44575),
            .I(\ppm_encoder_1.counterZ0Z_10 ));
    Odrv4 I__10484 (
            .O(N__44572),
            .I(\ppm_encoder_1.counterZ0Z_10 ));
    CascadeMux I__10483 (
            .O(N__44565),
            .I(N__44562));
    InMux I__10482 (
            .O(N__44562),
            .I(N__44559));
    LocalMux I__10481 (
            .O(N__44559),
            .I(\ppm_encoder_1.counter24_0_I_33_c_RNOZ0 ));
    InMux I__10480 (
            .O(N__44556),
            .I(N__44553));
    LocalMux I__10479 (
            .O(N__44553),
            .I(N__44549));
    CascadeMux I__10478 (
            .O(N__44552),
            .I(N__44545));
    Span4Mux_h I__10477 (
            .O(N__44549),
            .I(N__44542));
    InMux I__10476 (
            .O(N__44548),
            .I(N__44532));
    InMux I__10475 (
            .O(N__44545),
            .I(N__44532));
    Span4Mux_h I__10474 (
            .O(N__44542),
            .I(N__44529));
    InMux I__10473 (
            .O(N__44541),
            .I(N__44526));
    InMux I__10472 (
            .O(N__44540),
            .I(N__44523));
    InMux I__10471 (
            .O(N__44539),
            .I(N__44520));
    InMux I__10470 (
            .O(N__44538),
            .I(N__44515));
    InMux I__10469 (
            .O(N__44537),
            .I(N__44515));
    LocalMux I__10468 (
            .O(N__44532),
            .I(N__44512));
    Odrv4 I__10467 (
            .O(N__44529),
            .I(\uart_drone.stateZ0Z_3 ));
    LocalMux I__10466 (
            .O(N__44526),
            .I(\uart_drone.stateZ0Z_3 ));
    LocalMux I__10465 (
            .O(N__44523),
            .I(\uart_drone.stateZ0Z_3 ));
    LocalMux I__10464 (
            .O(N__44520),
            .I(\uart_drone.stateZ0Z_3 ));
    LocalMux I__10463 (
            .O(N__44515),
            .I(\uart_drone.stateZ0Z_3 ));
    Odrv4 I__10462 (
            .O(N__44512),
            .I(\uart_drone.stateZ0Z_3 ));
    CascadeMux I__10461 (
            .O(N__44499),
            .I(N__44496));
    InMux I__10460 (
            .O(N__44496),
            .I(N__44492));
    CascadeMux I__10459 (
            .O(N__44495),
            .I(N__44489));
    LocalMux I__10458 (
            .O(N__44492),
            .I(N__44486));
    InMux I__10457 (
            .O(N__44489),
            .I(N__44482));
    Span4Mux_h I__10456 (
            .O(N__44486),
            .I(N__44479));
    InMux I__10455 (
            .O(N__44485),
            .I(N__44476));
    LocalMux I__10454 (
            .O(N__44482),
            .I(\uart_drone.un1_state_4_0 ));
    Odrv4 I__10453 (
            .O(N__44479),
            .I(\uart_drone.un1_state_4_0 ));
    LocalMux I__10452 (
            .O(N__44476),
            .I(\uart_drone.un1_state_4_0 ));
    InMux I__10451 (
            .O(N__44469),
            .I(N__44465));
    InMux I__10450 (
            .O(N__44468),
            .I(N__44462));
    LocalMux I__10449 (
            .O(N__44465),
            .I(N__44458));
    LocalMux I__10448 (
            .O(N__44462),
            .I(N__44455));
    InMux I__10447 (
            .O(N__44461),
            .I(N__44452));
    Span4Mux_v I__10446 (
            .O(N__44458),
            .I(N__44448));
    Span4Mux_v I__10445 (
            .O(N__44455),
            .I(N__44445));
    LocalMux I__10444 (
            .O(N__44452),
            .I(N__44442));
    InMux I__10443 (
            .O(N__44451),
            .I(N__44439));
    Span4Mux_h I__10442 (
            .O(N__44448),
            .I(N__44436));
    Span4Mux_h I__10441 (
            .O(N__44445),
            .I(N__44429));
    Span4Mux_v I__10440 (
            .O(N__44442),
            .I(N__44429));
    LocalMux I__10439 (
            .O(N__44439),
            .I(N__44429));
    Odrv4 I__10438 (
            .O(N__44436),
            .I(\uart_drone.N_152 ));
    Odrv4 I__10437 (
            .O(N__44429),
            .I(\uart_drone.N_152 ));
    InMux I__10436 (
            .O(N__44424),
            .I(N__44415));
    InMux I__10435 (
            .O(N__44423),
            .I(N__44415));
    InMux I__10434 (
            .O(N__44422),
            .I(N__44410));
    InMux I__10433 (
            .O(N__44421),
            .I(N__44410));
    InMux I__10432 (
            .O(N__44420),
            .I(N__44407));
    LocalMux I__10431 (
            .O(N__44415),
            .I(N__44398));
    LocalMux I__10430 (
            .O(N__44410),
            .I(N__44398));
    LocalMux I__10429 (
            .O(N__44407),
            .I(N__44398));
    InMux I__10428 (
            .O(N__44406),
            .I(N__44393));
    InMux I__10427 (
            .O(N__44405),
            .I(N__44393));
    Span4Mux_v I__10426 (
            .O(N__44398),
            .I(N__44386));
    LocalMux I__10425 (
            .O(N__44393),
            .I(N__44386));
    InMux I__10424 (
            .O(N__44392),
            .I(N__44383));
    InMux I__10423 (
            .O(N__44391),
            .I(N__44379));
    Span4Mux_h I__10422 (
            .O(N__44386),
            .I(N__44375));
    LocalMux I__10421 (
            .O(N__44383),
            .I(N__44372));
    InMux I__10420 (
            .O(N__44382),
            .I(N__44369));
    LocalMux I__10419 (
            .O(N__44379),
            .I(N__44366));
    InMux I__10418 (
            .O(N__44378),
            .I(N__44363));
    Span4Mux_h I__10417 (
            .O(N__44375),
            .I(N__44360));
    Span4Mux_v I__10416 (
            .O(N__44372),
            .I(N__44355));
    LocalMux I__10415 (
            .O(N__44369),
            .I(N__44355));
    Span12Mux_h I__10414 (
            .O(N__44366),
            .I(N__44352));
    LocalMux I__10413 (
            .O(N__44363),
            .I(\uart_drone.bit_CountZ0Z_0 ));
    Odrv4 I__10412 (
            .O(N__44360),
            .I(\uart_drone.bit_CountZ0Z_0 ));
    Odrv4 I__10411 (
            .O(N__44355),
            .I(\uart_drone.bit_CountZ0Z_0 ));
    Odrv12 I__10410 (
            .O(N__44352),
            .I(\uart_drone.bit_CountZ0Z_0 ));
    InMux I__10409 (
            .O(N__44343),
            .I(N__44340));
    LocalMux I__10408 (
            .O(N__44340),
            .I(N__44337));
    Span4Mux_h I__10407 (
            .O(N__44337),
            .I(N__44334));
    Span4Mux_h I__10406 (
            .O(N__44334),
            .I(N__44331));
    Span4Mux_h I__10405 (
            .O(N__44331),
            .I(N__44327));
    InMux I__10404 (
            .O(N__44330),
            .I(N__44324));
    Span4Mux_h I__10403 (
            .O(N__44327),
            .I(N__44321));
    LocalMux I__10402 (
            .O(N__44324),
            .I(N__44318));
    Span4Mux_h I__10401 (
            .O(N__44321),
            .I(N__44313));
    Span4Mux_v I__10400 (
            .O(N__44318),
            .I(N__44313));
    Span4Mux_v I__10399 (
            .O(N__44313),
            .I(N__44310));
    Odrv4 I__10398 (
            .O(N__44310),
            .I(\pid_alt.error_filt_21 ));
    InMux I__10397 (
            .O(N__44307),
            .I(N__44304));
    LocalMux I__10396 (
            .O(N__44304),
            .I(N__44301));
    Span4Mux_s0_h I__10395 (
            .O(N__44301),
            .I(N__44298));
    Span4Mux_h I__10394 (
            .O(N__44298),
            .I(N__44295));
    Odrv4 I__10393 (
            .O(N__44295),
            .I(\pid_alt.error_filt_prevZ0Z_21 ));
    InMux I__10392 (
            .O(N__44292),
            .I(N__44287));
    InMux I__10391 (
            .O(N__44291),
            .I(N__44284));
    InMux I__10390 (
            .O(N__44290),
            .I(N__44280));
    LocalMux I__10389 (
            .O(N__44287),
            .I(N__44275));
    LocalMux I__10388 (
            .O(N__44284),
            .I(N__44275));
    InMux I__10387 (
            .O(N__44283),
            .I(N__44272));
    LocalMux I__10386 (
            .O(N__44280),
            .I(N__44267));
    Span4Mux_v I__10385 (
            .O(N__44275),
            .I(N__44264));
    LocalMux I__10384 (
            .O(N__44272),
            .I(N__44259));
    CascadeMux I__10383 (
            .O(N__44271),
            .I(N__44255));
    InMux I__10382 (
            .O(N__44270),
            .I(N__44251));
    Span4Mux_v I__10381 (
            .O(N__44267),
            .I(N__44244));
    Span4Mux_h I__10380 (
            .O(N__44264),
            .I(N__44244));
    InMux I__10379 (
            .O(N__44263),
            .I(N__44241));
    InMux I__10378 (
            .O(N__44262),
            .I(N__44237));
    Span4Mux_v I__10377 (
            .O(N__44259),
            .I(N__44234));
    InMux I__10376 (
            .O(N__44258),
            .I(N__44227));
    InMux I__10375 (
            .O(N__44255),
            .I(N__44227));
    InMux I__10374 (
            .O(N__44254),
            .I(N__44227));
    LocalMux I__10373 (
            .O(N__44251),
            .I(N__44224));
    InMux I__10372 (
            .O(N__44250),
            .I(N__44221));
    InMux I__10371 (
            .O(N__44249),
            .I(N__44218));
    Span4Mux_v I__10370 (
            .O(N__44244),
            .I(N__44213));
    LocalMux I__10369 (
            .O(N__44241),
            .I(N__44213));
    InMux I__10368 (
            .O(N__44240),
            .I(N__44210));
    LocalMux I__10367 (
            .O(N__44237),
            .I(N__44207));
    Sp12to4 I__10366 (
            .O(N__44234),
            .I(N__44202));
    LocalMux I__10365 (
            .O(N__44227),
            .I(N__44199));
    Span4Mux_v I__10364 (
            .O(N__44224),
            .I(N__44190));
    LocalMux I__10363 (
            .O(N__44221),
            .I(N__44190));
    LocalMux I__10362 (
            .O(N__44218),
            .I(N__44190));
    Span4Mux_h I__10361 (
            .O(N__44213),
            .I(N__44190));
    LocalMux I__10360 (
            .O(N__44210),
            .I(N__44187));
    Span4Mux_h I__10359 (
            .O(N__44207),
            .I(N__44184));
    InMux I__10358 (
            .O(N__44206),
            .I(N__44181));
    InMux I__10357 (
            .O(N__44205),
            .I(N__44178));
    Span12Mux_v I__10356 (
            .O(N__44202),
            .I(N__44175));
    Span4Mux_h I__10355 (
            .O(N__44199),
            .I(N__44172));
    Span4Mux_v I__10354 (
            .O(N__44190),
            .I(N__44169));
    Odrv12 I__10353 (
            .O(N__44187),
            .I(uart_pc_data_5));
    Odrv4 I__10352 (
            .O(N__44184),
            .I(uart_pc_data_5));
    LocalMux I__10351 (
            .O(N__44181),
            .I(uart_pc_data_5));
    LocalMux I__10350 (
            .O(N__44178),
            .I(uart_pc_data_5));
    Odrv12 I__10349 (
            .O(N__44175),
            .I(uart_pc_data_5));
    Odrv4 I__10348 (
            .O(N__44172),
            .I(uart_pc_data_5));
    Odrv4 I__10347 (
            .O(N__44169),
            .I(uart_pc_data_5));
    InMux I__10346 (
            .O(N__44154),
            .I(N__44151));
    LocalMux I__10345 (
            .O(N__44151),
            .I(N__44148));
    Span4Mux_s0_h I__10344 (
            .O(N__44148),
            .I(N__44145));
    Span4Mux_h I__10343 (
            .O(N__44145),
            .I(N__44142));
    Odrv4 I__10342 (
            .O(N__44142),
            .I(alt_ki_5));
    CascadeMux I__10341 (
            .O(N__44139),
            .I(N__44132));
    CascadeMux I__10340 (
            .O(N__44138),
            .I(N__44129));
    CascadeMux I__10339 (
            .O(N__44137),
            .I(N__44119));
    CascadeMux I__10338 (
            .O(N__44136),
            .I(N__44113));
    CascadeMux I__10337 (
            .O(N__44135),
            .I(N__44093));
    InMux I__10336 (
            .O(N__44132),
            .I(N__44060));
    InMux I__10335 (
            .O(N__44129),
            .I(N__44060));
    InMux I__10334 (
            .O(N__44128),
            .I(N__44057));
    InMux I__10333 (
            .O(N__44127),
            .I(N__44052));
    InMux I__10332 (
            .O(N__44126),
            .I(N__44052));
    InMux I__10331 (
            .O(N__44125),
            .I(N__44049));
    InMux I__10330 (
            .O(N__44124),
            .I(N__44046));
    InMux I__10329 (
            .O(N__44123),
            .I(N__44043));
    InMux I__10328 (
            .O(N__44122),
            .I(N__44040));
    InMux I__10327 (
            .O(N__44119),
            .I(N__44037));
    InMux I__10326 (
            .O(N__44118),
            .I(N__44034));
    InMux I__10325 (
            .O(N__44117),
            .I(N__44031));
    InMux I__10324 (
            .O(N__44116),
            .I(N__44022));
    InMux I__10323 (
            .O(N__44113),
            .I(N__44022));
    InMux I__10322 (
            .O(N__44112),
            .I(N__44022));
    InMux I__10321 (
            .O(N__44111),
            .I(N__44022));
    InMux I__10320 (
            .O(N__44110),
            .I(N__44019));
    InMux I__10319 (
            .O(N__44109),
            .I(N__44014));
    InMux I__10318 (
            .O(N__44108),
            .I(N__44014));
    InMux I__10317 (
            .O(N__44107),
            .I(N__44009));
    InMux I__10316 (
            .O(N__44106),
            .I(N__44009));
    InMux I__10315 (
            .O(N__44105),
            .I(N__44004));
    InMux I__10314 (
            .O(N__44104),
            .I(N__44004));
    InMux I__10313 (
            .O(N__44103),
            .I(N__43999));
    InMux I__10312 (
            .O(N__44102),
            .I(N__43999));
    InMux I__10311 (
            .O(N__44101),
            .I(N__43996));
    InMux I__10310 (
            .O(N__44100),
            .I(N__43993));
    InMux I__10309 (
            .O(N__44099),
            .I(N__43990));
    InMux I__10308 (
            .O(N__44098),
            .I(N__43983));
    InMux I__10307 (
            .O(N__44097),
            .I(N__43983));
    InMux I__10306 (
            .O(N__44096),
            .I(N__43983));
    InMux I__10305 (
            .O(N__44093),
            .I(N__43980));
    InMux I__10304 (
            .O(N__44092),
            .I(N__43977));
    InMux I__10303 (
            .O(N__44091),
            .I(N__43974));
    InMux I__10302 (
            .O(N__44090),
            .I(N__43971));
    InMux I__10301 (
            .O(N__44089),
            .I(N__43968));
    InMux I__10300 (
            .O(N__44088),
            .I(N__43965));
    InMux I__10299 (
            .O(N__44087),
            .I(N__43960));
    InMux I__10298 (
            .O(N__44086),
            .I(N__43960));
    InMux I__10297 (
            .O(N__44085),
            .I(N__43957));
    InMux I__10296 (
            .O(N__44084),
            .I(N__43954));
    InMux I__10295 (
            .O(N__44083),
            .I(N__43951));
    InMux I__10294 (
            .O(N__44082),
            .I(N__43948));
    InMux I__10293 (
            .O(N__44081),
            .I(N__43941));
    InMux I__10292 (
            .O(N__44080),
            .I(N__43941));
    InMux I__10291 (
            .O(N__44079),
            .I(N__43941));
    InMux I__10290 (
            .O(N__44078),
            .I(N__43938));
    InMux I__10289 (
            .O(N__44077),
            .I(N__43933));
    InMux I__10288 (
            .O(N__44076),
            .I(N__43933));
    InMux I__10287 (
            .O(N__44075),
            .I(N__43930));
    InMux I__10286 (
            .O(N__44074),
            .I(N__43927));
    InMux I__10285 (
            .O(N__44073),
            .I(N__43922));
    InMux I__10284 (
            .O(N__44072),
            .I(N__43922));
    InMux I__10283 (
            .O(N__44071),
            .I(N__43919));
    InMux I__10282 (
            .O(N__44070),
            .I(N__43916));
    InMux I__10281 (
            .O(N__44069),
            .I(N__43913));
    InMux I__10280 (
            .O(N__44068),
            .I(N__43908));
    InMux I__10279 (
            .O(N__44067),
            .I(N__43908));
    InMux I__10278 (
            .O(N__44066),
            .I(N__43905));
    InMux I__10277 (
            .O(N__44065),
            .I(N__43902));
    LocalMux I__10276 (
            .O(N__44060),
            .I(N__43796));
    LocalMux I__10275 (
            .O(N__44057),
            .I(N__43793));
    LocalMux I__10274 (
            .O(N__44052),
            .I(N__43790));
    LocalMux I__10273 (
            .O(N__44049),
            .I(N__43787));
    LocalMux I__10272 (
            .O(N__44046),
            .I(N__43784));
    LocalMux I__10271 (
            .O(N__44043),
            .I(N__43781));
    LocalMux I__10270 (
            .O(N__44040),
            .I(N__43778));
    LocalMux I__10269 (
            .O(N__44037),
            .I(N__43775));
    LocalMux I__10268 (
            .O(N__44034),
            .I(N__43772));
    LocalMux I__10267 (
            .O(N__44031),
            .I(N__43769));
    LocalMux I__10266 (
            .O(N__44022),
            .I(N__43766));
    LocalMux I__10265 (
            .O(N__44019),
            .I(N__43763));
    LocalMux I__10264 (
            .O(N__44014),
            .I(N__43760));
    LocalMux I__10263 (
            .O(N__44009),
            .I(N__43757));
    LocalMux I__10262 (
            .O(N__44004),
            .I(N__43754));
    LocalMux I__10261 (
            .O(N__43999),
            .I(N__43751));
    LocalMux I__10260 (
            .O(N__43996),
            .I(N__43748));
    LocalMux I__10259 (
            .O(N__43993),
            .I(N__43745));
    LocalMux I__10258 (
            .O(N__43990),
            .I(N__43742));
    LocalMux I__10257 (
            .O(N__43983),
            .I(N__43739));
    LocalMux I__10256 (
            .O(N__43980),
            .I(N__43736));
    LocalMux I__10255 (
            .O(N__43977),
            .I(N__43733));
    LocalMux I__10254 (
            .O(N__43974),
            .I(N__43730));
    LocalMux I__10253 (
            .O(N__43971),
            .I(N__43727));
    LocalMux I__10252 (
            .O(N__43968),
            .I(N__43724));
    LocalMux I__10251 (
            .O(N__43965),
            .I(N__43721));
    LocalMux I__10250 (
            .O(N__43960),
            .I(N__43718));
    LocalMux I__10249 (
            .O(N__43957),
            .I(N__43715));
    LocalMux I__10248 (
            .O(N__43954),
            .I(N__43712));
    LocalMux I__10247 (
            .O(N__43951),
            .I(N__43709));
    LocalMux I__10246 (
            .O(N__43948),
            .I(N__43706));
    LocalMux I__10245 (
            .O(N__43941),
            .I(N__43703));
    LocalMux I__10244 (
            .O(N__43938),
            .I(N__43700));
    LocalMux I__10243 (
            .O(N__43933),
            .I(N__43697));
    LocalMux I__10242 (
            .O(N__43930),
            .I(N__43694));
    LocalMux I__10241 (
            .O(N__43927),
            .I(N__43691));
    LocalMux I__10240 (
            .O(N__43922),
            .I(N__43688));
    LocalMux I__10239 (
            .O(N__43919),
            .I(N__43685));
    LocalMux I__10238 (
            .O(N__43916),
            .I(N__43682));
    LocalMux I__10237 (
            .O(N__43913),
            .I(N__43679));
    LocalMux I__10236 (
            .O(N__43908),
            .I(N__43676));
    LocalMux I__10235 (
            .O(N__43905),
            .I(N__43673));
    LocalMux I__10234 (
            .O(N__43902),
            .I(N__43670));
    SRMux I__10233 (
            .O(N__43901),
            .I(N__43377));
    SRMux I__10232 (
            .O(N__43900),
            .I(N__43377));
    SRMux I__10231 (
            .O(N__43899),
            .I(N__43377));
    SRMux I__10230 (
            .O(N__43898),
            .I(N__43377));
    SRMux I__10229 (
            .O(N__43897),
            .I(N__43377));
    SRMux I__10228 (
            .O(N__43896),
            .I(N__43377));
    SRMux I__10227 (
            .O(N__43895),
            .I(N__43377));
    SRMux I__10226 (
            .O(N__43894),
            .I(N__43377));
    SRMux I__10225 (
            .O(N__43893),
            .I(N__43377));
    SRMux I__10224 (
            .O(N__43892),
            .I(N__43377));
    SRMux I__10223 (
            .O(N__43891),
            .I(N__43377));
    SRMux I__10222 (
            .O(N__43890),
            .I(N__43377));
    SRMux I__10221 (
            .O(N__43889),
            .I(N__43377));
    SRMux I__10220 (
            .O(N__43888),
            .I(N__43377));
    SRMux I__10219 (
            .O(N__43887),
            .I(N__43377));
    SRMux I__10218 (
            .O(N__43886),
            .I(N__43377));
    SRMux I__10217 (
            .O(N__43885),
            .I(N__43377));
    SRMux I__10216 (
            .O(N__43884),
            .I(N__43377));
    SRMux I__10215 (
            .O(N__43883),
            .I(N__43377));
    SRMux I__10214 (
            .O(N__43882),
            .I(N__43377));
    SRMux I__10213 (
            .O(N__43881),
            .I(N__43377));
    SRMux I__10212 (
            .O(N__43880),
            .I(N__43377));
    SRMux I__10211 (
            .O(N__43879),
            .I(N__43377));
    SRMux I__10210 (
            .O(N__43878),
            .I(N__43377));
    SRMux I__10209 (
            .O(N__43877),
            .I(N__43377));
    SRMux I__10208 (
            .O(N__43876),
            .I(N__43377));
    SRMux I__10207 (
            .O(N__43875),
            .I(N__43377));
    SRMux I__10206 (
            .O(N__43874),
            .I(N__43377));
    SRMux I__10205 (
            .O(N__43873),
            .I(N__43377));
    SRMux I__10204 (
            .O(N__43872),
            .I(N__43377));
    SRMux I__10203 (
            .O(N__43871),
            .I(N__43377));
    SRMux I__10202 (
            .O(N__43870),
            .I(N__43377));
    SRMux I__10201 (
            .O(N__43869),
            .I(N__43377));
    SRMux I__10200 (
            .O(N__43868),
            .I(N__43377));
    SRMux I__10199 (
            .O(N__43867),
            .I(N__43377));
    SRMux I__10198 (
            .O(N__43866),
            .I(N__43377));
    SRMux I__10197 (
            .O(N__43865),
            .I(N__43377));
    SRMux I__10196 (
            .O(N__43864),
            .I(N__43377));
    SRMux I__10195 (
            .O(N__43863),
            .I(N__43377));
    SRMux I__10194 (
            .O(N__43862),
            .I(N__43377));
    SRMux I__10193 (
            .O(N__43861),
            .I(N__43377));
    SRMux I__10192 (
            .O(N__43860),
            .I(N__43377));
    SRMux I__10191 (
            .O(N__43859),
            .I(N__43377));
    SRMux I__10190 (
            .O(N__43858),
            .I(N__43377));
    SRMux I__10189 (
            .O(N__43857),
            .I(N__43377));
    SRMux I__10188 (
            .O(N__43856),
            .I(N__43377));
    SRMux I__10187 (
            .O(N__43855),
            .I(N__43377));
    SRMux I__10186 (
            .O(N__43854),
            .I(N__43377));
    SRMux I__10185 (
            .O(N__43853),
            .I(N__43377));
    SRMux I__10184 (
            .O(N__43852),
            .I(N__43377));
    SRMux I__10183 (
            .O(N__43851),
            .I(N__43377));
    SRMux I__10182 (
            .O(N__43850),
            .I(N__43377));
    SRMux I__10181 (
            .O(N__43849),
            .I(N__43377));
    SRMux I__10180 (
            .O(N__43848),
            .I(N__43377));
    SRMux I__10179 (
            .O(N__43847),
            .I(N__43377));
    SRMux I__10178 (
            .O(N__43846),
            .I(N__43377));
    SRMux I__10177 (
            .O(N__43845),
            .I(N__43377));
    SRMux I__10176 (
            .O(N__43844),
            .I(N__43377));
    SRMux I__10175 (
            .O(N__43843),
            .I(N__43377));
    SRMux I__10174 (
            .O(N__43842),
            .I(N__43377));
    SRMux I__10173 (
            .O(N__43841),
            .I(N__43377));
    SRMux I__10172 (
            .O(N__43840),
            .I(N__43377));
    SRMux I__10171 (
            .O(N__43839),
            .I(N__43377));
    SRMux I__10170 (
            .O(N__43838),
            .I(N__43377));
    SRMux I__10169 (
            .O(N__43837),
            .I(N__43377));
    SRMux I__10168 (
            .O(N__43836),
            .I(N__43377));
    SRMux I__10167 (
            .O(N__43835),
            .I(N__43377));
    SRMux I__10166 (
            .O(N__43834),
            .I(N__43377));
    SRMux I__10165 (
            .O(N__43833),
            .I(N__43377));
    SRMux I__10164 (
            .O(N__43832),
            .I(N__43377));
    SRMux I__10163 (
            .O(N__43831),
            .I(N__43377));
    SRMux I__10162 (
            .O(N__43830),
            .I(N__43377));
    SRMux I__10161 (
            .O(N__43829),
            .I(N__43377));
    SRMux I__10160 (
            .O(N__43828),
            .I(N__43377));
    SRMux I__10159 (
            .O(N__43827),
            .I(N__43377));
    SRMux I__10158 (
            .O(N__43826),
            .I(N__43377));
    SRMux I__10157 (
            .O(N__43825),
            .I(N__43377));
    SRMux I__10156 (
            .O(N__43824),
            .I(N__43377));
    SRMux I__10155 (
            .O(N__43823),
            .I(N__43377));
    SRMux I__10154 (
            .O(N__43822),
            .I(N__43377));
    SRMux I__10153 (
            .O(N__43821),
            .I(N__43377));
    SRMux I__10152 (
            .O(N__43820),
            .I(N__43377));
    SRMux I__10151 (
            .O(N__43819),
            .I(N__43377));
    SRMux I__10150 (
            .O(N__43818),
            .I(N__43377));
    SRMux I__10149 (
            .O(N__43817),
            .I(N__43377));
    SRMux I__10148 (
            .O(N__43816),
            .I(N__43377));
    SRMux I__10147 (
            .O(N__43815),
            .I(N__43377));
    SRMux I__10146 (
            .O(N__43814),
            .I(N__43377));
    SRMux I__10145 (
            .O(N__43813),
            .I(N__43377));
    SRMux I__10144 (
            .O(N__43812),
            .I(N__43377));
    SRMux I__10143 (
            .O(N__43811),
            .I(N__43377));
    SRMux I__10142 (
            .O(N__43810),
            .I(N__43377));
    SRMux I__10141 (
            .O(N__43809),
            .I(N__43377));
    SRMux I__10140 (
            .O(N__43808),
            .I(N__43377));
    SRMux I__10139 (
            .O(N__43807),
            .I(N__43377));
    SRMux I__10138 (
            .O(N__43806),
            .I(N__43377));
    SRMux I__10137 (
            .O(N__43805),
            .I(N__43377));
    SRMux I__10136 (
            .O(N__43804),
            .I(N__43377));
    SRMux I__10135 (
            .O(N__43803),
            .I(N__43377));
    SRMux I__10134 (
            .O(N__43802),
            .I(N__43377));
    SRMux I__10133 (
            .O(N__43801),
            .I(N__43377));
    SRMux I__10132 (
            .O(N__43800),
            .I(N__43377));
    SRMux I__10131 (
            .O(N__43799),
            .I(N__43377));
    Glb2LocalMux I__10130 (
            .O(N__43796),
            .I(N__43377));
    Glb2LocalMux I__10129 (
            .O(N__43793),
            .I(N__43377));
    Glb2LocalMux I__10128 (
            .O(N__43790),
            .I(N__43377));
    Glb2LocalMux I__10127 (
            .O(N__43787),
            .I(N__43377));
    Glb2LocalMux I__10126 (
            .O(N__43784),
            .I(N__43377));
    Glb2LocalMux I__10125 (
            .O(N__43781),
            .I(N__43377));
    Glb2LocalMux I__10124 (
            .O(N__43778),
            .I(N__43377));
    Glb2LocalMux I__10123 (
            .O(N__43775),
            .I(N__43377));
    Glb2LocalMux I__10122 (
            .O(N__43772),
            .I(N__43377));
    Glb2LocalMux I__10121 (
            .O(N__43769),
            .I(N__43377));
    Glb2LocalMux I__10120 (
            .O(N__43766),
            .I(N__43377));
    Glb2LocalMux I__10119 (
            .O(N__43763),
            .I(N__43377));
    Glb2LocalMux I__10118 (
            .O(N__43760),
            .I(N__43377));
    Glb2LocalMux I__10117 (
            .O(N__43757),
            .I(N__43377));
    Glb2LocalMux I__10116 (
            .O(N__43754),
            .I(N__43377));
    Glb2LocalMux I__10115 (
            .O(N__43751),
            .I(N__43377));
    Glb2LocalMux I__10114 (
            .O(N__43748),
            .I(N__43377));
    Glb2LocalMux I__10113 (
            .O(N__43745),
            .I(N__43377));
    Glb2LocalMux I__10112 (
            .O(N__43742),
            .I(N__43377));
    Glb2LocalMux I__10111 (
            .O(N__43739),
            .I(N__43377));
    Glb2LocalMux I__10110 (
            .O(N__43736),
            .I(N__43377));
    Glb2LocalMux I__10109 (
            .O(N__43733),
            .I(N__43377));
    Glb2LocalMux I__10108 (
            .O(N__43730),
            .I(N__43377));
    Glb2LocalMux I__10107 (
            .O(N__43727),
            .I(N__43377));
    Glb2LocalMux I__10106 (
            .O(N__43724),
            .I(N__43377));
    Glb2LocalMux I__10105 (
            .O(N__43721),
            .I(N__43377));
    Glb2LocalMux I__10104 (
            .O(N__43718),
            .I(N__43377));
    Glb2LocalMux I__10103 (
            .O(N__43715),
            .I(N__43377));
    Glb2LocalMux I__10102 (
            .O(N__43712),
            .I(N__43377));
    Glb2LocalMux I__10101 (
            .O(N__43709),
            .I(N__43377));
    Glb2LocalMux I__10100 (
            .O(N__43706),
            .I(N__43377));
    Glb2LocalMux I__10099 (
            .O(N__43703),
            .I(N__43377));
    Glb2LocalMux I__10098 (
            .O(N__43700),
            .I(N__43377));
    Glb2LocalMux I__10097 (
            .O(N__43697),
            .I(N__43377));
    Glb2LocalMux I__10096 (
            .O(N__43694),
            .I(N__43377));
    Glb2LocalMux I__10095 (
            .O(N__43691),
            .I(N__43377));
    Glb2LocalMux I__10094 (
            .O(N__43688),
            .I(N__43377));
    Glb2LocalMux I__10093 (
            .O(N__43685),
            .I(N__43377));
    Glb2LocalMux I__10092 (
            .O(N__43682),
            .I(N__43377));
    Glb2LocalMux I__10091 (
            .O(N__43679),
            .I(N__43377));
    Glb2LocalMux I__10090 (
            .O(N__43676),
            .I(N__43377));
    Glb2LocalMux I__10089 (
            .O(N__43673),
            .I(N__43377));
    Glb2LocalMux I__10088 (
            .O(N__43670),
            .I(N__43377));
    GlobalMux I__10087 (
            .O(N__43377),
            .I(N__43374));
    gio2CtrlBuf I__10086 (
            .O(N__43374),
            .I(reset_system_g));
    IoInMux I__10085 (
            .O(N__43371),
            .I(N__43368));
    LocalMux I__10084 (
            .O(N__43368),
            .I(GB_BUFFER_reset_system_g_THRU_CO));
    InMux I__10083 (
            .O(N__43365),
            .I(N__43361));
    InMux I__10082 (
            .O(N__43364),
            .I(N__43358));
    LocalMux I__10081 (
            .O(N__43361),
            .I(N__43355));
    LocalMux I__10080 (
            .O(N__43358),
            .I(N__43350));
    Span4Mux_v I__10079 (
            .O(N__43355),
            .I(N__43346));
    InMux I__10078 (
            .O(N__43354),
            .I(N__43343));
    InMux I__10077 (
            .O(N__43353),
            .I(N__43336));
    Span4Mux_v I__10076 (
            .O(N__43350),
            .I(N__43333));
    InMux I__10075 (
            .O(N__43349),
            .I(N__43330));
    Span4Mux_h I__10074 (
            .O(N__43346),
            .I(N__43325));
    LocalMux I__10073 (
            .O(N__43343),
            .I(N__43325));
    InMux I__10072 (
            .O(N__43342),
            .I(N__43322));
    InMux I__10071 (
            .O(N__43341),
            .I(N__43319));
    InMux I__10070 (
            .O(N__43340),
            .I(N__43316));
    InMux I__10069 (
            .O(N__43339),
            .I(N__43313));
    LocalMux I__10068 (
            .O(N__43336),
            .I(N__43309));
    Span4Mux_h I__10067 (
            .O(N__43333),
            .I(N__43305));
    LocalMux I__10066 (
            .O(N__43330),
            .I(N__43298));
    Span4Mux_h I__10065 (
            .O(N__43325),
            .I(N__43298));
    LocalMux I__10064 (
            .O(N__43322),
            .I(N__43298));
    LocalMux I__10063 (
            .O(N__43319),
            .I(N__43293));
    LocalMux I__10062 (
            .O(N__43316),
            .I(N__43293));
    LocalMux I__10061 (
            .O(N__43313),
            .I(N__43290));
    InMux I__10060 (
            .O(N__43312),
            .I(N__43287));
    Span4Mux_h I__10059 (
            .O(N__43309),
            .I(N__43283));
    InMux I__10058 (
            .O(N__43308),
            .I(N__43280));
    Span4Mux_h I__10057 (
            .O(N__43305),
            .I(N__43277));
    Span4Mux_v I__10056 (
            .O(N__43298),
            .I(N__43274));
    Span4Mux_v I__10055 (
            .O(N__43293),
            .I(N__43267));
    Span4Mux_h I__10054 (
            .O(N__43290),
            .I(N__43267));
    LocalMux I__10053 (
            .O(N__43287),
            .I(N__43267));
    InMux I__10052 (
            .O(N__43286),
            .I(N__43263));
    Span4Mux_h I__10051 (
            .O(N__43283),
            .I(N__43258));
    LocalMux I__10050 (
            .O(N__43280),
            .I(N__43258));
    Span4Mux_v I__10049 (
            .O(N__43277),
            .I(N__43253));
    Span4Mux_h I__10048 (
            .O(N__43274),
            .I(N__43253));
    Span4Mux_v I__10047 (
            .O(N__43267),
            .I(N__43250));
    InMux I__10046 (
            .O(N__43266),
            .I(N__43247));
    LocalMux I__10045 (
            .O(N__43263),
            .I(N__43244));
    Span4Mux_h I__10044 (
            .O(N__43258),
            .I(N__43239));
    Span4Mux_v I__10043 (
            .O(N__43253),
            .I(N__43239));
    Odrv4 I__10042 (
            .O(N__43250),
            .I(uart_pc_data_3));
    LocalMux I__10041 (
            .O(N__43247),
            .I(uart_pc_data_3));
    Odrv12 I__10040 (
            .O(N__43244),
            .I(uart_pc_data_3));
    Odrv4 I__10039 (
            .O(N__43239),
            .I(uart_pc_data_3));
    InMux I__10038 (
            .O(N__43230),
            .I(N__43227));
    LocalMux I__10037 (
            .O(N__43227),
            .I(N__43224));
    Span4Mux_v I__10036 (
            .O(N__43224),
            .I(N__43221));
    Odrv4 I__10035 (
            .O(N__43221),
            .I(alt_ki_3));
    InMux I__10034 (
            .O(N__43218),
            .I(N__43215));
    LocalMux I__10033 (
            .O(N__43215),
            .I(N__43212));
    Span4Mux_h I__10032 (
            .O(N__43212),
            .I(N__43209));
    Odrv4 I__10031 (
            .O(N__43209),
            .I(\pid_alt.O_0_8 ));
    CascadeMux I__10030 (
            .O(N__43206),
            .I(N__43203));
    InMux I__10029 (
            .O(N__43203),
            .I(N__43200));
    LocalMux I__10028 (
            .O(N__43200),
            .I(N__43197));
    Span12Mux_h I__10027 (
            .O(N__43197),
            .I(N__43194));
    Odrv12 I__10026 (
            .O(N__43194),
            .I(\pid_alt.error_i_regZ0Z_4 ));
    InMux I__10025 (
            .O(N__43191),
            .I(N__43188));
    LocalMux I__10024 (
            .O(N__43188),
            .I(N__43185));
    Span4Mux_h I__10023 (
            .O(N__43185),
            .I(N__43182));
    Odrv4 I__10022 (
            .O(N__43182),
            .I(\ppm_encoder_1.counter24_0_I_15_c_RNOZ0 ));
    CascadeMux I__10021 (
            .O(N__43179),
            .I(N__43176));
    InMux I__10020 (
            .O(N__43176),
            .I(N__43173));
    LocalMux I__10019 (
            .O(N__43173),
            .I(N__43170));
    Odrv4 I__10018 (
            .O(N__43170),
            .I(\ppm_encoder_1.counter24_0_I_21_c_RNOZ0 ));
    InMux I__10017 (
            .O(N__43167),
            .I(N__43164));
    LocalMux I__10016 (
            .O(N__43164),
            .I(\ppm_encoder_1.counter24_0_I_27_c_RNOZ0 ));
    InMux I__10015 (
            .O(N__43161),
            .I(N__43158));
    LocalMux I__10014 (
            .O(N__43158),
            .I(\ppm_encoder_1.counter24_0_I_39_c_RNOZ0 ));
    CascadeMux I__10013 (
            .O(N__43155),
            .I(N__43152));
    InMux I__10012 (
            .O(N__43152),
            .I(N__43149));
    LocalMux I__10011 (
            .O(N__43149),
            .I(\ppm_encoder_1.counter24_0_I_45_c_RNOZ0 ));
    InMux I__10010 (
            .O(N__43146),
            .I(N__43143));
    LocalMux I__10009 (
            .O(N__43143),
            .I(\ppm_encoder_1.counter24_0_I_51_c_RNOZ0 ));
    InMux I__10008 (
            .O(N__43140),
            .I(N__43135));
    InMux I__10007 (
            .O(N__43139),
            .I(N__43132));
    InMux I__10006 (
            .O(N__43138),
            .I(N__43119));
    LocalMux I__10005 (
            .O(N__43135),
            .I(N__43111));
    LocalMux I__10004 (
            .O(N__43132),
            .I(N__43111));
    InMux I__10003 (
            .O(N__43131),
            .I(N__43107));
    InMux I__10002 (
            .O(N__43130),
            .I(N__43104));
    InMux I__10001 (
            .O(N__43129),
            .I(N__43101));
    InMux I__10000 (
            .O(N__43128),
            .I(N__43098));
    InMux I__9999 (
            .O(N__43127),
            .I(N__43093));
    InMux I__9998 (
            .O(N__43126),
            .I(N__43093));
    InMux I__9997 (
            .O(N__43125),
            .I(N__43088));
    InMux I__9996 (
            .O(N__43124),
            .I(N__43088));
    CascadeMux I__9995 (
            .O(N__43123),
            .I(N__43082));
    InMux I__9994 (
            .O(N__43122),
            .I(N__43078));
    LocalMux I__9993 (
            .O(N__43119),
            .I(N__43075));
    CascadeMux I__9992 (
            .O(N__43118),
            .I(N__43071));
    InMux I__9991 (
            .O(N__43117),
            .I(N__43065));
    InMux I__9990 (
            .O(N__43116),
            .I(N__43062));
    Span4Mux_v I__9989 (
            .O(N__43111),
            .I(N__43059));
    InMux I__9988 (
            .O(N__43110),
            .I(N__43056));
    LocalMux I__9987 (
            .O(N__43107),
            .I(N__43047));
    LocalMux I__9986 (
            .O(N__43104),
            .I(N__43042));
    LocalMux I__9985 (
            .O(N__43101),
            .I(N__43042));
    LocalMux I__9984 (
            .O(N__43098),
            .I(N__43035));
    LocalMux I__9983 (
            .O(N__43093),
            .I(N__43035));
    LocalMux I__9982 (
            .O(N__43088),
            .I(N__43035));
    InMux I__9981 (
            .O(N__43087),
            .I(N__43030));
    InMux I__9980 (
            .O(N__43086),
            .I(N__43030));
    InMux I__9979 (
            .O(N__43085),
            .I(N__43027));
    InMux I__9978 (
            .O(N__43082),
            .I(N__43024));
    CascadeMux I__9977 (
            .O(N__43081),
            .I(N__43021));
    LocalMux I__9976 (
            .O(N__43078),
            .I(N__43017));
    Span4Mux_s2_h I__9975 (
            .O(N__43075),
            .I(N__43014));
    InMux I__9974 (
            .O(N__43074),
            .I(N__43009));
    InMux I__9973 (
            .O(N__43071),
            .I(N__43009));
    CascadeMux I__9972 (
            .O(N__43070),
            .I(N__43004));
    CascadeMux I__9971 (
            .O(N__43069),
            .I(N__43000));
    CascadeMux I__9970 (
            .O(N__43068),
            .I(N__42996));
    LocalMux I__9969 (
            .O(N__43065),
            .I(N__42989));
    LocalMux I__9968 (
            .O(N__43062),
            .I(N__42989));
    Span4Mux_h I__9967 (
            .O(N__43059),
            .I(N__42984));
    LocalMux I__9966 (
            .O(N__43056),
            .I(N__42984));
    InMux I__9965 (
            .O(N__43055),
            .I(N__42979));
    InMux I__9964 (
            .O(N__43054),
            .I(N__42979));
    InMux I__9963 (
            .O(N__43053),
            .I(N__42976));
    InMux I__9962 (
            .O(N__43052),
            .I(N__42971));
    InMux I__9961 (
            .O(N__43051),
            .I(N__42971));
    CascadeMux I__9960 (
            .O(N__43050),
            .I(N__42968));
    Span4Mux_v I__9959 (
            .O(N__43047),
            .I(N__42963));
    Span4Mux_v I__9958 (
            .O(N__43042),
            .I(N__42963));
    Span4Mux_v I__9957 (
            .O(N__43035),
            .I(N__42956));
    LocalMux I__9956 (
            .O(N__43030),
            .I(N__42956));
    LocalMux I__9955 (
            .O(N__43027),
            .I(N__42956));
    LocalMux I__9954 (
            .O(N__43024),
            .I(N__42953));
    InMux I__9953 (
            .O(N__43021),
            .I(N__42950));
    CascadeMux I__9952 (
            .O(N__43020),
            .I(N__42947));
    Span4Mux_s3_h I__9951 (
            .O(N__43017),
            .I(N__42944));
    Span4Mux_h I__9950 (
            .O(N__43014),
            .I(N__42939));
    LocalMux I__9949 (
            .O(N__43009),
            .I(N__42939));
    InMux I__9948 (
            .O(N__43008),
            .I(N__42924));
    InMux I__9947 (
            .O(N__43007),
            .I(N__42924));
    InMux I__9946 (
            .O(N__43004),
            .I(N__42924));
    InMux I__9945 (
            .O(N__43003),
            .I(N__42924));
    InMux I__9944 (
            .O(N__43000),
            .I(N__42924));
    InMux I__9943 (
            .O(N__42999),
            .I(N__42924));
    InMux I__9942 (
            .O(N__42996),
            .I(N__42924));
    CascadeMux I__9941 (
            .O(N__42995),
            .I(N__42920));
    CascadeMux I__9940 (
            .O(N__42994),
            .I(N__42917));
    Span4Mux_v I__9939 (
            .O(N__42989),
            .I(N__42913));
    Span4Mux_v I__9938 (
            .O(N__42984),
            .I(N__42908));
    LocalMux I__9937 (
            .O(N__42979),
            .I(N__42908));
    LocalMux I__9936 (
            .O(N__42976),
            .I(N__42903));
    LocalMux I__9935 (
            .O(N__42971),
            .I(N__42903));
    InMux I__9934 (
            .O(N__42968),
            .I(N__42900));
    Span4Mux_v I__9933 (
            .O(N__42963),
            .I(N__42895));
    Span4Mux_v I__9932 (
            .O(N__42956),
            .I(N__42895));
    Span4Mux_v I__9931 (
            .O(N__42953),
            .I(N__42890));
    LocalMux I__9930 (
            .O(N__42950),
            .I(N__42890));
    InMux I__9929 (
            .O(N__42947),
            .I(N__42887));
    Span4Mux_v I__9928 (
            .O(N__42944),
            .I(N__42882));
    Span4Mux_v I__9927 (
            .O(N__42939),
            .I(N__42877));
    LocalMux I__9926 (
            .O(N__42924),
            .I(N__42877));
    InMux I__9925 (
            .O(N__42923),
            .I(N__42870));
    InMux I__9924 (
            .O(N__42920),
            .I(N__42870));
    InMux I__9923 (
            .O(N__42917),
            .I(N__42870));
    CascadeMux I__9922 (
            .O(N__42916),
            .I(N__42867));
    Span4Mux_v I__9921 (
            .O(N__42913),
            .I(N__42862));
    Span4Mux_v I__9920 (
            .O(N__42908),
            .I(N__42862));
    Span4Mux_v I__9919 (
            .O(N__42903),
            .I(N__42859));
    LocalMux I__9918 (
            .O(N__42900),
            .I(N__42856));
    Span4Mux_h I__9917 (
            .O(N__42895),
            .I(N__42853));
    Span4Mux_v I__9916 (
            .O(N__42890),
            .I(N__42848));
    LocalMux I__9915 (
            .O(N__42887),
            .I(N__42848));
    InMux I__9914 (
            .O(N__42886),
            .I(N__42845));
    CascadeMux I__9913 (
            .O(N__42885),
            .I(N__42842));
    Span4Mux_h I__9912 (
            .O(N__42882),
            .I(N__42838));
    Span4Mux_h I__9911 (
            .O(N__42877),
            .I(N__42835));
    LocalMux I__9910 (
            .O(N__42870),
            .I(N__42832));
    InMux I__9909 (
            .O(N__42867),
            .I(N__42829));
    Span4Mux_h I__9908 (
            .O(N__42862),
            .I(N__42824));
    Span4Mux_h I__9907 (
            .O(N__42859),
            .I(N__42824));
    Span4Mux_v I__9906 (
            .O(N__42856),
            .I(N__42821));
    Span4Mux_h I__9905 (
            .O(N__42853),
            .I(N__42816));
    Span4Mux_v I__9904 (
            .O(N__42848),
            .I(N__42816));
    LocalMux I__9903 (
            .O(N__42845),
            .I(N__42813));
    InMux I__9902 (
            .O(N__42842),
            .I(N__42810));
    CascadeMux I__9901 (
            .O(N__42841),
            .I(N__42807));
    Span4Mux_h I__9900 (
            .O(N__42838),
            .I(N__42802));
    Span4Mux_h I__9899 (
            .O(N__42835),
            .I(N__42802));
    Span4Mux_h I__9898 (
            .O(N__42832),
            .I(N__42797));
    LocalMux I__9897 (
            .O(N__42829),
            .I(N__42797));
    Span4Mux_h I__9896 (
            .O(N__42824),
            .I(N__42788));
    Span4Mux_h I__9895 (
            .O(N__42821),
            .I(N__42788));
    Span4Mux_h I__9894 (
            .O(N__42816),
            .I(N__42788));
    Span4Mux_v I__9893 (
            .O(N__42813),
            .I(N__42788));
    LocalMux I__9892 (
            .O(N__42810),
            .I(N__42785));
    InMux I__9891 (
            .O(N__42807),
            .I(N__42782));
    Odrv4 I__9890 (
            .O(N__42802),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__9889 (
            .O(N__42797),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__9888 (
            .O(N__42788),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__9887 (
            .O(N__42785),
            .I(CONSTANT_ONE_NET));
    LocalMux I__9886 (
            .O(N__42782),
            .I(CONSTANT_ONE_NET));
    CascadeMux I__9885 (
            .O(N__42771),
            .I(N__42768));
    InMux I__9884 (
            .O(N__42768),
            .I(N__42765));
    LocalMux I__9883 (
            .O(N__42765),
            .I(\ppm_encoder_1.counter24_0_I_57_c_RNOZ0 ));
    InMux I__9882 (
            .O(N__42762),
            .I(N__42759));
    LocalMux I__9881 (
            .O(N__42759),
            .I(N__42756));
    Span12Mux_v I__9880 (
            .O(N__42756),
            .I(N__42753));
    Odrv12 I__9879 (
            .O(N__42753),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_7 ));
    InMux I__9878 (
            .O(N__42750),
            .I(N__42747));
    LocalMux I__9877 (
            .O(N__42747),
            .I(N__42744));
    Odrv12 I__9876 (
            .O(N__42744),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_7 ));
    CascadeMux I__9875 (
            .O(N__42741),
            .I(N__42737));
    InMux I__9874 (
            .O(N__42740),
            .I(N__42733));
    InMux I__9873 (
            .O(N__42737),
            .I(N__42730));
    InMux I__9872 (
            .O(N__42736),
            .I(N__42727));
    LocalMux I__9871 (
            .O(N__42733),
            .I(N__42720));
    LocalMux I__9870 (
            .O(N__42730),
            .I(N__42720));
    LocalMux I__9869 (
            .O(N__42727),
            .I(N__42720));
    Odrv4 I__9868 (
            .O(N__42720),
            .I(\ppm_encoder_1.counterZ0Z_7 ));
    CascadeMux I__9867 (
            .O(N__42717),
            .I(N__42714));
    InMux I__9866 (
            .O(N__42714),
            .I(N__42711));
    LocalMux I__9865 (
            .O(N__42711),
            .I(\ppm_encoder_1.pulses2countZ0Z_7 ));
    InMux I__9864 (
            .O(N__42708),
            .I(N__42703));
    InMux I__9863 (
            .O(N__42707),
            .I(N__42700));
    InMux I__9862 (
            .O(N__42706),
            .I(N__42697));
    LocalMux I__9861 (
            .O(N__42703),
            .I(N__42692));
    LocalMux I__9860 (
            .O(N__42700),
            .I(N__42692));
    LocalMux I__9859 (
            .O(N__42697),
            .I(\ppm_encoder_1.counterZ0Z_6 ));
    Odrv4 I__9858 (
            .O(N__42692),
            .I(\ppm_encoder_1.counterZ0Z_6 ));
    InMux I__9857 (
            .O(N__42687),
            .I(N__42684));
    LocalMux I__9856 (
            .O(N__42684),
            .I(N__42681));
    Span4Mux_v I__9855 (
            .O(N__42681),
            .I(N__42678));
    Span4Mux_h I__9854 (
            .O(N__42678),
            .I(N__42675));
    Odrv4 I__9853 (
            .O(N__42675),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_6 ));
    InMux I__9852 (
            .O(N__42672),
            .I(N__42669));
    LocalMux I__9851 (
            .O(N__42669),
            .I(N__42666));
    Span4Mux_h I__9850 (
            .O(N__42666),
            .I(N__42663));
    Odrv4 I__9849 (
            .O(N__42663),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_6 ));
    InMux I__9848 (
            .O(N__42660),
            .I(N__42657));
    LocalMux I__9847 (
            .O(N__42657),
            .I(\ppm_encoder_1.pulses2countZ0Z_6 ));
    InMux I__9846 (
            .O(N__42654),
            .I(N__42651));
    LocalMux I__9845 (
            .O(N__42651),
            .I(N__42648));
    Span4Mux_h I__9844 (
            .O(N__42648),
            .I(N__42645));
    Odrv4 I__9843 (
            .O(N__42645),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_11 ));
    InMux I__9842 (
            .O(N__42642),
            .I(N__42639));
    LocalMux I__9841 (
            .O(N__42639),
            .I(N__42636));
    Span4Mux_v I__9840 (
            .O(N__42636),
            .I(N__42633));
    Odrv4 I__9839 (
            .O(N__42633),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_11 ));
    InMux I__9838 (
            .O(N__42630),
            .I(N__42627));
    LocalMux I__9837 (
            .O(N__42627),
            .I(N__42624));
    Span4Mux_h I__9836 (
            .O(N__42624),
            .I(N__42621));
    Odrv4 I__9835 (
            .O(N__42621),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_12 ));
    CascadeMux I__9834 (
            .O(N__42618),
            .I(N__42613));
    CascadeMux I__9833 (
            .O(N__42617),
            .I(N__42600));
    InMux I__9832 (
            .O(N__42616),
            .I(N__42591));
    InMux I__9831 (
            .O(N__42613),
            .I(N__42591));
    InMux I__9830 (
            .O(N__42612),
            .I(N__42591));
    InMux I__9829 (
            .O(N__42611),
            .I(N__42580));
    InMux I__9828 (
            .O(N__42610),
            .I(N__42580));
    InMux I__9827 (
            .O(N__42609),
            .I(N__42580));
    InMux I__9826 (
            .O(N__42608),
            .I(N__42580));
    InMux I__9825 (
            .O(N__42607),
            .I(N__42580));
    InMux I__9824 (
            .O(N__42606),
            .I(N__42573));
    InMux I__9823 (
            .O(N__42605),
            .I(N__42573));
    InMux I__9822 (
            .O(N__42604),
            .I(N__42573));
    InMux I__9821 (
            .O(N__42603),
            .I(N__42564));
    InMux I__9820 (
            .O(N__42600),
            .I(N__42564));
    InMux I__9819 (
            .O(N__42599),
            .I(N__42564));
    InMux I__9818 (
            .O(N__42598),
            .I(N__42564));
    LocalMux I__9817 (
            .O(N__42591),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_11_mux ));
    LocalMux I__9816 (
            .O(N__42580),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_11_mux ));
    LocalMux I__9815 (
            .O(N__42573),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_11_mux ));
    LocalMux I__9814 (
            .O(N__42564),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_11_mux ));
    InMux I__9813 (
            .O(N__42555),
            .I(N__42552));
    LocalMux I__9812 (
            .O(N__42552),
            .I(N__42549));
    Span4Mux_v I__9811 (
            .O(N__42549),
            .I(N__42546));
    Span4Mux_h I__9810 (
            .O(N__42546),
            .I(N__42543));
    Odrv4 I__9809 (
            .O(N__42543),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_12 ));
    CEMux I__9808 (
            .O(N__42540),
            .I(N__42535));
    CEMux I__9807 (
            .O(N__42539),
            .I(N__42532));
    CEMux I__9806 (
            .O(N__42538),
            .I(N__42528));
    LocalMux I__9805 (
            .O(N__42535),
            .I(N__42525));
    LocalMux I__9804 (
            .O(N__42532),
            .I(N__42522));
    CEMux I__9803 (
            .O(N__42531),
            .I(N__42519));
    LocalMux I__9802 (
            .O(N__42528),
            .I(N__42516));
    Span4Mux_v I__9801 (
            .O(N__42525),
            .I(N__42513));
    Span4Mux_v I__9800 (
            .O(N__42522),
            .I(N__42510));
    LocalMux I__9799 (
            .O(N__42519),
            .I(N__42507));
    Span4Mux_h I__9798 (
            .O(N__42516),
            .I(N__42504));
    Span4Mux_h I__9797 (
            .O(N__42513),
            .I(N__42501));
    Span4Mux_h I__9796 (
            .O(N__42510),
            .I(N__42496));
    Span4Mux_h I__9795 (
            .O(N__42507),
            .I(N__42496));
    Odrv4 I__9794 (
            .O(N__42504),
            .I(\ppm_encoder_1.N_1330_0 ));
    Odrv4 I__9793 (
            .O(N__42501),
            .I(\ppm_encoder_1.N_1330_0 ));
    Odrv4 I__9792 (
            .O(N__42496),
            .I(\ppm_encoder_1.N_1330_0 ));
    InMux I__9791 (
            .O(N__42489),
            .I(N__42486));
    LocalMux I__9790 (
            .O(N__42486),
            .I(N__42481));
    InMux I__9789 (
            .O(N__42485),
            .I(N__42478));
    InMux I__9788 (
            .O(N__42484),
            .I(N__42475));
    Span4Mux_h I__9787 (
            .O(N__42481),
            .I(N__42472));
    LocalMux I__9786 (
            .O(N__42478),
            .I(\ppm_encoder_1.counterZ0Z_13 ));
    LocalMux I__9785 (
            .O(N__42475),
            .I(\ppm_encoder_1.counterZ0Z_13 ));
    Odrv4 I__9784 (
            .O(N__42472),
            .I(\ppm_encoder_1.counterZ0Z_13 ));
    InMux I__9783 (
            .O(N__42465),
            .I(N__42462));
    LocalMux I__9782 (
            .O(N__42462),
            .I(\ppm_encoder_1.pulses2countZ0Z_12 ));
    CascadeMux I__9781 (
            .O(N__42459),
            .I(N__42456));
    InMux I__9780 (
            .O(N__42456),
            .I(N__42453));
    LocalMux I__9779 (
            .O(N__42453),
            .I(\ppm_encoder_1.pulses2countZ0Z_13 ));
    InMux I__9778 (
            .O(N__42450),
            .I(N__42447));
    LocalMux I__9777 (
            .O(N__42447),
            .I(N__42442));
    InMux I__9776 (
            .O(N__42446),
            .I(N__42439));
    InMux I__9775 (
            .O(N__42445),
            .I(N__42436));
    Span4Mux_h I__9774 (
            .O(N__42442),
            .I(N__42433));
    LocalMux I__9773 (
            .O(N__42439),
            .I(\ppm_encoder_1.counterZ0Z_12 ));
    LocalMux I__9772 (
            .O(N__42436),
            .I(\ppm_encoder_1.counterZ0Z_12 ));
    Odrv4 I__9771 (
            .O(N__42433),
            .I(\ppm_encoder_1.counterZ0Z_12 ));
    InMux I__9770 (
            .O(N__42426),
            .I(N__42423));
    LocalMux I__9769 (
            .O(N__42423),
            .I(N__42420));
    Odrv4 I__9768 (
            .O(N__42420),
            .I(\ppm_encoder_1.counter24_0_I_1_c_RNOZ0 ));
    CascadeMux I__9767 (
            .O(N__42417),
            .I(N__42414));
    InMux I__9766 (
            .O(N__42414),
            .I(N__42411));
    LocalMux I__9765 (
            .O(N__42411),
            .I(N__42408));
    Odrv4 I__9764 (
            .O(N__42408),
            .I(\ppm_encoder_1.counter24_0_I_9_c_RNOZ0 ));
    InMux I__9763 (
            .O(N__42405),
            .I(N__42402));
    LocalMux I__9762 (
            .O(N__42402),
            .I(N__42399));
    Odrv4 I__9761 (
            .O(N__42399),
            .I(\ppm_encoder_1.init_pulses_RNI5ATG1Z0Z_15 ));
    InMux I__9760 (
            .O(N__42396),
            .I(N__42393));
    LocalMux I__9759 (
            .O(N__42393),
            .I(N__42390));
    Odrv12 I__9758 (
            .O(N__42390),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_15 ));
    InMux I__9757 (
            .O(N__42387),
            .I(N__42384));
    LocalMux I__9756 (
            .O(N__42384),
            .I(N__42381));
    Odrv12 I__9755 (
            .O(N__42381),
            .I(\ppm_encoder_1.un1_init_pulses_11_15 ));
    InMux I__9754 (
            .O(N__42378),
            .I(N__42375));
    LocalMux I__9753 (
            .O(N__42375),
            .I(N__42372));
    Odrv4 I__9752 (
            .O(N__42372),
            .I(\ppm_encoder_1.un1_init_pulses_10_15 ));
    InMux I__9751 (
            .O(N__42369),
            .I(N__42366));
    LocalMux I__9750 (
            .O(N__42366),
            .I(N__42363));
    Span4Mux_h I__9749 (
            .O(N__42363),
            .I(N__42358));
    InMux I__9748 (
            .O(N__42362),
            .I(N__42353));
    InMux I__9747 (
            .O(N__42361),
            .I(N__42353));
    Odrv4 I__9746 (
            .O(N__42358),
            .I(\ppm_encoder_1.init_pulsesZ0Z_15 ));
    LocalMux I__9745 (
            .O(N__42353),
            .I(\ppm_encoder_1.init_pulsesZ0Z_15 ));
    InMux I__9744 (
            .O(N__42348),
            .I(N__42343));
    InMux I__9743 (
            .O(N__42347),
            .I(N__42338));
    InMux I__9742 (
            .O(N__42346),
            .I(N__42338));
    LocalMux I__9741 (
            .O(N__42343),
            .I(N__42334));
    LocalMux I__9740 (
            .O(N__42338),
            .I(N__42331));
    InMux I__9739 (
            .O(N__42337),
            .I(N__42328));
    Span4Mux_v I__9738 (
            .O(N__42334),
            .I(N__42320));
    Span4Mux_h I__9737 (
            .O(N__42331),
            .I(N__42317));
    LocalMux I__9736 (
            .O(N__42328),
            .I(N__42314));
    InMux I__9735 (
            .O(N__42327),
            .I(N__42311));
    InMux I__9734 (
            .O(N__42326),
            .I(N__42302));
    InMux I__9733 (
            .O(N__42325),
            .I(N__42302));
    InMux I__9732 (
            .O(N__42324),
            .I(N__42302));
    InMux I__9731 (
            .O(N__42323),
            .I(N__42302));
    Odrv4 I__9730 (
            .O(N__42320),
            .I(\ppm_encoder_1.un1_init_pulses_0Z0Z_1 ));
    Odrv4 I__9729 (
            .O(N__42317),
            .I(\ppm_encoder_1.un1_init_pulses_0Z0Z_1 ));
    Odrv12 I__9728 (
            .O(N__42314),
            .I(\ppm_encoder_1.un1_init_pulses_0Z0Z_1 ));
    LocalMux I__9727 (
            .O(N__42311),
            .I(\ppm_encoder_1.un1_init_pulses_0Z0Z_1 ));
    LocalMux I__9726 (
            .O(N__42302),
            .I(\ppm_encoder_1.un1_init_pulses_0Z0Z_1 ));
    CascadeMux I__9725 (
            .O(N__42291),
            .I(N__42281));
    CascadeMux I__9724 (
            .O(N__42290),
            .I(N__42278));
    InMux I__9723 (
            .O(N__42289),
            .I(N__42267));
    InMux I__9722 (
            .O(N__42288),
            .I(N__42260));
    InMux I__9721 (
            .O(N__42287),
            .I(N__42260));
    InMux I__9720 (
            .O(N__42286),
            .I(N__42260));
    CascadeMux I__9719 (
            .O(N__42285),
            .I(N__42255));
    CascadeMux I__9718 (
            .O(N__42284),
            .I(N__42251));
    InMux I__9717 (
            .O(N__42281),
            .I(N__42238));
    InMux I__9716 (
            .O(N__42278),
            .I(N__42238));
    InMux I__9715 (
            .O(N__42277),
            .I(N__42238));
    InMux I__9714 (
            .O(N__42276),
            .I(N__42238));
    InMux I__9713 (
            .O(N__42275),
            .I(N__42235));
    InMux I__9712 (
            .O(N__42274),
            .I(N__42225));
    InMux I__9711 (
            .O(N__42273),
            .I(N__42222));
    InMux I__9710 (
            .O(N__42272),
            .I(N__42219));
    InMux I__9709 (
            .O(N__42271),
            .I(N__42214));
    InMux I__9708 (
            .O(N__42270),
            .I(N__42214));
    LocalMux I__9707 (
            .O(N__42267),
            .I(N__42209));
    LocalMux I__9706 (
            .O(N__42260),
            .I(N__42209));
    InMux I__9705 (
            .O(N__42259),
            .I(N__42204));
    InMux I__9704 (
            .O(N__42258),
            .I(N__42204));
    InMux I__9703 (
            .O(N__42255),
            .I(N__42195));
    InMux I__9702 (
            .O(N__42254),
            .I(N__42195));
    InMux I__9701 (
            .O(N__42251),
            .I(N__42195));
    InMux I__9700 (
            .O(N__42250),
            .I(N__42195));
    InMux I__9699 (
            .O(N__42249),
            .I(N__42188));
    InMux I__9698 (
            .O(N__42248),
            .I(N__42188));
    InMux I__9697 (
            .O(N__42247),
            .I(N__42188));
    LocalMux I__9696 (
            .O(N__42238),
            .I(N__42185));
    LocalMux I__9695 (
            .O(N__42235),
            .I(N__42182));
    InMux I__9694 (
            .O(N__42234),
            .I(N__42179));
    InMux I__9693 (
            .O(N__42233),
            .I(N__42176));
    CascadeMux I__9692 (
            .O(N__42232),
            .I(N__42173));
    CascadeMux I__9691 (
            .O(N__42231),
            .I(N__42168));
    CascadeMux I__9690 (
            .O(N__42230),
            .I(N__42159));
    InMux I__9689 (
            .O(N__42229),
            .I(N__42155));
    CascadeMux I__9688 (
            .O(N__42228),
            .I(N__42152));
    LocalMux I__9687 (
            .O(N__42225),
            .I(N__42148));
    LocalMux I__9686 (
            .O(N__42222),
            .I(N__42133));
    LocalMux I__9685 (
            .O(N__42219),
            .I(N__42133));
    LocalMux I__9684 (
            .O(N__42214),
            .I(N__42133));
    Span4Mux_v I__9683 (
            .O(N__42209),
            .I(N__42133));
    LocalMux I__9682 (
            .O(N__42204),
            .I(N__42133));
    LocalMux I__9681 (
            .O(N__42195),
            .I(N__42133));
    LocalMux I__9680 (
            .O(N__42188),
            .I(N__42133));
    Span4Mux_v I__9679 (
            .O(N__42185),
            .I(N__42130));
    Span4Mux_v I__9678 (
            .O(N__42182),
            .I(N__42127));
    LocalMux I__9677 (
            .O(N__42179),
            .I(N__42122));
    LocalMux I__9676 (
            .O(N__42176),
            .I(N__42122));
    InMux I__9675 (
            .O(N__42173),
            .I(N__42115));
    InMux I__9674 (
            .O(N__42172),
            .I(N__42115));
    InMux I__9673 (
            .O(N__42171),
            .I(N__42115));
    InMux I__9672 (
            .O(N__42168),
            .I(N__42111));
    InMux I__9671 (
            .O(N__42167),
            .I(N__42106));
    InMux I__9670 (
            .O(N__42166),
            .I(N__42106));
    InMux I__9669 (
            .O(N__42165),
            .I(N__42097));
    InMux I__9668 (
            .O(N__42164),
            .I(N__42097));
    InMux I__9667 (
            .O(N__42163),
            .I(N__42097));
    InMux I__9666 (
            .O(N__42162),
            .I(N__42097));
    InMux I__9665 (
            .O(N__42159),
            .I(N__42092));
    InMux I__9664 (
            .O(N__42158),
            .I(N__42092));
    LocalMux I__9663 (
            .O(N__42155),
            .I(N__42089));
    InMux I__9662 (
            .O(N__42152),
            .I(N__42084));
    InMux I__9661 (
            .O(N__42151),
            .I(N__42084));
    Span4Mux_h I__9660 (
            .O(N__42148),
            .I(N__42077));
    Span4Mux_v I__9659 (
            .O(N__42133),
            .I(N__42077));
    Span4Mux_v I__9658 (
            .O(N__42130),
            .I(N__42077));
    Span4Mux_h I__9657 (
            .O(N__42127),
            .I(N__42070));
    Span4Mux_v I__9656 (
            .O(N__42122),
            .I(N__42070));
    LocalMux I__9655 (
            .O(N__42115),
            .I(N__42070));
    InMux I__9654 (
            .O(N__42114),
            .I(N__42067));
    LocalMux I__9653 (
            .O(N__42111),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_d_12 ));
    LocalMux I__9652 (
            .O(N__42106),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_d_12 ));
    LocalMux I__9651 (
            .O(N__42097),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_d_12 ));
    LocalMux I__9650 (
            .O(N__42092),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_d_12 ));
    Odrv4 I__9649 (
            .O(N__42089),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_d_12 ));
    LocalMux I__9648 (
            .O(N__42084),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_d_12 ));
    Odrv4 I__9647 (
            .O(N__42077),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_d_12 ));
    Odrv4 I__9646 (
            .O(N__42070),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_d_12 ));
    LocalMux I__9645 (
            .O(N__42067),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_d_12 ));
    CascadeMux I__9644 (
            .O(N__42048),
            .I(N__42044));
    CascadeMux I__9643 (
            .O(N__42047),
            .I(N__42031));
    InMux I__9642 (
            .O(N__42044),
            .I(N__42024));
    InMux I__9641 (
            .O(N__42043),
            .I(N__42024));
    InMux I__9640 (
            .O(N__42042),
            .I(N__42024));
    CascadeMux I__9639 (
            .O(N__42041),
            .I(N__42015));
    CascadeMux I__9638 (
            .O(N__42040),
            .I(N__42012));
    CascadeMux I__9637 (
            .O(N__42039),
            .I(N__42004));
    InMux I__9636 (
            .O(N__42038),
            .I(N__41999));
    CascadeMux I__9635 (
            .O(N__42037),
            .I(N__41988));
    CascadeMux I__9634 (
            .O(N__42036),
            .I(N__41985));
    InMux I__9633 (
            .O(N__42035),
            .I(N__41979));
    InMux I__9632 (
            .O(N__42034),
            .I(N__41979));
    InMux I__9631 (
            .O(N__42031),
            .I(N__41972));
    LocalMux I__9630 (
            .O(N__42024),
            .I(N__41969));
    InMux I__9629 (
            .O(N__42023),
            .I(N__41964));
    InMux I__9628 (
            .O(N__42022),
            .I(N__41964));
    InMux I__9627 (
            .O(N__42021),
            .I(N__41955));
    InMux I__9626 (
            .O(N__42020),
            .I(N__41955));
    InMux I__9625 (
            .O(N__42019),
            .I(N__41955));
    InMux I__9624 (
            .O(N__42018),
            .I(N__41955));
    InMux I__9623 (
            .O(N__42015),
            .I(N__41948));
    InMux I__9622 (
            .O(N__42012),
            .I(N__41948));
    InMux I__9621 (
            .O(N__42011),
            .I(N__41948));
    InMux I__9620 (
            .O(N__42010),
            .I(N__41933));
    InMux I__9619 (
            .O(N__42009),
            .I(N__41930));
    InMux I__9618 (
            .O(N__42008),
            .I(N__41925));
    InMux I__9617 (
            .O(N__42007),
            .I(N__41925));
    InMux I__9616 (
            .O(N__42004),
            .I(N__41916));
    InMux I__9615 (
            .O(N__42003),
            .I(N__41916));
    InMux I__9614 (
            .O(N__42002),
            .I(N__41913));
    LocalMux I__9613 (
            .O(N__41999),
            .I(N__41910));
    InMux I__9612 (
            .O(N__41998),
            .I(N__41905));
    InMux I__9611 (
            .O(N__41997),
            .I(N__41905));
    InMux I__9610 (
            .O(N__41996),
            .I(N__41900));
    InMux I__9609 (
            .O(N__41995),
            .I(N__41900));
    InMux I__9608 (
            .O(N__41994),
            .I(N__41893));
    InMux I__9607 (
            .O(N__41993),
            .I(N__41893));
    InMux I__9606 (
            .O(N__41992),
            .I(N__41893));
    InMux I__9605 (
            .O(N__41991),
            .I(N__41883));
    InMux I__9604 (
            .O(N__41988),
            .I(N__41883));
    InMux I__9603 (
            .O(N__41985),
            .I(N__41883));
    InMux I__9602 (
            .O(N__41984),
            .I(N__41883));
    LocalMux I__9601 (
            .O(N__41979),
            .I(N__41880));
    InMux I__9600 (
            .O(N__41978),
            .I(N__41871));
    InMux I__9599 (
            .O(N__41977),
            .I(N__41871));
    InMux I__9598 (
            .O(N__41976),
            .I(N__41871));
    InMux I__9597 (
            .O(N__41975),
            .I(N__41871));
    LocalMux I__9596 (
            .O(N__41972),
            .I(N__41864));
    Span4Mux_v I__9595 (
            .O(N__41969),
            .I(N__41864));
    LocalMux I__9594 (
            .O(N__41964),
            .I(N__41864));
    LocalMux I__9593 (
            .O(N__41955),
            .I(N__41859));
    LocalMux I__9592 (
            .O(N__41948),
            .I(N__41859));
    InMux I__9591 (
            .O(N__41947),
            .I(N__41848));
    InMux I__9590 (
            .O(N__41946),
            .I(N__41848));
    InMux I__9589 (
            .O(N__41945),
            .I(N__41848));
    InMux I__9588 (
            .O(N__41944),
            .I(N__41848));
    InMux I__9587 (
            .O(N__41943),
            .I(N__41848));
    InMux I__9586 (
            .O(N__41942),
            .I(N__41841));
    InMux I__9585 (
            .O(N__41941),
            .I(N__41841));
    InMux I__9584 (
            .O(N__41940),
            .I(N__41841));
    InMux I__9583 (
            .O(N__41939),
            .I(N__41837));
    InMux I__9582 (
            .O(N__41938),
            .I(N__41830));
    InMux I__9581 (
            .O(N__41937),
            .I(N__41830));
    InMux I__9580 (
            .O(N__41936),
            .I(N__41830));
    LocalMux I__9579 (
            .O(N__41933),
            .I(N__41827));
    LocalMux I__9578 (
            .O(N__41930),
            .I(N__41822));
    LocalMux I__9577 (
            .O(N__41925),
            .I(N__41822));
    InMux I__9576 (
            .O(N__41924),
            .I(N__41817));
    InMux I__9575 (
            .O(N__41923),
            .I(N__41817));
    InMux I__9574 (
            .O(N__41922),
            .I(N__41811));
    InMux I__9573 (
            .O(N__41921),
            .I(N__41808));
    LocalMux I__9572 (
            .O(N__41916),
            .I(N__41795));
    LocalMux I__9571 (
            .O(N__41913),
            .I(N__41795));
    Span4Mux_v I__9570 (
            .O(N__41910),
            .I(N__41795));
    LocalMux I__9569 (
            .O(N__41905),
            .I(N__41795));
    LocalMux I__9568 (
            .O(N__41900),
            .I(N__41795));
    LocalMux I__9567 (
            .O(N__41893),
            .I(N__41795));
    InMux I__9566 (
            .O(N__41892),
            .I(N__41792));
    LocalMux I__9565 (
            .O(N__41883),
            .I(N__41785));
    Span4Mux_v I__9564 (
            .O(N__41880),
            .I(N__41785));
    LocalMux I__9563 (
            .O(N__41871),
            .I(N__41785));
    Span4Mux_v I__9562 (
            .O(N__41864),
            .I(N__41778));
    Span4Mux_v I__9561 (
            .O(N__41859),
            .I(N__41778));
    LocalMux I__9560 (
            .O(N__41848),
            .I(N__41778));
    LocalMux I__9559 (
            .O(N__41841),
            .I(N__41767));
    InMux I__9558 (
            .O(N__41840),
            .I(N__41764));
    LocalMux I__9557 (
            .O(N__41837),
            .I(N__41759));
    LocalMux I__9556 (
            .O(N__41830),
            .I(N__41759));
    Span4Mux_h I__9555 (
            .O(N__41827),
            .I(N__41752));
    Span4Mux_v I__9554 (
            .O(N__41822),
            .I(N__41752));
    LocalMux I__9553 (
            .O(N__41817),
            .I(N__41752));
    InMux I__9552 (
            .O(N__41816),
            .I(N__41747));
    InMux I__9551 (
            .O(N__41815),
            .I(N__41747));
    InMux I__9550 (
            .O(N__41814),
            .I(N__41744));
    LocalMux I__9549 (
            .O(N__41811),
            .I(N__41741));
    LocalMux I__9548 (
            .O(N__41808),
            .I(N__41736));
    Span4Mux_v I__9547 (
            .O(N__41795),
            .I(N__41736));
    LocalMux I__9546 (
            .O(N__41792),
            .I(N__41729));
    Span4Mux_h I__9545 (
            .O(N__41785),
            .I(N__41729));
    Span4Mux_h I__9544 (
            .O(N__41778),
            .I(N__41729));
    InMux I__9543 (
            .O(N__41777),
            .I(N__41726));
    InMux I__9542 (
            .O(N__41776),
            .I(N__41723));
    InMux I__9541 (
            .O(N__41775),
            .I(N__41710));
    InMux I__9540 (
            .O(N__41774),
            .I(N__41710));
    InMux I__9539 (
            .O(N__41773),
            .I(N__41710));
    InMux I__9538 (
            .O(N__41772),
            .I(N__41710));
    InMux I__9537 (
            .O(N__41771),
            .I(N__41710));
    InMux I__9536 (
            .O(N__41770),
            .I(N__41710));
    Span4Mux_h I__9535 (
            .O(N__41767),
            .I(N__41701));
    LocalMux I__9534 (
            .O(N__41764),
            .I(N__41701));
    Span4Mux_h I__9533 (
            .O(N__41759),
            .I(N__41701));
    Span4Mux_v I__9532 (
            .O(N__41752),
            .I(N__41701));
    LocalMux I__9531 (
            .O(N__41747),
            .I(N__41698));
    LocalMux I__9530 (
            .O(N__41744),
            .I(N__41691));
    Span4Mux_v I__9529 (
            .O(N__41741),
            .I(N__41691));
    Span4Mux_v I__9528 (
            .O(N__41736),
            .I(N__41691));
    Span4Mux_v I__9527 (
            .O(N__41729),
            .I(N__41688));
    LocalMux I__9526 (
            .O(N__41726),
            .I(\ppm_encoder_1.PPM_STATE_59_d ));
    LocalMux I__9525 (
            .O(N__41723),
            .I(\ppm_encoder_1.PPM_STATE_59_d ));
    LocalMux I__9524 (
            .O(N__41710),
            .I(\ppm_encoder_1.PPM_STATE_59_d ));
    Odrv4 I__9523 (
            .O(N__41701),
            .I(\ppm_encoder_1.PPM_STATE_59_d ));
    Odrv12 I__9522 (
            .O(N__41698),
            .I(\ppm_encoder_1.PPM_STATE_59_d ));
    Odrv4 I__9521 (
            .O(N__41691),
            .I(\ppm_encoder_1.PPM_STATE_59_d ));
    Odrv4 I__9520 (
            .O(N__41688),
            .I(\ppm_encoder_1.PPM_STATE_59_d ));
    InMux I__9519 (
            .O(N__41673),
            .I(N__41670));
    LocalMux I__9518 (
            .O(N__41670),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_18 ));
    InMux I__9517 (
            .O(N__41667),
            .I(N__41664));
    LocalMux I__9516 (
            .O(N__41664),
            .I(N__41661));
    Odrv12 I__9515 (
            .O(N__41661),
            .I(\ppm_encoder_1.un1_init_pulses_11_18 ));
    InMux I__9514 (
            .O(N__41658),
            .I(N__41655));
    LocalMux I__9513 (
            .O(N__41655),
            .I(\ppm_encoder_1.un1_init_pulses_10_18 ));
    CascadeMux I__9512 (
            .O(N__41652),
            .I(N__41648));
    InMux I__9511 (
            .O(N__41651),
            .I(N__41645));
    InMux I__9510 (
            .O(N__41648),
            .I(N__41642));
    LocalMux I__9509 (
            .O(N__41645),
            .I(N__41638));
    LocalMux I__9508 (
            .O(N__41642),
            .I(N__41635));
    CascadeMux I__9507 (
            .O(N__41641),
            .I(N__41632));
    Span4Mux_v I__9506 (
            .O(N__41638),
            .I(N__41627));
    Span4Mux_h I__9505 (
            .O(N__41635),
            .I(N__41627));
    InMux I__9504 (
            .O(N__41632),
            .I(N__41624));
    Odrv4 I__9503 (
            .O(N__41627),
            .I(\ppm_encoder_1.init_pulsesZ0Z_18 ));
    LocalMux I__9502 (
            .O(N__41624),
            .I(\ppm_encoder_1.init_pulsesZ0Z_18 ));
    CascadeMux I__9501 (
            .O(N__41619),
            .I(N__41603));
    CascadeMux I__9500 (
            .O(N__41618),
            .I(N__41596));
    InMux I__9499 (
            .O(N__41617),
            .I(N__41590));
    InMux I__9498 (
            .O(N__41616),
            .I(N__41590));
    InMux I__9497 (
            .O(N__41615),
            .I(N__41587));
    InMux I__9496 (
            .O(N__41614),
            .I(N__41584));
    InMux I__9495 (
            .O(N__41613),
            .I(N__41579));
    InMux I__9494 (
            .O(N__41612),
            .I(N__41579));
    InMux I__9493 (
            .O(N__41611),
            .I(N__41576));
    InMux I__9492 (
            .O(N__41610),
            .I(N__41573));
    InMux I__9491 (
            .O(N__41609),
            .I(N__41566));
    InMux I__9490 (
            .O(N__41608),
            .I(N__41566));
    InMux I__9489 (
            .O(N__41607),
            .I(N__41566));
    InMux I__9488 (
            .O(N__41606),
            .I(N__41557));
    InMux I__9487 (
            .O(N__41603),
            .I(N__41557));
    InMux I__9486 (
            .O(N__41602),
            .I(N__41557));
    InMux I__9485 (
            .O(N__41601),
            .I(N__41557));
    InMux I__9484 (
            .O(N__41600),
            .I(N__41552));
    InMux I__9483 (
            .O(N__41599),
            .I(N__41552));
    InMux I__9482 (
            .O(N__41596),
            .I(N__41547));
    InMux I__9481 (
            .O(N__41595),
            .I(N__41547));
    LocalMux I__9480 (
            .O(N__41590),
            .I(N__41542));
    LocalMux I__9479 (
            .O(N__41587),
            .I(N__41542));
    LocalMux I__9478 (
            .O(N__41584),
            .I(N__41537));
    LocalMux I__9477 (
            .O(N__41579),
            .I(N__41537));
    LocalMux I__9476 (
            .O(N__41576),
            .I(N__41534));
    LocalMux I__9475 (
            .O(N__41573),
            .I(N__41529));
    LocalMux I__9474 (
            .O(N__41566),
            .I(N__41529));
    LocalMux I__9473 (
            .O(N__41557),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_1 ));
    LocalMux I__9472 (
            .O(N__41552),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_1 ));
    LocalMux I__9471 (
            .O(N__41547),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_1 ));
    Odrv4 I__9470 (
            .O(N__41542),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_1 ));
    Odrv4 I__9469 (
            .O(N__41537),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_1 ));
    Odrv4 I__9468 (
            .O(N__41534),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_1 ));
    Odrv12 I__9467 (
            .O(N__41529),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_1 ));
    InMux I__9466 (
            .O(N__41514),
            .I(N__41511));
    LocalMux I__9465 (
            .O(N__41511),
            .I(N__41508));
    Span4Mux_v I__9464 (
            .O(N__41508),
            .I(N__41505));
    Odrv4 I__9463 (
            .O(N__41505),
            .I(\ppm_encoder_1.un1_init_pulses_11_13 ));
    CascadeMux I__9462 (
            .O(N__41502),
            .I(N__41493));
    CascadeMux I__9461 (
            .O(N__41501),
            .I(N__41490));
    CascadeMux I__9460 (
            .O(N__41500),
            .I(N__41487));
    CascadeMux I__9459 (
            .O(N__41499),
            .I(N__41484));
    CascadeMux I__9458 (
            .O(N__41498),
            .I(N__41481));
    CascadeMux I__9457 (
            .O(N__41497),
            .I(N__41478));
    CascadeMux I__9456 (
            .O(N__41496),
            .I(N__41475));
    InMux I__9455 (
            .O(N__41493),
            .I(N__41466));
    InMux I__9454 (
            .O(N__41490),
            .I(N__41466));
    InMux I__9453 (
            .O(N__41487),
            .I(N__41466));
    InMux I__9452 (
            .O(N__41484),
            .I(N__41463));
    InMux I__9451 (
            .O(N__41481),
            .I(N__41458));
    InMux I__9450 (
            .O(N__41478),
            .I(N__41458));
    InMux I__9449 (
            .O(N__41475),
            .I(N__41455));
    CascadeMux I__9448 (
            .O(N__41474),
            .I(N__41452));
    CascadeMux I__9447 (
            .O(N__41473),
            .I(N__41449));
    LocalMux I__9446 (
            .O(N__41466),
            .I(N__41435));
    LocalMux I__9445 (
            .O(N__41463),
            .I(N__41435));
    LocalMux I__9444 (
            .O(N__41458),
            .I(N__41435));
    LocalMux I__9443 (
            .O(N__41455),
            .I(N__41435));
    InMux I__9442 (
            .O(N__41452),
            .I(N__41430));
    InMux I__9441 (
            .O(N__41449),
            .I(N__41430));
    CascadeMux I__9440 (
            .O(N__41448),
            .I(N__41427));
    CascadeMux I__9439 (
            .O(N__41447),
            .I(N__41424));
    CascadeMux I__9438 (
            .O(N__41446),
            .I(N__41420));
    InMux I__9437 (
            .O(N__41445),
            .I(N__41416));
    CascadeMux I__9436 (
            .O(N__41444),
            .I(N__41413));
    Span4Mux_v I__9435 (
            .O(N__41435),
            .I(N__41406));
    LocalMux I__9434 (
            .O(N__41430),
            .I(N__41406));
    InMux I__9433 (
            .O(N__41427),
            .I(N__41403));
    InMux I__9432 (
            .O(N__41424),
            .I(N__41400));
    InMux I__9431 (
            .O(N__41423),
            .I(N__41393));
    InMux I__9430 (
            .O(N__41420),
            .I(N__41393));
    InMux I__9429 (
            .O(N__41419),
            .I(N__41393));
    LocalMux I__9428 (
            .O(N__41416),
            .I(N__41390));
    InMux I__9427 (
            .O(N__41413),
            .I(N__41387));
    CascadeMux I__9426 (
            .O(N__41412),
            .I(N__41384));
    CascadeMux I__9425 (
            .O(N__41411),
            .I(N__41381));
    Span4Mux_v I__9424 (
            .O(N__41406),
            .I(N__41377));
    LocalMux I__9423 (
            .O(N__41403),
            .I(N__41370));
    LocalMux I__9422 (
            .O(N__41400),
            .I(N__41370));
    LocalMux I__9421 (
            .O(N__41393),
            .I(N__41370));
    Span4Mux_h I__9420 (
            .O(N__41390),
            .I(N__41365));
    LocalMux I__9419 (
            .O(N__41387),
            .I(N__41365));
    InMux I__9418 (
            .O(N__41384),
            .I(N__41360));
    InMux I__9417 (
            .O(N__41381),
            .I(N__41360));
    InMux I__9416 (
            .O(N__41380),
            .I(N__41357));
    Odrv4 I__9415 (
            .O(N__41377),
            .I(\ppm_encoder_1.un1_init_pulses_4_sqmuxa_0 ));
    Odrv4 I__9414 (
            .O(N__41370),
            .I(\ppm_encoder_1.un1_init_pulses_4_sqmuxa_0 ));
    Odrv4 I__9413 (
            .O(N__41365),
            .I(\ppm_encoder_1.un1_init_pulses_4_sqmuxa_0 ));
    LocalMux I__9412 (
            .O(N__41360),
            .I(\ppm_encoder_1.un1_init_pulses_4_sqmuxa_0 ));
    LocalMux I__9411 (
            .O(N__41357),
            .I(\ppm_encoder_1.un1_init_pulses_4_sqmuxa_0 ));
    InMux I__9410 (
            .O(N__41346),
            .I(N__41343));
    LocalMux I__9409 (
            .O(N__41343),
            .I(N__41340));
    Odrv4 I__9408 (
            .O(N__41340),
            .I(\ppm_encoder_1.un1_init_pulses_10_13 ));
    InMux I__9407 (
            .O(N__41337),
            .I(N__41333));
    CascadeMux I__9406 (
            .O(N__41336),
            .I(N__41329));
    LocalMux I__9405 (
            .O(N__41333),
            .I(N__41326));
    InMux I__9404 (
            .O(N__41332),
            .I(N__41323));
    InMux I__9403 (
            .O(N__41329),
            .I(N__41320));
    Span4Mux_v I__9402 (
            .O(N__41326),
            .I(N__41317));
    LocalMux I__9401 (
            .O(N__41323),
            .I(N__41314));
    LocalMux I__9400 (
            .O(N__41320),
            .I(\ppm_encoder_1.init_pulsesZ0Z_13 ));
    Odrv4 I__9399 (
            .O(N__41317),
            .I(\ppm_encoder_1.init_pulsesZ0Z_13 ));
    Odrv4 I__9398 (
            .O(N__41314),
            .I(\ppm_encoder_1.init_pulsesZ0Z_13 ));
    InMux I__9397 (
            .O(N__41307),
            .I(N__41304));
    LocalMux I__9396 (
            .O(N__41304),
            .I(N__41301));
    Odrv4 I__9395 (
            .O(N__41301),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_14 ));
    InMux I__9394 (
            .O(N__41298),
            .I(N__41295));
    LocalMux I__9393 (
            .O(N__41295),
            .I(N__41292));
    Odrv4 I__9392 (
            .O(N__41292),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_14 ));
    InMux I__9391 (
            .O(N__41289),
            .I(N__41286));
    LocalMux I__9390 (
            .O(N__41286),
            .I(N__41283));
    Odrv4 I__9389 (
            .O(N__41283),
            .I(\ppm_encoder_1.pulses2countZ0Z_14 ));
    InMux I__9388 (
            .O(N__41280),
            .I(N__41277));
    LocalMux I__9387 (
            .O(N__41277),
            .I(N__41274));
    Span4Mux_h I__9386 (
            .O(N__41274),
            .I(N__41271));
    Odrv4 I__9385 (
            .O(N__41271),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_10 ));
    InMux I__9384 (
            .O(N__41268),
            .I(N__41265));
    LocalMux I__9383 (
            .O(N__41265),
            .I(N__41262));
    Span4Mux_h I__9382 (
            .O(N__41262),
            .I(N__41259));
    Odrv4 I__9381 (
            .O(N__41259),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_10 ));
    InMux I__9380 (
            .O(N__41256),
            .I(N__41253));
    LocalMux I__9379 (
            .O(N__41253),
            .I(N__41250));
    Odrv4 I__9378 (
            .O(N__41250),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_17 ));
    InMux I__9377 (
            .O(N__41247),
            .I(N__41243));
    InMux I__9376 (
            .O(N__41246),
            .I(N__41239));
    LocalMux I__9375 (
            .O(N__41243),
            .I(N__41236));
    InMux I__9374 (
            .O(N__41242),
            .I(N__41233));
    LocalMux I__9373 (
            .O(N__41239),
            .I(N__41230));
    Span4Mux_v I__9372 (
            .O(N__41236),
            .I(N__41227));
    LocalMux I__9371 (
            .O(N__41233),
            .I(N__41222));
    Span4Mux_v I__9370 (
            .O(N__41230),
            .I(N__41222));
    Odrv4 I__9369 (
            .O(N__41227),
            .I(\ppm_encoder_1.init_pulsesZ0Z_10 ));
    Odrv4 I__9368 (
            .O(N__41222),
            .I(\ppm_encoder_1.init_pulsesZ0Z_10 ));
    InMux I__9367 (
            .O(N__41217),
            .I(N__41214));
    LocalMux I__9366 (
            .O(N__41214),
            .I(N__41211));
    Span4Mux_v I__9365 (
            .O(N__41211),
            .I(N__41208));
    Odrv4 I__9364 (
            .O(N__41208),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_10 ));
    InMux I__9363 (
            .O(N__41205),
            .I(N__41202));
    LocalMux I__9362 (
            .O(N__41202),
            .I(N__41199));
    Odrv12 I__9361 (
            .O(N__41199),
            .I(\ppm_encoder_1.un1_init_pulses_11_14 ));
    InMux I__9360 (
            .O(N__41196),
            .I(N__41193));
    LocalMux I__9359 (
            .O(N__41193),
            .I(\ppm_encoder_1.un1_init_pulses_10_14 ));
    InMux I__9358 (
            .O(N__41190),
            .I(N__41187));
    LocalMux I__9357 (
            .O(N__41187),
            .I(N__41184));
    Span4Mux_v I__9356 (
            .O(N__41184),
            .I(N__41180));
    InMux I__9355 (
            .O(N__41183),
            .I(N__41177));
    Odrv4 I__9354 (
            .O(N__41180),
            .I(\ppm_encoder_1.un1_init_pulses_0_14 ));
    LocalMux I__9353 (
            .O(N__41177),
            .I(\ppm_encoder_1.un1_init_pulses_0_14 ));
    InMux I__9352 (
            .O(N__41172),
            .I(N__41169));
    LocalMux I__9351 (
            .O(N__41169),
            .I(N__41166));
    Span4Mux_v I__9350 (
            .O(N__41166),
            .I(N__41163));
    Odrv4 I__9349 (
            .O(N__41163),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_14 ));
    InMux I__9348 (
            .O(N__41160),
            .I(N__41151));
    InMux I__9347 (
            .O(N__41159),
            .I(N__41151));
    InMux I__9346 (
            .O(N__41158),
            .I(N__41151));
    LocalMux I__9345 (
            .O(N__41151),
            .I(\ppm_encoder_1.init_pulsesZ0Z_14 ));
    InMux I__9344 (
            .O(N__41148),
            .I(N__41142));
    InMux I__9343 (
            .O(N__41147),
            .I(N__41138));
    InMux I__9342 (
            .O(N__41146),
            .I(N__41133));
    InMux I__9341 (
            .O(N__41145),
            .I(N__41133));
    LocalMux I__9340 (
            .O(N__41142),
            .I(N__41129));
    InMux I__9339 (
            .O(N__41141),
            .I(N__41125));
    LocalMux I__9338 (
            .O(N__41138),
            .I(N__41118));
    LocalMux I__9337 (
            .O(N__41133),
            .I(N__41115));
    InMux I__9336 (
            .O(N__41132),
            .I(N__41112));
    Span4Mux_v I__9335 (
            .O(N__41129),
            .I(N__41109));
    InMux I__9334 (
            .O(N__41128),
            .I(N__41106));
    LocalMux I__9333 (
            .O(N__41125),
            .I(N__41103));
    InMux I__9332 (
            .O(N__41124),
            .I(N__41098));
    InMux I__9331 (
            .O(N__41123),
            .I(N__41098));
    InMux I__9330 (
            .O(N__41122),
            .I(N__41095));
    CascadeMux I__9329 (
            .O(N__41121),
            .I(N__41091));
    Span4Mux_v I__9328 (
            .O(N__41118),
            .I(N__41084));
    Span4Mux_h I__9327 (
            .O(N__41115),
            .I(N__41084));
    LocalMux I__9326 (
            .O(N__41112),
            .I(N__41084));
    Span4Mux_h I__9325 (
            .O(N__41109),
            .I(N__41079));
    LocalMux I__9324 (
            .O(N__41106),
            .I(N__41079));
    Span4Mux_v I__9323 (
            .O(N__41103),
            .I(N__41074));
    LocalMux I__9322 (
            .O(N__41098),
            .I(N__41074));
    LocalMux I__9321 (
            .O(N__41095),
            .I(N__41071));
    InMux I__9320 (
            .O(N__41094),
            .I(N__41068));
    InMux I__9319 (
            .O(N__41091),
            .I(N__41065));
    Span4Mux_v I__9318 (
            .O(N__41084),
            .I(N__41059));
    Span4Mux_v I__9317 (
            .O(N__41079),
            .I(N__41054));
    Span4Mux_h I__9316 (
            .O(N__41074),
            .I(N__41054));
    Span4Mux_h I__9315 (
            .O(N__41071),
            .I(N__41051));
    LocalMux I__9314 (
            .O(N__41068),
            .I(N__41046));
    LocalMux I__9313 (
            .O(N__41065),
            .I(N__41046));
    InMux I__9312 (
            .O(N__41064),
            .I(N__41041));
    InMux I__9311 (
            .O(N__41063),
            .I(N__41041));
    InMux I__9310 (
            .O(N__41062),
            .I(N__41038));
    Odrv4 I__9309 (
            .O(N__41059),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_7 ));
    Odrv4 I__9308 (
            .O(N__41054),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_7 ));
    Odrv4 I__9307 (
            .O(N__41051),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_7 ));
    Odrv12 I__9306 (
            .O(N__41046),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_7 ));
    LocalMux I__9305 (
            .O(N__41041),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_7 ));
    LocalMux I__9304 (
            .O(N__41038),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_7 ));
    CascadeMux I__9303 (
            .O(N__41025),
            .I(N__41022));
    InMux I__9302 (
            .O(N__41022),
            .I(N__41018));
    InMux I__9301 (
            .O(N__41021),
            .I(N__41015));
    LocalMux I__9300 (
            .O(N__41018),
            .I(N__41012));
    LocalMux I__9299 (
            .O(N__41015),
            .I(N__41009));
    Span4Mux_h I__9298 (
            .O(N__41012),
            .I(N__41006));
    Span4Mux_v I__9297 (
            .O(N__41009),
            .I(N__41003));
    Span4Mux_h I__9296 (
            .O(N__41006),
            .I(N__41000));
    Span4Mux_v I__9295 (
            .O(N__41003),
            .I(N__40997));
    Odrv4 I__9294 (
            .O(N__41000),
            .I(\ppm_encoder_1.rudderZ0Z_14 ));
    Odrv4 I__9293 (
            .O(N__40997),
            .I(\ppm_encoder_1.rudderZ0Z_14 ));
    CascadeMux I__9292 (
            .O(N__40992),
            .I(N__40985));
    CascadeMux I__9291 (
            .O(N__40991),
            .I(N__40979));
    InMux I__9290 (
            .O(N__40990),
            .I(N__40974));
    InMux I__9289 (
            .O(N__40989),
            .I(N__40971));
    InMux I__9288 (
            .O(N__40988),
            .I(N__40968));
    InMux I__9287 (
            .O(N__40985),
            .I(N__40965));
    CascadeMux I__9286 (
            .O(N__40984),
            .I(N__40962));
    CascadeMux I__9285 (
            .O(N__40983),
            .I(N__40959));
    InMux I__9284 (
            .O(N__40982),
            .I(N__40955));
    InMux I__9283 (
            .O(N__40979),
            .I(N__40952));
    InMux I__9282 (
            .O(N__40978),
            .I(N__40949));
    CascadeMux I__9281 (
            .O(N__40977),
            .I(N__40945));
    LocalMux I__9280 (
            .O(N__40974),
            .I(N__40936));
    LocalMux I__9279 (
            .O(N__40971),
            .I(N__40936));
    LocalMux I__9278 (
            .O(N__40968),
            .I(N__40936));
    LocalMux I__9277 (
            .O(N__40965),
            .I(N__40936));
    InMux I__9276 (
            .O(N__40962),
            .I(N__40931));
    InMux I__9275 (
            .O(N__40959),
            .I(N__40931));
    InMux I__9274 (
            .O(N__40958),
            .I(N__40923));
    LocalMux I__9273 (
            .O(N__40955),
            .I(N__40918));
    LocalMux I__9272 (
            .O(N__40952),
            .I(N__40918));
    LocalMux I__9271 (
            .O(N__40949),
            .I(N__40915));
    InMux I__9270 (
            .O(N__40948),
            .I(N__40910));
    InMux I__9269 (
            .O(N__40945),
            .I(N__40910));
    Span4Mux_v I__9268 (
            .O(N__40936),
            .I(N__40904));
    LocalMux I__9267 (
            .O(N__40931),
            .I(N__40904));
    CascadeMux I__9266 (
            .O(N__40930),
            .I(N__40901));
    CascadeMux I__9265 (
            .O(N__40929),
            .I(N__40898));
    InMux I__9264 (
            .O(N__40928),
            .I(N__40895));
    InMux I__9263 (
            .O(N__40927),
            .I(N__40892));
    CascadeMux I__9262 (
            .O(N__40926),
            .I(N__40889));
    LocalMux I__9261 (
            .O(N__40923),
            .I(N__40879));
    Span4Mux_v I__9260 (
            .O(N__40918),
            .I(N__40879));
    Span4Mux_h I__9259 (
            .O(N__40915),
            .I(N__40879));
    LocalMux I__9258 (
            .O(N__40910),
            .I(N__40879));
    InMux I__9257 (
            .O(N__40909),
            .I(N__40876));
    Span4Mux_v I__9256 (
            .O(N__40904),
            .I(N__40873));
    InMux I__9255 (
            .O(N__40901),
            .I(N__40870));
    InMux I__9254 (
            .O(N__40898),
            .I(N__40867));
    LocalMux I__9253 (
            .O(N__40895),
            .I(N__40864));
    LocalMux I__9252 (
            .O(N__40892),
            .I(N__40861));
    InMux I__9251 (
            .O(N__40889),
            .I(N__40858));
    InMux I__9250 (
            .O(N__40888),
            .I(N__40855));
    Span4Mux_v I__9249 (
            .O(N__40879),
            .I(N__40852));
    LocalMux I__9248 (
            .O(N__40876),
            .I(N__40849));
    Sp12to4 I__9247 (
            .O(N__40873),
            .I(N__40840));
    LocalMux I__9246 (
            .O(N__40870),
            .I(N__40840));
    LocalMux I__9245 (
            .O(N__40867),
            .I(N__40840));
    Span12Mux_v I__9244 (
            .O(N__40864),
            .I(N__40840));
    Span12Mux_v I__9243 (
            .O(N__40861),
            .I(N__40837));
    LocalMux I__9242 (
            .O(N__40858),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ));
    LocalMux I__9241 (
            .O(N__40855),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ));
    Odrv4 I__9240 (
            .O(N__40852),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ));
    Odrv4 I__9239 (
            .O(N__40849),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ));
    Odrv12 I__9238 (
            .O(N__40840),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ));
    Odrv12 I__9237 (
            .O(N__40837),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ));
    InMux I__9236 (
            .O(N__40824),
            .I(N__40821));
    LocalMux I__9235 (
            .O(N__40821),
            .I(N__40818));
    Odrv12 I__9234 (
            .O(N__40818),
            .I(\ppm_encoder_1.un1_init_pulses_11_16 ));
    InMux I__9233 (
            .O(N__40815),
            .I(N__40812));
    LocalMux I__9232 (
            .O(N__40812),
            .I(\ppm_encoder_1.un1_init_pulses_10_16 ));
    InMux I__9231 (
            .O(N__40809),
            .I(N__40806));
    LocalMux I__9230 (
            .O(N__40806),
            .I(N__40803));
    Span4Mux_h I__9229 (
            .O(N__40803),
            .I(N__40800));
    Span4Mux_h I__9228 (
            .O(N__40800),
            .I(N__40795));
    InMux I__9227 (
            .O(N__40799),
            .I(N__40792));
    InMux I__9226 (
            .O(N__40798),
            .I(N__40789));
    Odrv4 I__9225 (
            .O(N__40795),
            .I(\ppm_encoder_1.init_pulsesZ0Z_16 ));
    LocalMux I__9224 (
            .O(N__40792),
            .I(\ppm_encoder_1.init_pulsesZ0Z_16 ));
    LocalMux I__9223 (
            .O(N__40789),
            .I(\ppm_encoder_1.init_pulsesZ0Z_16 ));
    CascadeMux I__9222 (
            .O(N__40782),
            .I(N__40779));
    InMux I__9221 (
            .O(N__40779),
            .I(N__40776));
    LocalMux I__9220 (
            .O(N__40776),
            .I(N__40773));
    Odrv12 I__9219 (
            .O(N__40773),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_16 ));
    InMux I__9218 (
            .O(N__40770),
            .I(N__40767));
    LocalMux I__9217 (
            .O(N__40767),
            .I(N__40764));
    Odrv12 I__9216 (
            .O(N__40764),
            .I(\ppm_encoder_1.un1_init_pulses_11_17 ));
    InMux I__9215 (
            .O(N__40761),
            .I(N__40758));
    LocalMux I__9214 (
            .O(N__40758),
            .I(\ppm_encoder_1.un1_init_pulses_10_17 ));
    InMux I__9213 (
            .O(N__40755),
            .I(N__40751));
    InMux I__9212 (
            .O(N__40754),
            .I(N__40748));
    LocalMux I__9211 (
            .O(N__40751),
            .I(N__40745));
    LocalMux I__9210 (
            .O(N__40748),
            .I(N__40742));
    Span4Mux_h I__9209 (
            .O(N__40745),
            .I(N__40738));
    Span4Mux_v I__9208 (
            .O(N__40742),
            .I(N__40735));
    InMux I__9207 (
            .O(N__40741),
            .I(N__40732));
    Span4Mux_h I__9206 (
            .O(N__40738),
            .I(N__40729));
    Odrv4 I__9205 (
            .O(N__40735),
            .I(\ppm_encoder_1.init_pulsesZ0Z_17 ));
    LocalMux I__9204 (
            .O(N__40732),
            .I(\ppm_encoder_1.init_pulsesZ0Z_17 ));
    Odrv4 I__9203 (
            .O(N__40729),
            .I(\ppm_encoder_1.init_pulsesZ0Z_17 ));
    CascadeMux I__9202 (
            .O(N__40722),
            .I(N__40719));
    InMux I__9201 (
            .O(N__40719),
            .I(N__40716));
    LocalMux I__9200 (
            .O(N__40716),
            .I(N__40713));
    Odrv4 I__9199 (
            .O(N__40713),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_7 ));
    InMux I__9198 (
            .O(N__40710),
            .I(N__40701));
    InMux I__9197 (
            .O(N__40709),
            .I(N__40701));
    InMux I__9196 (
            .O(N__40708),
            .I(N__40701));
    LocalMux I__9195 (
            .O(N__40701),
            .I(N__40698));
    Odrv4 I__9194 (
            .O(N__40698),
            .I(\ppm_encoder_1.init_pulsesZ0Z_7 ));
    InMux I__9193 (
            .O(N__40695),
            .I(N__40692));
    LocalMux I__9192 (
            .O(N__40692),
            .I(N__40687));
    InMux I__9191 (
            .O(N__40691),
            .I(N__40684));
    CascadeMux I__9190 (
            .O(N__40690),
            .I(N__40681));
    Span4Mux_v I__9189 (
            .O(N__40687),
            .I(N__40678));
    LocalMux I__9188 (
            .O(N__40684),
            .I(N__40675));
    InMux I__9187 (
            .O(N__40681),
            .I(N__40672));
    Span4Mux_h I__9186 (
            .O(N__40678),
            .I(N__40669));
    Span4Mux_h I__9185 (
            .O(N__40675),
            .I(N__40666));
    LocalMux I__9184 (
            .O(N__40672),
            .I(\ppm_encoder_1.rudderZ0Z_7 ));
    Odrv4 I__9183 (
            .O(N__40669),
            .I(\ppm_encoder_1.rudderZ0Z_7 ));
    Odrv4 I__9182 (
            .O(N__40666),
            .I(\ppm_encoder_1.rudderZ0Z_7 ));
    InMux I__9181 (
            .O(N__40659),
            .I(N__40656));
    LocalMux I__9180 (
            .O(N__40656),
            .I(N__40653));
    Odrv4 I__9179 (
            .O(N__40653),
            .I(\ppm_encoder_1.un1_init_pulses_11_8 ));
    InMux I__9178 (
            .O(N__40650),
            .I(N__40647));
    LocalMux I__9177 (
            .O(N__40647),
            .I(\ppm_encoder_1.un1_init_pulses_10_8 ));
    InMux I__9176 (
            .O(N__40644),
            .I(N__40641));
    LocalMux I__9175 (
            .O(N__40641),
            .I(N__40636));
    InMux I__9174 (
            .O(N__40640),
            .I(N__40633));
    InMux I__9173 (
            .O(N__40639),
            .I(N__40630));
    Odrv4 I__9172 (
            .O(N__40636),
            .I(\ppm_encoder_1.init_pulsesZ0Z_8 ));
    LocalMux I__9171 (
            .O(N__40633),
            .I(\ppm_encoder_1.init_pulsesZ0Z_8 ));
    LocalMux I__9170 (
            .O(N__40630),
            .I(\ppm_encoder_1.init_pulsesZ0Z_8 ));
    InMux I__9169 (
            .O(N__40623),
            .I(N__40619));
    CascadeMux I__9168 (
            .O(N__40622),
            .I(N__40616));
    LocalMux I__9167 (
            .O(N__40619),
            .I(N__40613));
    InMux I__9166 (
            .O(N__40616),
            .I(N__40610));
    Span4Mux_v I__9165 (
            .O(N__40613),
            .I(N__40607));
    LocalMux I__9164 (
            .O(N__40610),
            .I(N__40604));
    Odrv4 I__9163 (
            .O(N__40607),
            .I(\ppm_encoder_1.un1_init_pulses_0_8 ));
    Odrv4 I__9162 (
            .O(N__40604),
            .I(\ppm_encoder_1.un1_init_pulses_0_8 ));
    InMux I__9161 (
            .O(N__40599),
            .I(N__40596));
    LocalMux I__9160 (
            .O(N__40596),
            .I(\ppm_encoder_1.un1_init_pulses_10_9 ));
    InMux I__9159 (
            .O(N__40593),
            .I(N__40590));
    LocalMux I__9158 (
            .O(N__40590),
            .I(N__40587));
    Odrv12 I__9157 (
            .O(N__40587),
            .I(\ppm_encoder_1.un1_init_pulses_11_9 ));
    InMux I__9156 (
            .O(N__40584),
            .I(N__40581));
    LocalMux I__9155 (
            .O(N__40581),
            .I(N__40578));
    Odrv4 I__9154 (
            .O(N__40578),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_9 ));
    CascadeMux I__9153 (
            .O(N__40575),
            .I(N__40571));
    InMux I__9152 (
            .O(N__40574),
            .I(N__40568));
    InMux I__9151 (
            .O(N__40571),
            .I(N__40565));
    LocalMux I__9150 (
            .O(N__40568),
            .I(N__40562));
    LocalMux I__9149 (
            .O(N__40565),
            .I(N__40559));
    Odrv12 I__9148 (
            .O(N__40562),
            .I(\ppm_encoder_1.un1_init_pulses_0_9 ));
    Odrv4 I__9147 (
            .O(N__40559),
            .I(\ppm_encoder_1.un1_init_pulses_0_9 ));
    InMux I__9146 (
            .O(N__40554),
            .I(N__40545));
    InMux I__9145 (
            .O(N__40553),
            .I(N__40545));
    InMux I__9144 (
            .O(N__40552),
            .I(N__40545));
    LocalMux I__9143 (
            .O(N__40545),
            .I(\ppm_encoder_1.init_pulsesZ0Z_9 ));
    CascadeMux I__9142 (
            .O(N__40542),
            .I(N__40539));
    InMux I__9141 (
            .O(N__40539),
            .I(N__40536));
    LocalMux I__9140 (
            .O(N__40536),
            .I(N__40532));
    InMux I__9139 (
            .O(N__40535),
            .I(N__40528));
    Span12Mux_h I__9138 (
            .O(N__40532),
            .I(N__40525));
    InMux I__9137 (
            .O(N__40531),
            .I(N__40522));
    LocalMux I__9136 (
            .O(N__40528),
            .I(\ppm_encoder_1.rudderZ0Z_9 ));
    Odrv12 I__9135 (
            .O(N__40525),
            .I(\ppm_encoder_1.rudderZ0Z_9 ));
    LocalMux I__9134 (
            .O(N__40522),
            .I(\ppm_encoder_1.rudderZ0Z_9 ));
    InMux I__9133 (
            .O(N__40515),
            .I(N__40512));
    LocalMux I__9132 (
            .O(N__40512),
            .I(N__40509));
    Span4Mux_v I__9131 (
            .O(N__40509),
            .I(N__40506));
    Odrv4 I__9130 (
            .O(N__40506),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_9 ));
    InMux I__9129 (
            .O(N__40503),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_14 ));
    InMux I__9128 (
            .O(N__40500),
            .I(bfn_18_13_0_));
    InMux I__9127 (
            .O(N__40497),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_16 ));
    InMux I__9126 (
            .O(N__40494),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_17 ));
    InMux I__9125 (
            .O(N__40491),
            .I(N__40486));
    InMux I__9124 (
            .O(N__40490),
            .I(N__40482));
    InMux I__9123 (
            .O(N__40489),
            .I(N__40479));
    LocalMux I__9122 (
            .O(N__40486),
            .I(N__40476));
    InMux I__9121 (
            .O(N__40485),
            .I(N__40473));
    LocalMux I__9120 (
            .O(N__40482),
            .I(N__40468));
    LocalMux I__9119 (
            .O(N__40479),
            .I(N__40465));
    Span4Mux_v I__9118 (
            .O(N__40476),
            .I(N__40460));
    LocalMux I__9117 (
            .O(N__40473),
            .I(N__40460));
    InMux I__9116 (
            .O(N__40472),
            .I(N__40455));
    InMux I__9115 (
            .O(N__40471),
            .I(N__40455));
    Span4Mux_h I__9114 (
            .O(N__40468),
            .I(N__40451));
    Span4Mux_v I__9113 (
            .O(N__40465),
            .I(N__40448));
    Span4Mux_h I__9112 (
            .O(N__40460),
            .I(N__40443));
    LocalMux I__9111 (
            .O(N__40455),
            .I(N__40443));
    InMux I__9110 (
            .O(N__40454),
            .I(N__40440));
    Span4Mux_v I__9109 (
            .O(N__40451),
            .I(N__40437));
    Span4Mux_h I__9108 (
            .O(N__40448),
            .I(N__40432));
    Span4Mux_v I__9107 (
            .O(N__40443),
            .I(N__40432));
    LocalMux I__9106 (
            .O(N__40440),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1 ));
    Odrv4 I__9105 (
            .O(N__40437),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1 ));
    Odrv4 I__9104 (
            .O(N__40432),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1 ));
    InMux I__9103 (
            .O(N__40425),
            .I(N__40422));
    LocalMux I__9102 (
            .O(N__40422),
            .I(N__40418));
    InMux I__9101 (
            .O(N__40421),
            .I(N__40415));
    Span4Mux_h I__9100 (
            .O(N__40418),
            .I(N__40412));
    LocalMux I__9099 (
            .O(N__40415),
            .I(N__40409));
    Span4Mux_v I__9098 (
            .O(N__40412),
            .I(N__40403));
    Span4Mux_h I__9097 (
            .O(N__40409),
            .I(N__40400));
    InMux I__9096 (
            .O(N__40408),
            .I(N__40397));
    InMux I__9095 (
            .O(N__40407),
            .I(N__40392));
    InMux I__9094 (
            .O(N__40406),
            .I(N__40392));
    Odrv4 I__9093 (
            .O(N__40403),
            .I(\ppm_encoder_1.N_227 ));
    Odrv4 I__9092 (
            .O(N__40400),
            .I(\ppm_encoder_1.N_227 ));
    LocalMux I__9091 (
            .O(N__40397),
            .I(\ppm_encoder_1.N_227 ));
    LocalMux I__9090 (
            .O(N__40392),
            .I(\ppm_encoder_1.N_227 ));
    CascadeMux I__9089 (
            .O(N__40383),
            .I(N__40380));
    InMux I__9088 (
            .O(N__40380),
            .I(N__40374));
    CascadeMux I__9087 (
            .O(N__40379),
            .I(N__40370));
    CascadeMux I__9086 (
            .O(N__40378),
            .I(N__40367));
    CascadeMux I__9085 (
            .O(N__40377),
            .I(N__40364));
    LocalMux I__9084 (
            .O(N__40374),
            .I(N__40359));
    InMux I__9083 (
            .O(N__40373),
            .I(N__40352));
    InMux I__9082 (
            .O(N__40370),
            .I(N__40352));
    InMux I__9081 (
            .O(N__40367),
            .I(N__40352));
    InMux I__9080 (
            .O(N__40364),
            .I(N__40349));
    InMux I__9079 (
            .O(N__40363),
            .I(N__40346));
    InMux I__9078 (
            .O(N__40362),
            .I(N__40343));
    Span4Mux_h I__9077 (
            .O(N__40359),
            .I(N__40340));
    LocalMux I__9076 (
            .O(N__40352),
            .I(N__40337));
    LocalMux I__9075 (
            .O(N__40349),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1 ));
    LocalMux I__9074 (
            .O(N__40346),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1 ));
    LocalMux I__9073 (
            .O(N__40343),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1 ));
    Odrv4 I__9072 (
            .O(N__40340),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1 ));
    Odrv4 I__9071 (
            .O(N__40337),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1 ));
    InMux I__9070 (
            .O(N__40326),
            .I(N__40322));
    InMux I__9069 (
            .O(N__40325),
            .I(N__40318));
    LocalMux I__9068 (
            .O(N__40322),
            .I(N__40315));
    CascadeMux I__9067 (
            .O(N__40321),
            .I(N__40312));
    LocalMux I__9066 (
            .O(N__40318),
            .I(N__40309));
    Span4Mux_v I__9065 (
            .O(N__40315),
            .I(N__40306));
    InMux I__9064 (
            .O(N__40312),
            .I(N__40303));
    Span4Mux_h I__9063 (
            .O(N__40309),
            .I(N__40296));
    Span4Mux_v I__9062 (
            .O(N__40306),
            .I(N__40291));
    LocalMux I__9061 (
            .O(N__40303),
            .I(N__40291));
    InMux I__9060 (
            .O(N__40302),
            .I(N__40282));
    InMux I__9059 (
            .O(N__40301),
            .I(N__40282));
    InMux I__9058 (
            .O(N__40300),
            .I(N__40282));
    InMux I__9057 (
            .O(N__40299),
            .I(N__40282));
    Odrv4 I__9056 (
            .O(N__40296),
            .I(\ppm_encoder_1.PPM_STATEZ0Z_0 ));
    Odrv4 I__9055 (
            .O(N__40291),
            .I(\ppm_encoder_1.PPM_STATEZ0Z_0 ));
    LocalMux I__9054 (
            .O(N__40282),
            .I(\ppm_encoder_1.PPM_STATEZ0Z_0 ));
    CascadeMux I__9053 (
            .O(N__40275),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_1_0_cascade_ ));
    InMux I__9052 (
            .O(N__40272),
            .I(N__40269));
    LocalMux I__9051 (
            .O(N__40269),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_8 ));
    InMux I__9050 (
            .O(N__40266),
            .I(N__40263));
    LocalMux I__9049 (
            .O(N__40263),
            .I(N__40260));
    Odrv4 I__9048 (
            .O(N__40260),
            .I(\ppm_encoder_1.un1_init_pulses_11_7 ));
    InMux I__9047 (
            .O(N__40257),
            .I(N__40254));
    LocalMux I__9046 (
            .O(N__40254),
            .I(\ppm_encoder_1.un1_init_pulses_10_7 ));
    InMux I__9045 (
            .O(N__40251),
            .I(N__40248));
    LocalMux I__9044 (
            .O(N__40248),
            .I(N__40244));
    CascadeMux I__9043 (
            .O(N__40247),
            .I(N__40241));
    Span4Mux_h I__9042 (
            .O(N__40244),
            .I(N__40238));
    InMux I__9041 (
            .O(N__40241),
            .I(N__40235));
    Odrv4 I__9040 (
            .O(N__40238),
            .I(\ppm_encoder_1.un1_init_pulses_0_7 ));
    LocalMux I__9039 (
            .O(N__40235),
            .I(\ppm_encoder_1.un1_init_pulses_0_7 ));
    InMux I__9038 (
            .O(N__40230),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_6 ));
    InMux I__9037 (
            .O(N__40227),
            .I(bfn_18_12_0_));
    InMux I__9036 (
            .O(N__40224),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_8 ));
    InMux I__9035 (
            .O(N__40221),
            .I(N__40218));
    LocalMux I__9034 (
            .O(N__40218),
            .I(\ppm_encoder_1.un1_init_pulses_11_10 ));
    InMux I__9033 (
            .O(N__40215),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_9 ));
    InMux I__9032 (
            .O(N__40212),
            .I(N__40209));
    LocalMux I__9031 (
            .O(N__40209),
            .I(N__40206));
    Span4Mux_h I__9030 (
            .O(N__40206),
            .I(N__40203));
    Span4Mux_h I__9029 (
            .O(N__40203),
            .I(N__40200));
    Span4Mux_v I__9028 (
            .O(N__40200),
            .I(N__40197));
    Odrv4 I__9027 (
            .O(N__40197),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_11 ));
    InMux I__9026 (
            .O(N__40194),
            .I(N__40191));
    LocalMux I__9025 (
            .O(N__40191),
            .I(\ppm_encoder_1.un1_init_pulses_11_11 ));
    InMux I__9024 (
            .O(N__40188),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_10 ));
    InMux I__9023 (
            .O(N__40185),
            .I(N__40182));
    LocalMux I__9022 (
            .O(N__40182),
            .I(N__40179));
    Span12Mux_s11_h I__9021 (
            .O(N__40179),
            .I(N__40176));
    Odrv12 I__9020 (
            .O(N__40176),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_12 ));
    InMux I__9019 (
            .O(N__40173),
            .I(N__40170));
    LocalMux I__9018 (
            .O(N__40170),
            .I(\ppm_encoder_1.un1_init_pulses_11_12 ));
    InMux I__9017 (
            .O(N__40167),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_11 ));
    InMux I__9016 (
            .O(N__40164),
            .I(N__40161));
    LocalMux I__9015 (
            .O(N__40161),
            .I(\ppm_encoder_1.init_pulses_RNIUPKO2Z0Z_13 ));
    CascadeMux I__9014 (
            .O(N__40158),
            .I(N__40155));
    InMux I__9013 (
            .O(N__40155),
            .I(N__40152));
    LocalMux I__9012 (
            .O(N__40152),
            .I(N__40149));
    Odrv4 I__9011 (
            .O(N__40149),
            .I(\ppm_encoder_1.PPM_STATE_RNI2APU1Z0Z_1 ));
    InMux I__9010 (
            .O(N__40146),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_12 ));
    InMux I__9009 (
            .O(N__40143),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_13 ));
    InMux I__9008 (
            .O(N__40140),
            .I(N__40137));
    LocalMux I__9007 (
            .O(N__40137),
            .I(N__40122));
    InMux I__9006 (
            .O(N__40136),
            .I(N__40118));
    InMux I__9005 (
            .O(N__40135),
            .I(N__40115));
    InMux I__9004 (
            .O(N__40134),
            .I(N__40110));
    InMux I__9003 (
            .O(N__40133),
            .I(N__40105));
    InMux I__9002 (
            .O(N__40132),
            .I(N__40105));
    InMux I__9001 (
            .O(N__40131),
            .I(N__40102));
    InMux I__9000 (
            .O(N__40130),
            .I(N__40099));
    InMux I__8999 (
            .O(N__40129),
            .I(N__40096));
    InMux I__8998 (
            .O(N__40128),
            .I(N__40093));
    InMux I__8997 (
            .O(N__40127),
            .I(N__40088));
    InMux I__8996 (
            .O(N__40126),
            .I(N__40083));
    InMux I__8995 (
            .O(N__40125),
            .I(N__40083));
    Span4Mux_v I__8994 (
            .O(N__40122),
            .I(N__40080));
    InMux I__8993 (
            .O(N__40121),
            .I(N__40077));
    LocalMux I__8992 (
            .O(N__40118),
            .I(N__40072));
    LocalMux I__8991 (
            .O(N__40115),
            .I(N__40072));
    InMux I__8990 (
            .O(N__40114),
            .I(N__40069));
    InMux I__8989 (
            .O(N__40113),
            .I(N__40066));
    LocalMux I__8988 (
            .O(N__40110),
            .I(N__40059));
    LocalMux I__8987 (
            .O(N__40105),
            .I(N__40059));
    LocalMux I__8986 (
            .O(N__40102),
            .I(N__40059));
    LocalMux I__8985 (
            .O(N__40099),
            .I(N__40056));
    LocalMux I__8984 (
            .O(N__40096),
            .I(N__40052));
    LocalMux I__8983 (
            .O(N__40093),
            .I(N__40049));
    InMux I__8982 (
            .O(N__40092),
            .I(N__40044));
    InMux I__8981 (
            .O(N__40091),
            .I(N__40044));
    LocalMux I__8980 (
            .O(N__40088),
            .I(N__40041));
    LocalMux I__8979 (
            .O(N__40083),
            .I(N__40036));
    Span4Mux_v I__8978 (
            .O(N__40080),
            .I(N__40036));
    LocalMux I__8977 (
            .O(N__40077),
            .I(N__40033));
    Span4Mux_h I__8976 (
            .O(N__40072),
            .I(N__40022));
    LocalMux I__8975 (
            .O(N__40069),
            .I(N__40022));
    LocalMux I__8974 (
            .O(N__40066),
            .I(N__40022));
    Span4Mux_v I__8973 (
            .O(N__40059),
            .I(N__40022));
    Span4Mux_h I__8972 (
            .O(N__40056),
            .I(N__40022));
    InMux I__8971 (
            .O(N__40055),
            .I(N__40019));
    Span4Mux_v I__8970 (
            .O(N__40052),
            .I(N__40014));
    Span4Mux_v I__8969 (
            .O(N__40049),
            .I(N__40014));
    LocalMux I__8968 (
            .O(N__40044),
            .I(N__40007));
    Span4Mux_v I__8967 (
            .O(N__40041),
            .I(N__40007));
    Span4Mux_h I__8966 (
            .O(N__40036),
            .I(N__40007));
    Span4Mux_v I__8965 (
            .O(N__40033),
            .I(N__40002));
    Span4Mux_v I__8964 (
            .O(N__40022),
            .I(N__40002));
    LocalMux I__8963 (
            .O(N__40019),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_1 ));
    Odrv4 I__8962 (
            .O(N__40014),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_1 ));
    Odrv4 I__8961 (
            .O(N__40007),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_1 ));
    Odrv4 I__8960 (
            .O(N__40002),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_1 ));
    InMux I__8959 (
            .O(N__39993),
            .I(N__39988));
    InMux I__8958 (
            .O(N__39992),
            .I(N__39985));
    CascadeMux I__8957 (
            .O(N__39991),
            .I(N__39982));
    LocalMux I__8956 (
            .O(N__39988),
            .I(N__39976));
    LocalMux I__8955 (
            .O(N__39985),
            .I(N__39976));
    InMux I__8954 (
            .O(N__39982),
            .I(N__39971));
    InMux I__8953 (
            .O(N__39981),
            .I(N__39968));
    Span4Mux_h I__8952 (
            .O(N__39976),
            .I(N__39965));
    InMux I__8951 (
            .O(N__39975),
            .I(N__39960));
    InMux I__8950 (
            .O(N__39974),
            .I(N__39960));
    LocalMux I__8949 (
            .O(N__39971),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_3 ));
    LocalMux I__8948 (
            .O(N__39968),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_3 ));
    Odrv4 I__8947 (
            .O(N__39965),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_3 ));
    LocalMux I__8946 (
            .O(N__39960),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_3 ));
    InMux I__8945 (
            .O(N__39951),
            .I(N__39948));
    LocalMux I__8944 (
            .O(N__39948),
            .I(N__39945));
    Odrv12 I__8943 (
            .O(N__39945),
            .I(\ppm_encoder_1.PPM_STATE_RNI2APU1_2Z0Z_1 ));
    CascadeMux I__8942 (
            .O(N__39942),
            .I(N__39939));
    InMux I__8941 (
            .O(N__39939),
            .I(N__39936));
    LocalMux I__8940 (
            .O(N__39936),
            .I(N__39933));
    Odrv4 I__8939 (
            .O(N__39933),
            .I(\ppm_encoder_1.init_pulses_RNIAVNR2Z0Z_0 ));
    InMux I__8938 (
            .O(N__39930),
            .I(N__39927));
    LocalMux I__8937 (
            .O(N__39927),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_1 ));
    InMux I__8936 (
            .O(N__39924),
            .I(N__39921));
    LocalMux I__8935 (
            .O(N__39921),
            .I(\ppm_encoder_1.un1_init_pulses_11_1 ));
    InMux I__8934 (
            .O(N__39918),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_0 ));
    InMux I__8933 (
            .O(N__39915),
            .I(N__39912));
    LocalMux I__8932 (
            .O(N__39912),
            .I(N__39909));
    Odrv4 I__8931 (
            .O(N__39909),
            .I(\ppm_encoder_1.PPM_STATE_RNI2APU1_1Z0Z_1 ));
    CascadeMux I__8930 (
            .O(N__39906),
            .I(N__39903));
    InMux I__8929 (
            .O(N__39903),
            .I(N__39900));
    LocalMux I__8928 (
            .O(N__39900),
            .I(N__39897));
    Odrv4 I__8927 (
            .O(N__39897),
            .I(\ppm_encoder_1.init_pulses_RNIC1OR2Z0Z_2 ));
    InMux I__8926 (
            .O(N__39894),
            .I(N__39891));
    LocalMux I__8925 (
            .O(N__39891),
            .I(N__39888));
    Span4Mux_v I__8924 (
            .O(N__39888),
            .I(N__39885));
    Odrv4 I__8923 (
            .O(N__39885),
            .I(\ppm_encoder_1.un1_init_pulses_11_2 ));
    InMux I__8922 (
            .O(N__39882),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_1 ));
    InMux I__8921 (
            .O(N__39879),
            .I(N__39876));
    LocalMux I__8920 (
            .O(N__39876),
            .I(N__39873));
    Span4Mux_h I__8919 (
            .O(N__39873),
            .I(N__39870));
    Odrv4 I__8918 (
            .O(N__39870),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_3 ));
    InMux I__8917 (
            .O(N__39867),
            .I(N__39864));
    LocalMux I__8916 (
            .O(N__39864),
            .I(N__39861));
    Span4Mux_v I__8915 (
            .O(N__39861),
            .I(N__39858));
    Odrv4 I__8914 (
            .O(N__39858),
            .I(\ppm_encoder_1.un1_init_pulses_11_3 ));
    InMux I__8913 (
            .O(N__39855),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_2 ));
    InMux I__8912 (
            .O(N__39852),
            .I(N__39849));
    LocalMux I__8911 (
            .O(N__39849),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_4 ));
    InMux I__8910 (
            .O(N__39846),
            .I(N__39843));
    LocalMux I__8909 (
            .O(N__39843),
            .I(\ppm_encoder_1.un1_init_pulses_11_4 ));
    InMux I__8908 (
            .O(N__39840),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_3 ));
    InMux I__8907 (
            .O(N__39837),
            .I(N__39834));
    LocalMux I__8906 (
            .O(N__39834),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_5 ));
    InMux I__8905 (
            .O(N__39831),
            .I(N__39828));
    LocalMux I__8904 (
            .O(N__39828),
            .I(\ppm_encoder_1.un1_init_pulses_11_5 ));
    InMux I__8903 (
            .O(N__39825),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_4 ));
    InMux I__8902 (
            .O(N__39822),
            .I(N__39819));
    LocalMux I__8901 (
            .O(N__39819),
            .I(N__39816));
    Span4Mux_h I__8900 (
            .O(N__39816),
            .I(N__39813));
    Span4Mux_v I__8899 (
            .O(N__39813),
            .I(N__39810));
    Span4Mux_v I__8898 (
            .O(N__39810),
            .I(N__39807));
    Odrv4 I__8897 (
            .O(N__39807),
            .I(\ppm_encoder_1.PPM_STATE_RNI2APU1_0Z0Z_1 ));
    CascadeMux I__8896 (
            .O(N__39804),
            .I(N__39801));
    InMux I__8895 (
            .O(N__39801),
            .I(N__39798));
    LocalMux I__8894 (
            .O(N__39798),
            .I(N__39795));
    Odrv4 I__8893 (
            .O(N__39795),
            .I(\ppm_encoder_1.init_pulses_RNIG5OR2Z0Z_6 ));
    InMux I__8892 (
            .O(N__39792),
            .I(N__39789));
    LocalMux I__8891 (
            .O(N__39789),
            .I(N__39786));
    Odrv4 I__8890 (
            .O(N__39786),
            .I(\ppm_encoder_1.un1_init_pulses_11_6 ));
    InMux I__8889 (
            .O(N__39783),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_5 ));
    InMux I__8888 (
            .O(N__39780),
            .I(N__39777));
    LocalMux I__8887 (
            .O(N__39777),
            .I(N__39774));
    Span4Mux_v I__8886 (
            .O(N__39774),
            .I(N__39770));
    InMux I__8885 (
            .O(N__39773),
            .I(N__39767));
    Span4Mux_h I__8884 (
            .O(N__39770),
            .I(N__39764));
    LocalMux I__8883 (
            .O(N__39767),
            .I(\ppm_encoder_1.pulses2countZ0Z_16 ));
    Odrv4 I__8882 (
            .O(N__39764),
            .I(\ppm_encoder_1.pulses2countZ0Z_16 ));
    CascadeMux I__8881 (
            .O(N__39759),
            .I(N__39756));
    InMux I__8880 (
            .O(N__39756),
            .I(N__39750));
    InMux I__8879 (
            .O(N__39755),
            .I(N__39750));
    LocalMux I__8878 (
            .O(N__39750),
            .I(\ppm_encoder_1.pulses2countZ0Z_17 ));
    CascadeMux I__8877 (
            .O(N__39747),
            .I(N__39743));
    CascadeMux I__8876 (
            .O(N__39746),
            .I(N__39739));
    InMux I__8875 (
            .O(N__39743),
            .I(N__39731));
    InMux I__8874 (
            .O(N__39742),
            .I(N__39731));
    InMux I__8873 (
            .O(N__39739),
            .I(N__39731));
    CascadeMux I__8872 (
            .O(N__39738),
            .I(N__39728));
    LocalMux I__8871 (
            .O(N__39731),
            .I(N__39725));
    InMux I__8870 (
            .O(N__39728),
            .I(N__39722));
    Span4Mux_h I__8869 (
            .O(N__39725),
            .I(N__39719));
    LocalMux I__8868 (
            .O(N__39722),
            .I(N__39716));
    Span4Mux_v I__8867 (
            .O(N__39719),
            .I(N__39713));
    Span4Mux_h I__8866 (
            .O(N__39716),
            .I(N__39710));
    Span4Mux_v I__8865 (
            .O(N__39713),
            .I(N__39707));
    Span4Mux_v I__8864 (
            .O(N__39710),
            .I(N__39704));
    Odrv4 I__8863 (
            .O(N__39707),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_159_d ));
    Odrv4 I__8862 (
            .O(N__39704),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_159_d ));
    InMux I__8861 (
            .O(N__39699),
            .I(N__39694));
    InMux I__8860 (
            .O(N__39698),
            .I(N__39689));
    InMux I__8859 (
            .O(N__39697),
            .I(N__39689));
    LocalMux I__8858 (
            .O(N__39694),
            .I(\ppm_encoder_1.counterZ0Z_15 ));
    LocalMux I__8857 (
            .O(N__39689),
            .I(\ppm_encoder_1.counterZ0Z_15 ));
    InMux I__8856 (
            .O(N__39684),
            .I(N__39679));
    CascadeMux I__8855 (
            .O(N__39683),
            .I(N__39676));
    InMux I__8854 (
            .O(N__39682),
            .I(N__39673));
    LocalMux I__8853 (
            .O(N__39679),
            .I(N__39670));
    InMux I__8852 (
            .O(N__39676),
            .I(N__39667));
    LocalMux I__8851 (
            .O(N__39673),
            .I(\ppm_encoder_1.counterZ0Z_17 ));
    Odrv4 I__8850 (
            .O(N__39670),
            .I(\ppm_encoder_1.counterZ0Z_17 ));
    LocalMux I__8849 (
            .O(N__39667),
            .I(\ppm_encoder_1.counterZ0Z_17 ));
    CascadeMux I__8848 (
            .O(N__39660),
            .I(N__39656));
    InMux I__8847 (
            .O(N__39659),
            .I(N__39652));
    InMux I__8846 (
            .O(N__39656),
            .I(N__39647));
    InMux I__8845 (
            .O(N__39655),
            .I(N__39647));
    LocalMux I__8844 (
            .O(N__39652),
            .I(\ppm_encoder_1.counterZ0Z_16 ));
    LocalMux I__8843 (
            .O(N__39647),
            .I(\ppm_encoder_1.counterZ0Z_16 ));
    InMux I__8842 (
            .O(N__39642),
            .I(N__39638));
    InMux I__8841 (
            .O(N__39641),
            .I(N__39635));
    LocalMux I__8840 (
            .O(N__39638),
            .I(N__39630));
    LocalMux I__8839 (
            .O(N__39635),
            .I(N__39630));
    Span4Mux_h I__8838 (
            .O(N__39630),
            .I(N__39627));
    Odrv4 I__8837 (
            .O(N__39627),
            .I(\ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_4_0 ));
    InMux I__8836 (
            .O(N__39624),
            .I(N__39620));
    InMux I__8835 (
            .O(N__39623),
            .I(N__39617));
    LocalMux I__8834 (
            .O(N__39620),
            .I(\ppm_encoder_1.pulses2countZ0Z_18 ));
    LocalMux I__8833 (
            .O(N__39617),
            .I(\ppm_encoder_1.pulses2countZ0Z_18 ));
    InMux I__8832 (
            .O(N__39612),
            .I(N__39607));
    InMux I__8831 (
            .O(N__39611),
            .I(N__39604));
    InMux I__8830 (
            .O(N__39610),
            .I(N__39601));
    LocalMux I__8829 (
            .O(N__39607),
            .I(\ppm_encoder_1.counterZ0Z_18 ));
    LocalMux I__8828 (
            .O(N__39604),
            .I(\ppm_encoder_1.counterZ0Z_18 ));
    LocalMux I__8827 (
            .O(N__39601),
            .I(\ppm_encoder_1.counterZ0Z_18 ));
    InMux I__8826 (
            .O(N__39594),
            .I(N__39591));
    LocalMux I__8825 (
            .O(N__39591),
            .I(N__39588));
    Odrv12 I__8824 (
            .O(N__39588),
            .I(\pid_alt.O_0_4 ));
    CascadeMux I__8823 (
            .O(N__39585),
            .I(N__39582));
    InMux I__8822 (
            .O(N__39582),
            .I(N__39578));
    InMux I__8821 (
            .O(N__39581),
            .I(N__39575));
    LocalMux I__8820 (
            .O(N__39578),
            .I(N__39572));
    LocalMux I__8819 (
            .O(N__39575),
            .I(N__39569));
    Span4Mux_h I__8818 (
            .O(N__39572),
            .I(N__39566));
    Odrv4 I__8817 (
            .O(N__39569),
            .I(\pid_alt.error_i_regZ0Z_0 ));
    Odrv4 I__8816 (
            .O(N__39566),
            .I(\pid_alt.error_i_regZ0Z_0 ));
    InMux I__8815 (
            .O(N__39561),
            .I(N__39558));
    LocalMux I__8814 (
            .O(N__39558),
            .I(N__39555));
    Odrv12 I__8813 (
            .O(N__39555),
            .I(\pid_alt.O_0_7 ));
    CascadeMux I__8812 (
            .O(N__39552),
            .I(N__39549));
    InMux I__8811 (
            .O(N__39549),
            .I(N__39546));
    LocalMux I__8810 (
            .O(N__39546),
            .I(N__39543));
    Span4Mux_h I__8809 (
            .O(N__39543),
            .I(N__39540));
    Odrv4 I__8808 (
            .O(N__39540),
            .I(\pid_alt.error_i_regZ0Z_3 ));
    InMux I__8807 (
            .O(N__39537),
            .I(N__39534));
    LocalMux I__8806 (
            .O(N__39534),
            .I(\uart_drone.CO0 ));
    InMux I__8805 (
            .O(N__39531),
            .I(N__39527));
    InMux I__8804 (
            .O(N__39530),
            .I(N__39524));
    LocalMux I__8803 (
            .O(N__39527),
            .I(\uart_drone.un1_state_7_0 ));
    LocalMux I__8802 (
            .O(N__39524),
            .I(\uart_drone.un1_state_7_0 ));
    CascadeMux I__8801 (
            .O(N__39519),
            .I(N__39513));
    InMux I__8800 (
            .O(N__39518),
            .I(N__39509));
    InMux I__8799 (
            .O(N__39517),
            .I(N__39504));
    InMux I__8798 (
            .O(N__39516),
            .I(N__39504));
    InMux I__8797 (
            .O(N__39513),
            .I(N__39497));
    InMux I__8796 (
            .O(N__39512),
            .I(N__39497));
    LocalMux I__8795 (
            .O(N__39509),
            .I(N__39491));
    LocalMux I__8794 (
            .O(N__39504),
            .I(N__39488));
    InMux I__8793 (
            .O(N__39503),
            .I(N__39483));
    InMux I__8792 (
            .O(N__39502),
            .I(N__39483));
    LocalMux I__8791 (
            .O(N__39497),
            .I(N__39480));
    InMux I__8790 (
            .O(N__39496),
            .I(N__39477));
    InMux I__8789 (
            .O(N__39495),
            .I(N__39474));
    InMux I__8788 (
            .O(N__39494),
            .I(N__39471));
    Span12Mux_h I__8787 (
            .O(N__39491),
            .I(N__39468));
    Span12Mux_v I__8786 (
            .O(N__39488),
            .I(N__39463));
    LocalMux I__8785 (
            .O(N__39483),
            .I(N__39463));
    Span4Mux_v I__8784 (
            .O(N__39480),
            .I(N__39458));
    LocalMux I__8783 (
            .O(N__39477),
            .I(N__39458));
    LocalMux I__8782 (
            .O(N__39474),
            .I(\uart_drone.bit_CountZ0Z_1 ));
    LocalMux I__8781 (
            .O(N__39471),
            .I(\uart_drone.bit_CountZ0Z_1 ));
    Odrv12 I__8780 (
            .O(N__39468),
            .I(\uart_drone.bit_CountZ0Z_1 ));
    Odrv12 I__8779 (
            .O(N__39463),
            .I(\uart_drone.bit_CountZ0Z_1 ));
    Odrv4 I__8778 (
            .O(N__39458),
            .I(\uart_drone.bit_CountZ0Z_1 ));
    InMux I__8777 (
            .O(N__39447),
            .I(N__39444));
    LocalMux I__8776 (
            .O(N__39444),
            .I(N__39441));
    Span4Mux_h I__8775 (
            .O(N__39441),
            .I(N__39438));
    Span4Mux_v I__8774 (
            .O(N__39438),
            .I(N__39435));
    Odrv4 I__8773 (
            .O(N__39435),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_9 ));
    InMux I__8772 (
            .O(N__39432),
            .I(N__39429));
    LocalMux I__8771 (
            .O(N__39429),
            .I(N__39426));
    Span4Mux_v I__8770 (
            .O(N__39426),
            .I(N__39423));
    Span4Mux_h I__8769 (
            .O(N__39423),
            .I(N__39420));
    Odrv4 I__8768 (
            .O(N__39420),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_13 ));
    InMux I__8767 (
            .O(N__39417),
            .I(N__39414));
    LocalMux I__8766 (
            .O(N__39414),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_13 ));
    InMux I__8765 (
            .O(N__39411),
            .I(N__39408));
    LocalMux I__8764 (
            .O(N__39408),
            .I(N__39405));
    Span4Mux_v I__8763 (
            .O(N__39405),
            .I(N__39402));
    Odrv4 I__8762 (
            .O(N__39402),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_2 ));
    InMux I__8761 (
            .O(N__39399),
            .I(N__39396));
    LocalMux I__8760 (
            .O(N__39396),
            .I(N__39393));
    Span4Mux_v I__8759 (
            .O(N__39393),
            .I(N__39390));
    Odrv4 I__8758 (
            .O(N__39390),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_2 ));
    CascadeMux I__8757 (
            .O(N__39387),
            .I(N__39382));
    InMux I__8756 (
            .O(N__39386),
            .I(N__39378));
    InMux I__8755 (
            .O(N__39385),
            .I(N__39373));
    InMux I__8754 (
            .O(N__39382),
            .I(N__39373));
    InMux I__8753 (
            .O(N__39381),
            .I(N__39370));
    LocalMux I__8752 (
            .O(N__39378),
            .I(\ppm_encoder_1.counterZ0Z_3 ));
    LocalMux I__8751 (
            .O(N__39373),
            .I(\ppm_encoder_1.counterZ0Z_3 ));
    LocalMux I__8750 (
            .O(N__39370),
            .I(\ppm_encoder_1.counterZ0Z_3 ));
    InMux I__8749 (
            .O(N__39363),
            .I(N__39360));
    LocalMux I__8748 (
            .O(N__39360),
            .I(\ppm_encoder_1.pulses2countZ0Z_2 ));
    InMux I__8747 (
            .O(N__39357),
            .I(N__39351));
    InMux I__8746 (
            .O(N__39356),
            .I(N__39346));
    InMux I__8745 (
            .O(N__39355),
            .I(N__39346));
    InMux I__8744 (
            .O(N__39354),
            .I(N__39343));
    LocalMux I__8743 (
            .O(N__39351),
            .I(\ppm_encoder_1.counterZ0Z_2 ));
    LocalMux I__8742 (
            .O(N__39346),
            .I(\ppm_encoder_1.counterZ0Z_2 ));
    LocalMux I__8741 (
            .O(N__39343),
            .I(\ppm_encoder_1.counterZ0Z_2 ));
    InMux I__8740 (
            .O(N__39336),
            .I(N__39333));
    LocalMux I__8739 (
            .O(N__39333),
            .I(N__39330));
    Span4Mux_v I__8738 (
            .O(N__39330),
            .I(N__39327));
    Span4Mux_v I__8737 (
            .O(N__39327),
            .I(N__39324));
    Odrv4 I__8736 (
            .O(N__39324),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_3 ));
    InMux I__8735 (
            .O(N__39321),
            .I(N__39318));
    LocalMux I__8734 (
            .O(N__39318),
            .I(N__39315));
    Span4Mux_v I__8733 (
            .O(N__39315),
            .I(N__39312));
    Odrv4 I__8732 (
            .O(N__39312),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_3 ));
    CascadeMux I__8731 (
            .O(N__39309),
            .I(N__39306));
    InMux I__8730 (
            .O(N__39306),
            .I(N__39303));
    LocalMux I__8729 (
            .O(N__39303),
            .I(\ppm_encoder_1.pulses2countZ0Z_3 ));
    InMux I__8728 (
            .O(N__39300),
            .I(N__39297));
    LocalMux I__8727 (
            .O(N__39297),
            .I(\ppm_encoder_1.pulses2countZ0Z_8 ));
    CascadeMux I__8726 (
            .O(N__39294),
            .I(N__39290));
    InMux I__8725 (
            .O(N__39293),
            .I(N__39286));
    InMux I__8724 (
            .O(N__39290),
            .I(N__39283));
    InMux I__8723 (
            .O(N__39289),
            .I(N__39280));
    LocalMux I__8722 (
            .O(N__39286),
            .I(\ppm_encoder_1.counterZ0Z_9 ));
    LocalMux I__8721 (
            .O(N__39283),
            .I(\ppm_encoder_1.counterZ0Z_9 ));
    LocalMux I__8720 (
            .O(N__39280),
            .I(\ppm_encoder_1.counterZ0Z_9 ));
    CascadeMux I__8719 (
            .O(N__39273),
            .I(N__39270));
    InMux I__8718 (
            .O(N__39270),
            .I(N__39267));
    LocalMux I__8717 (
            .O(N__39267),
            .I(\ppm_encoder_1.pulses2countZ0Z_9 ));
    InMux I__8716 (
            .O(N__39264),
            .I(N__39259));
    InMux I__8715 (
            .O(N__39263),
            .I(N__39256));
    InMux I__8714 (
            .O(N__39262),
            .I(N__39253));
    LocalMux I__8713 (
            .O(N__39259),
            .I(\ppm_encoder_1.counterZ0Z_8 ));
    LocalMux I__8712 (
            .O(N__39256),
            .I(\ppm_encoder_1.counterZ0Z_8 ));
    LocalMux I__8711 (
            .O(N__39253),
            .I(\ppm_encoder_1.counterZ0Z_8 ));
    InMux I__8710 (
            .O(N__39246),
            .I(N__39241));
    InMux I__8709 (
            .O(N__39245),
            .I(N__39238));
    InMux I__8708 (
            .O(N__39244),
            .I(N__39235));
    LocalMux I__8707 (
            .O(N__39241),
            .I(\ppm_encoder_1.counterZ0Z_14 ));
    LocalMux I__8706 (
            .O(N__39238),
            .I(\ppm_encoder_1.counterZ0Z_14 ));
    LocalMux I__8705 (
            .O(N__39235),
            .I(\ppm_encoder_1.counterZ0Z_14 ));
    CascadeMux I__8704 (
            .O(N__39228),
            .I(N__39224));
    InMux I__8703 (
            .O(N__39227),
            .I(N__39219));
    InMux I__8702 (
            .O(N__39224),
            .I(N__39219));
    LocalMux I__8701 (
            .O(N__39219),
            .I(\ppm_encoder_1.pulses2countZ0Z_15 ));
    InMux I__8700 (
            .O(N__39216),
            .I(N__39213));
    LocalMux I__8699 (
            .O(N__39213),
            .I(N__39210));
    Span4Mux_v I__8698 (
            .O(N__39210),
            .I(N__39207));
    Span4Mux_h I__8697 (
            .O(N__39207),
            .I(N__39204));
    Span4Mux_h I__8696 (
            .O(N__39204),
            .I(N__39201));
    Span4Mux_v I__8695 (
            .O(N__39201),
            .I(N__39198));
    Odrv4 I__8694 (
            .O(N__39198),
            .I(\pid_alt.un9_error_filt_2_9 ));
    CascadeMux I__8693 (
            .O(N__39195),
            .I(N__39192));
    InMux I__8692 (
            .O(N__39192),
            .I(N__39189));
    LocalMux I__8691 (
            .O(N__39189),
            .I(N__39186));
    Span12Mux_h I__8690 (
            .O(N__39186),
            .I(N__39183));
    Odrv12 I__8689 (
            .O(N__39183),
            .I(\pid_alt.un9_error_filt_add_1_cry_9_sZ0 ));
    InMux I__8688 (
            .O(N__39180),
            .I(\pid_alt.un9_error_filt_add_1_cry_8 ));
    CascadeMux I__8687 (
            .O(N__39177),
            .I(N__39174));
    InMux I__8686 (
            .O(N__39174),
            .I(N__39171));
    LocalMux I__8685 (
            .O(N__39171),
            .I(N__39168));
    Span4Mux_h I__8684 (
            .O(N__39168),
            .I(N__39165));
    Span4Mux_h I__8683 (
            .O(N__39165),
            .I(N__39162));
    Span4Mux_v I__8682 (
            .O(N__39162),
            .I(N__39159));
    Odrv4 I__8681 (
            .O(N__39159),
            .I(\pid_alt.un9_error_filt_2_10 ));
    InMux I__8680 (
            .O(N__39156),
            .I(N__39153));
    LocalMux I__8679 (
            .O(N__39153),
            .I(N__39150));
    Span4Mux_s2_h I__8678 (
            .O(N__39150),
            .I(N__39147));
    Span4Mux_h I__8677 (
            .O(N__39147),
            .I(N__39144));
    Span4Mux_h I__8676 (
            .O(N__39144),
            .I(N__39141));
    Span4Mux_h I__8675 (
            .O(N__39141),
            .I(N__39138));
    Odrv4 I__8674 (
            .O(N__39138),
            .I(\pid_alt.un9_error_filt_add_1_cry_10_sZ0 ));
    InMux I__8673 (
            .O(N__39135),
            .I(\pid_alt.un9_error_filt_add_1_cry_9 ));
    CascadeMux I__8672 (
            .O(N__39132),
            .I(N__39127));
    InMux I__8671 (
            .O(N__39131),
            .I(N__39115));
    InMux I__8670 (
            .O(N__39130),
            .I(N__39115));
    InMux I__8669 (
            .O(N__39127),
            .I(N__39115));
    InMux I__8668 (
            .O(N__39126),
            .I(N__39115));
    CascadeMux I__8667 (
            .O(N__39125),
            .I(N__39112));
    CascadeMux I__8666 (
            .O(N__39124),
            .I(N__39108));
    LocalMux I__8665 (
            .O(N__39115),
            .I(N__39104));
    InMux I__8664 (
            .O(N__39112),
            .I(N__39095));
    InMux I__8663 (
            .O(N__39111),
            .I(N__39095));
    InMux I__8662 (
            .O(N__39108),
            .I(N__39095));
    InMux I__8661 (
            .O(N__39107),
            .I(N__39095));
    Span4Mux_v I__8660 (
            .O(N__39104),
            .I(N__39090));
    LocalMux I__8659 (
            .O(N__39095),
            .I(N__39090));
    Span4Mux_h I__8658 (
            .O(N__39090),
            .I(N__39087));
    Span4Mux_h I__8657 (
            .O(N__39087),
            .I(N__39084));
    Odrv4 I__8656 (
            .O(N__39084),
            .I(\pid_alt.un9_error_filt_1_19 ));
    InMux I__8655 (
            .O(N__39081),
            .I(N__39078));
    LocalMux I__8654 (
            .O(N__39078),
            .I(N__39075));
    Span4Mux_h I__8653 (
            .O(N__39075),
            .I(N__39072));
    Span4Mux_h I__8652 (
            .O(N__39072),
            .I(N__39069));
    Span4Mux_v I__8651 (
            .O(N__39069),
            .I(N__39066));
    Odrv4 I__8650 (
            .O(N__39066),
            .I(\pid_alt.un9_error_filt_2_11 ));
    InMux I__8649 (
            .O(N__39063),
            .I(\pid_alt.un9_error_filt_add_1_cry_10 ));
    CascadeMux I__8648 (
            .O(N__39060),
            .I(N__39056));
    InMux I__8647 (
            .O(N__39059),
            .I(N__39051));
    InMux I__8646 (
            .O(N__39056),
            .I(N__39051));
    LocalMux I__8645 (
            .O(N__39051),
            .I(N__39048));
    Span12Mux_s10_h I__8644 (
            .O(N__39048),
            .I(N__39045));
    Odrv12 I__8643 (
            .O(N__39045),
            .I(\pid_alt.un9_error_filt_add_1_sZ0Z_11 ));
    InMux I__8642 (
            .O(N__39042),
            .I(N__39039));
    LocalMux I__8641 (
            .O(N__39039),
            .I(N__39036));
    Span4Mux_h I__8640 (
            .O(N__39036),
            .I(N__39033));
    Odrv4 I__8639 (
            .O(N__39033),
            .I(\ppm_encoder_1.N_140_0 ));
    InMux I__8638 (
            .O(N__39030),
            .I(N__39026));
    CascadeMux I__8637 (
            .O(N__39029),
            .I(N__39023));
    LocalMux I__8636 (
            .O(N__39026),
            .I(N__39020));
    InMux I__8635 (
            .O(N__39023),
            .I(N__39017));
    Span4Mux_v I__8634 (
            .O(N__39020),
            .I(N__39014));
    LocalMux I__8633 (
            .O(N__39017),
            .I(N__39011));
    Odrv4 I__8632 (
            .O(N__39014),
            .I(\ppm_encoder_1.un1_init_pulses_0_10 ));
    Odrv12 I__8631 (
            .O(N__39011),
            .I(\ppm_encoder_1.un1_init_pulses_0_10 ));
    InMux I__8630 (
            .O(N__39006),
            .I(N__39002));
    InMux I__8629 (
            .O(N__39005),
            .I(N__38998));
    LocalMux I__8628 (
            .O(N__39002),
            .I(N__38995));
    InMux I__8627 (
            .O(N__39001),
            .I(N__38992));
    LocalMux I__8626 (
            .O(N__38998),
            .I(\ppm_encoder_1.rudderZ0Z_13 ));
    Odrv4 I__8625 (
            .O(N__38995),
            .I(\ppm_encoder_1.rudderZ0Z_13 ));
    LocalMux I__8624 (
            .O(N__38992),
            .I(\ppm_encoder_1.rudderZ0Z_13 ));
    CascadeMux I__8623 (
            .O(N__38985),
            .I(N__38980));
    CascadeMux I__8622 (
            .O(N__38984),
            .I(N__38977));
    InMux I__8621 (
            .O(N__38983),
            .I(N__38968));
    InMux I__8620 (
            .O(N__38980),
            .I(N__38965));
    InMux I__8619 (
            .O(N__38977),
            .I(N__38958));
    InMux I__8618 (
            .O(N__38976),
            .I(N__38958));
    InMux I__8617 (
            .O(N__38975),
            .I(N__38958));
    InMux I__8616 (
            .O(N__38974),
            .I(N__38953));
    InMux I__8615 (
            .O(N__38973),
            .I(N__38953));
    InMux I__8614 (
            .O(N__38972),
            .I(N__38950));
    CascadeMux I__8613 (
            .O(N__38971),
            .I(N__38942));
    LocalMux I__8612 (
            .O(N__38968),
            .I(N__38939));
    LocalMux I__8611 (
            .O(N__38965),
            .I(N__38932));
    LocalMux I__8610 (
            .O(N__38958),
            .I(N__38932));
    LocalMux I__8609 (
            .O(N__38953),
            .I(N__38932));
    LocalMux I__8608 (
            .O(N__38950),
            .I(N__38929));
    InMux I__8607 (
            .O(N__38949),
            .I(N__38926));
    InMux I__8606 (
            .O(N__38948),
            .I(N__38922));
    InMux I__8605 (
            .O(N__38947),
            .I(N__38919));
    CascadeMux I__8604 (
            .O(N__38946),
            .I(N__38913));
    InMux I__8603 (
            .O(N__38945),
            .I(N__38910));
    InMux I__8602 (
            .O(N__38942),
            .I(N__38907));
    Span4Mux_h I__8601 (
            .O(N__38939),
            .I(N__38898));
    Span4Mux_v I__8600 (
            .O(N__38932),
            .I(N__38898));
    Span4Mux_h I__8599 (
            .O(N__38929),
            .I(N__38898));
    LocalMux I__8598 (
            .O(N__38926),
            .I(N__38898));
    InMux I__8597 (
            .O(N__38925),
            .I(N__38895));
    LocalMux I__8596 (
            .O(N__38922),
            .I(N__38892));
    LocalMux I__8595 (
            .O(N__38919),
            .I(N__38889));
    InMux I__8594 (
            .O(N__38918),
            .I(N__38886));
    InMux I__8593 (
            .O(N__38917),
            .I(N__38879));
    InMux I__8592 (
            .O(N__38916),
            .I(N__38879));
    InMux I__8591 (
            .O(N__38913),
            .I(N__38879));
    LocalMux I__8590 (
            .O(N__38910),
            .I(N__38876));
    LocalMux I__8589 (
            .O(N__38907),
            .I(N__38869));
    Span4Mux_v I__8588 (
            .O(N__38898),
            .I(N__38869));
    LocalMux I__8587 (
            .O(N__38895),
            .I(N__38869));
    Span4Mux_v I__8586 (
            .O(N__38892),
            .I(N__38864));
    Span4Mux_v I__8585 (
            .O(N__38889),
            .I(N__38864));
    LocalMux I__8584 (
            .O(N__38886),
            .I(N__38861));
    LocalMux I__8583 (
            .O(N__38879),
            .I(N__38852));
    Span4Mux_v I__8582 (
            .O(N__38876),
            .I(N__38852));
    Span4Mux_h I__8581 (
            .O(N__38869),
            .I(N__38849));
    Span4Mux_v I__8580 (
            .O(N__38864),
            .I(N__38844));
    Span4Mux_h I__8579 (
            .O(N__38861),
            .I(N__38844));
    InMux I__8578 (
            .O(N__38860),
            .I(N__38841));
    InMux I__8577 (
            .O(N__38859),
            .I(N__38834));
    InMux I__8576 (
            .O(N__38858),
            .I(N__38834));
    InMux I__8575 (
            .O(N__38857),
            .I(N__38834));
    Odrv4 I__8574 (
            .O(N__38852),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_0 ));
    Odrv4 I__8573 (
            .O(N__38849),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_0 ));
    Odrv4 I__8572 (
            .O(N__38844),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_0 ));
    LocalMux I__8571 (
            .O(N__38841),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_0 ));
    LocalMux I__8570 (
            .O(N__38834),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_0 ));
    InMux I__8569 (
            .O(N__38823),
            .I(N__38820));
    LocalMux I__8568 (
            .O(N__38820),
            .I(N__38817));
    Span4Mux_h I__8567 (
            .O(N__38817),
            .I(N__38814));
    Span4Mux_v I__8566 (
            .O(N__38814),
            .I(N__38811));
    Odrv4 I__8565 (
            .O(N__38811),
            .I(\ppm_encoder_1.N_300 ));
    InMux I__8564 (
            .O(N__38808),
            .I(N__38805));
    LocalMux I__8563 (
            .O(N__38805),
            .I(N__38802));
    Span4Mux_v I__8562 (
            .O(N__38802),
            .I(N__38797));
    InMux I__8561 (
            .O(N__38801),
            .I(N__38792));
    InMux I__8560 (
            .O(N__38800),
            .I(N__38792));
    Odrv4 I__8559 (
            .O(N__38797),
            .I(\ppm_encoder_1.aileronZ0Z_8 ));
    LocalMux I__8558 (
            .O(N__38792),
            .I(\ppm_encoder_1.aileronZ0Z_8 ));
    CascadeMux I__8557 (
            .O(N__38787),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_8_cascade_ ));
    InMux I__8556 (
            .O(N__38784),
            .I(N__38781));
    LocalMux I__8555 (
            .O(N__38781),
            .I(N__38778));
    Odrv4 I__8554 (
            .O(N__38778),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_8 ));
    InMux I__8553 (
            .O(N__38775),
            .I(N__38772));
    LocalMux I__8552 (
            .O(N__38772),
            .I(N__38769));
    Span4Mux_h I__8551 (
            .O(N__38769),
            .I(N__38766));
    Span4Mux_h I__8550 (
            .O(N__38766),
            .I(N__38763));
    Odrv4 I__8549 (
            .O(N__38763),
            .I(\pid_alt.un9_error_filt_1_17 ));
    CascadeMux I__8548 (
            .O(N__38760),
            .I(N__38757));
    InMux I__8547 (
            .O(N__38757),
            .I(N__38754));
    LocalMux I__8546 (
            .O(N__38754),
            .I(N__38751));
    Span4Mux_h I__8545 (
            .O(N__38751),
            .I(N__38748));
    Span4Mux_h I__8544 (
            .O(N__38748),
            .I(N__38745));
    Span4Mux_v I__8543 (
            .O(N__38745),
            .I(N__38742));
    Odrv4 I__8542 (
            .O(N__38742),
            .I(\pid_alt.un9_error_filt_2_2 ));
    InMux I__8541 (
            .O(N__38739),
            .I(N__38736));
    LocalMux I__8540 (
            .O(N__38736),
            .I(N__38733));
    Span4Mux_s2_h I__8539 (
            .O(N__38733),
            .I(N__38730));
    Span4Mux_h I__8538 (
            .O(N__38730),
            .I(N__38727));
    Span4Mux_h I__8537 (
            .O(N__38727),
            .I(N__38724));
    Span4Mux_h I__8536 (
            .O(N__38724),
            .I(N__38721));
    Odrv4 I__8535 (
            .O(N__38721),
            .I(\pid_alt.un9_error_filt_add_1_cry_2_sZ0 ));
    InMux I__8534 (
            .O(N__38718),
            .I(\pid_alt.un9_error_filt_add_1_cry_1 ));
    InMux I__8533 (
            .O(N__38715),
            .I(N__38712));
    LocalMux I__8532 (
            .O(N__38712),
            .I(N__38709));
    Span4Mux_h I__8531 (
            .O(N__38709),
            .I(N__38706));
    Span4Mux_h I__8530 (
            .O(N__38706),
            .I(N__38703));
    Odrv4 I__8529 (
            .O(N__38703),
            .I(\pid_alt.un9_error_filt_1_18 ));
    CascadeMux I__8528 (
            .O(N__38700),
            .I(N__38697));
    InMux I__8527 (
            .O(N__38697),
            .I(N__38694));
    LocalMux I__8526 (
            .O(N__38694),
            .I(N__38691));
    Span4Mux_h I__8525 (
            .O(N__38691),
            .I(N__38688));
    Span4Mux_h I__8524 (
            .O(N__38688),
            .I(N__38685));
    Span4Mux_v I__8523 (
            .O(N__38685),
            .I(N__38682));
    Odrv4 I__8522 (
            .O(N__38682),
            .I(\pid_alt.un9_error_filt_2_3 ));
    InMux I__8521 (
            .O(N__38679),
            .I(N__38676));
    LocalMux I__8520 (
            .O(N__38676),
            .I(N__38673));
    Span4Mux_s2_h I__8519 (
            .O(N__38673),
            .I(N__38670));
    Span4Mux_h I__8518 (
            .O(N__38670),
            .I(N__38667));
    Span4Mux_h I__8517 (
            .O(N__38667),
            .I(N__38664));
    Span4Mux_h I__8516 (
            .O(N__38664),
            .I(N__38661));
    Odrv4 I__8515 (
            .O(N__38661),
            .I(\pid_alt.un9_error_filt_add_1_cry_3_sZ0 ));
    InMux I__8514 (
            .O(N__38658),
            .I(\pid_alt.un9_error_filt_add_1_cry_2 ));
    CascadeMux I__8513 (
            .O(N__38655),
            .I(N__38652));
    InMux I__8512 (
            .O(N__38652),
            .I(N__38649));
    LocalMux I__8511 (
            .O(N__38649),
            .I(N__38646));
    Span12Mux_v I__8510 (
            .O(N__38646),
            .I(N__38643));
    Odrv12 I__8509 (
            .O(N__38643),
            .I(\pid_alt.un9_error_filt_2_4 ));
    CascadeMux I__8508 (
            .O(N__38640),
            .I(N__38637));
    InMux I__8507 (
            .O(N__38637),
            .I(N__38634));
    LocalMux I__8506 (
            .O(N__38634),
            .I(N__38631));
    Span12Mux_s9_h I__8505 (
            .O(N__38631),
            .I(N__38628));
    Odrv12 I__8504 (
            .O(N__38628),
            .I(\pid_alt.un9_error_filt_add_1_cry_4_sZ0 ));
    InMux I__8503 (
            .O(N__38625),
            .I(\pid_alt.un9_error_filt_add_1_cry_3 ));
    InMux I__8502 (
            .O(N__38622),
            .I(N__38619));
    LocalMux I__8501 (
            .O(N__38619),
            .I(N__38616));
    Span4Mux_h I__8500 (
            .O(N__38616),
            .I(N__38613));
    Span4Mux_h I__8499 (
            .O(N__38613),
            .I(N__38610));
    Span4Mux_v I__8498 (
            .O(N__38610),
            .I(N__38607));
    Odrv4 I__8497 (
            .O(N__38607),
            .I(\pid_alt.un9_error_filt_2_5 ));
    InMux I__8496 (
            .O(N__38604),
            .I(N__38601));
    LocalMux I__8495 (
            .O(N__38601),
            .I(N__38598));
    Span12Mux_s8_h I__8494 (
            .O(N__38598),
            .I(N__38595));
    Odrv12 I__8493 (
            .O(N__38595),
            .I(\pid_alt.un9_error_filt_add_1_cry_5_sZ0 ));
    InMux I__8492 (
            .O(N__38592),
            .I(\pid_alt.un9_error_filt_add_1_cry_4 ));
    CascadeMux I__8491 (
            .O(N__38589),
            .I(N__38586));
    InMux I__8490 (
            .O(N__38586),
            .I(N__38583));
    LocalMux I__8489 (
            .O(N__38583),
            .I(N__38580));
    Span4Mux_v I__8488 (
            .O(N__38580),
            .I(N__38577));
    Span4Mux_h I__8487 (
            .O(N__38577),
            .I(N__38574));
    Span4Mux_h I__8486 (
            .O(N__38574),
            .I(N__38571));
    Odrv4 I__8485 (
            .O(N__38571),
            .I(\pid_alt.un9_error_filt_2_6 ));
    InMux I__8484 (
            .O(N__38568),
            .I(N__38565));
    LocalMux I__8483 (
            .O(N__38565),
            .I(N__38562));
    Span4Mux_h I__8482 (
            .O(N__38562),
            .I(N__38559));
    Span4Mux_h I__8481 (
            .O(N__38559),
            .I(N__38556));
    Span4Mux_h I__8480 (
            .O(N__38556),
            .I(N__38553));
    Span4Mux_h I__8479 (
            .O(N__38553),
            .I(N__38550));
    Odrv4 I__8478 (
            .O(N__38550),
            .I(\pid_alt.un9_error_filt_add_1_cry_6_sZ0 ));
    InMux I__8477 (
            .O(N__38547),
            .I(\pid_alt.un9_error_filt_add_1_cry_5 ));
    InMux I__8476 (
            .O(N__38544),
            .I(N__38541));
    LocalMux I__8475 (
            .O(N__38541),
            .I(N__38538));
    Span4Mux_h I__8474 (
            .O(N__38538),
            .I(N__38535));
    Span4Mux_h I__8473 (
            .O(N__38535),
            .I(N__38532));
    Span4Mux_v I__8472 (
            .O(N__38532),
            .I(N__38529));
    Odrv4 I__8471 (
            .O(N__38529),
            .I(\pid_alt.un9_error_filt_2_7 ));
    CascadeMux I__8470 (
            .O(N__38526),
            .I(N__38523));
    InMux I__8469 (
            .O(N__38523),
            .I(N__38520));
    LocalMux I__8468 (
            .O(N__38520),
            .I(N__38517));
    Span4Mux_h I__8467 (
            .O(N__38517),
            .I(N__38514));
    Span4Mux_h I__8466 (
            .O(N__38514),
            .I(N__38511));
    Span4Mux_h I__8465 (
            .O(N__38511),
            .I(N__38508));
    Span4Mux_h I__8464 (
            .O(N__38508),
            .I(N__38505));
    Odrv4 I__8463 (
            .O(N__38505),
            .I(\pid_alt.un9_error_filt_add_1_cry_7_sZ0 ));
    InMux I__8462 (
            .O(N__38502),
            .I(\pid_alt.un9_error_filt_add_1_cry_6 ));
    CascadeMux I__8461 (
            .O(N__38499),
            .I(N__38496));
    InMux I__8460 (
            .O(N__38496),
            .I(N__38493));
    LocalMux I__8459 (
            .O(N__38493),
            .I(N__38490));
    Span4Mux_v I__8458 (
            .O(N__38490),
            .I(N__38487));
    Span4Mux_h I__8457 (
            .O(N__38487),
            .I(N__38484));
    Span4Mux_h I__8456 (
            .O(N__38484),
            .I(N__38481));
    Span4Mux_v I__8455 (
            .O(N__38481),
            .I(N__38478));
    Odrv4 I__8454 (
            .O(N__38478),
            .I(\pid_alt.un9_error_filt_2_8 ));
    InMux I__8453 (
            .O(N__38475),
            .I(N__38472));
    LocalMux I__8452 (
            .O(N__38472),
            .I(N__38469));
    Span4Mux_s3_h I__8451 (
            .O(N__38469),
            .I(N__38466));
    Span4Mux_h I__8450 (
            .O(N__38466),
            .I(N__38463));
    Span4Mux_h I__8449 (
            .O(N__38463),
            .I(N__38460));
    Span4Mux_h I__8448 (
            .O(N__38460),
            .I(N__38457));
    Odrv4 I__8447 (
            .O(N__38457),
            .I(\pid_alt.un9_error_filt_add_1_cry_8_sZ0 ));
    InMux I__8446 (
            .O(N__38454),
            .I(bfn_17_18_0_));
    CascadeMux I__8445 (
            .O(N__38451),
            .I(N__38448));
    InMux I__8444 (
            .O(N__38448),
            .I(N__38445));
    LocalMux I__8443 (
            .O(N__38445),
            .I(N__38442));
    Span4Mux_h I__8442 (
            .O(N__38442),
            .I(N__38439));
    Span4Mux_h I__8441 (
            .O(N__38439),
            .I(N__38436));
    Odrv4 I__8440 (
            .O(N__38436),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI7O1NZ0Z_2 ));
    InMux I__8439 (
            .O(N__38433),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_14 ));
    InMux I__8438 (
            .O(N__38430),
            .I(bfn_17_16_0_));
    InMux I__8437 (
            .O(N__38427),
            .I(N__38424));
    LocalMux I__8436 (
            .O(N__38424),
            .I(N__38421));
    Span4Mux_h I__8435 (
            .O(N__38421),
            .I(N__38418));
    Span4Mux_h I__8434 (
            .O(N__38418),
            .I(N__38415));
    Odrv4 I__8433 (
            .O(N__38415),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_17 ));
    InMux I__8432 (
            .O(N__38412),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_16 ));
    InMux I__8431 (
            .O(N__38409),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_17 ));
    InMux I__8430 (
            .O(N__38406),
            .I(N__38402));
    InMux I__8429 (
            .O(N__38405),
            .I(N__38398));
    LocalMux I__8428 (
            .O(N__38402),
            .I(N__38395));
    InMux I__8427 (
            .O(N__38401),
            .I(N__38392));
    LocalMux I__8426 (
            .O(N__38398),
            .I(N__38387));
    Span4Mux_v I__8425 (
            .O(N__38395),
            .I(N__38387));
    LocalMux I__8424 (
            .O(N__38392),
            .I(N__38384));
    Odrv4 I__8423 (
            .O(N__38387),
            .I(\ppm_encoder_1.rudderZ0Z_8 ));
    Odrv12 I__8422 (
            .O(N__38384),
            .I(\ppm_encoder_1.rudderZ0Z_8 ));
    InMux I__8421 (
            .O(N__38379),
            .I(N__38376));
    LocalMux I__8420 (
            .O(N__38376),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_16 ));
    InMux I__8419 (
            .O(N__38373),
            .I(N__38369));
    InMux I__8418 (
            .O(N__38372),
            .I(N__38366));
    LocalMux I__8417 (
            .O(N__38369),
            .I(N__38363));
    LocalMux I__8416 (
            .O(N__38366),
            .I(\ppm_encoder_1.aileronZ0Z_14 ));
    Odrv4 I__8415 (
            .O(N__38363),
            .I(\ppm_encoder_1.aileronZ0Z_14 ));
    InMux I__8414 (
            .O(N__38358),
            .I(N__38355));
    LocalMux I__8413 (
            .O(N__38355),
            .I(N__38352));
    Odrv4 I__8412 (
            .O(N__38352),
            .I(\ppm_encoder_1.N_306 ));
    InMux I__8411 (
            .O(N__38349),
            .I(N__38346));
    LocalMux I__8410 (
            .O(N__38346),
            .I(N__38343));
    Span4Mux_h I__8409 (
            .O(N__38343),
            .I(N__38340));
    Span4Mux_h I__8408 (
            .O(N__38340),
            .I(N__38337));
    Odrv4 I__8407 (
            .O(N__38337),
            .I(\pid_alt.un9_error_filt_1_15 ));
    CascadeMux I__8406 (
            .O(N__38334),
            .I(N__38331));
    InMux I__8405 (
            .O(N__38331),
            .I(N__38328));
    LocalMux I__8404 (
            .O(N__38328),
            .I(N__38325));
    Span4Mux_v I__8403 (
            .O(N__38325),
            .I(N__38322));
    Span4Mux_h I__8402 (
            .O(N__38322),
            .I(N__38319));
    Span4Mux_h I__8401 (
            .O(N__38319),
            .I(N__38316));
    Span4Mux_v I__8400 (
            .O(N__38316),
            .I(N__38313));
    Odrv4 I__8399 (
            .O(N__38313),
            .I(\pid_alt.un9_error_filt_2_0 ));
    InMux I__8398 (
            .O(N__38310),
            .I(N__38307));
    LocalMux I__8397 (
            .O(N__38307),
            .I(N__38304));
    Span4Mux_h I__8396 (
            .O(N__38304),
            .I(N__38301));
    Span4Mux_h I__8395 (
            .O(N__38301),
            .I(N__38298));
    Span4Mux_h I__8394 (
            .O(N__38298),
            .I(N__38295));
    Span4Mux_h I__8393 (
            .O(N__38295),
            .I(N__38292));
    Odrv4 I__8392 (
            .O(N__38292),
            .I(\pid_alt.un9_error_filt_add_1_axbZ0Z_0 ));
    InMux I__8391 (
            .O(N__38289),
            .I(N__38286));
    LocalMux I__8390 (
            .O(N__38286),
            .I(N__38283));
    Span4Mux_h I__8389 (
            .O(N__38283),
            .I(N__38280));
    Span4Mux_h I__8388 (
            .O(N__38280),
            .I(N__38277));
    Odrv4 I__8387 (
            .O(N__38277),
            .I(\pid_alt.un9_error_filt_1_16 ));
    CascadeMux I__8386 (
            .O(N__38274),
            .I(N__38271));
    InMux I__8385 (
            .O(N__38271),
            .I(N__38268));
    LocalMux I__8384 (
            .O(N__38268),
            .I(N__38265));
    Span4Mux_v I__8383 (
            .O(N__38265),
            .I(N__38262));
    Span4Mux_h I__8382 (
            .O(N__38262),
            .I(N__38259));
    Span4Mux_h I__8381 (
            .O(N__38259),
            .I(N__38256));
    Span4Mux_v I__8380 (
            .O(N__38256),
            .I(N__38253));
    Odrv4 I__8379 (
            .O(N__38253),
            .I(\pid_alt.un9_error_filt_2_1 ));
    InMux I__8378 (
            .O(N__38250),
            .I(N__38247));
    LocalMux I__8377 (
            .O(N__38247),
            .I(N__38244));
    Span4Mux_s3_h I__8376 (
            .O(N__38244),
            .I(N__38241));
    Span4Mux_h I__8375 (
            .O(N__38241),
            .I(N__38238));
    Span4Mux_h I__8374 (
            .O(N__38238),
            .I(N__38235));
    Span4Mux_h I__8373 (
            .O(N__38235),
            .I(N__38232));
    Odrv4 I__8372 (
            .O(N__38232),
            .I(\pid_alt.un9_error_filt_add_1_cry_1_sZ0 ));
    InMux I__8371 (
            .O(N__38229),
            .I(\pid_alt.un9_error_filt_add_1_cry_0 ));
    InMux I__8370 (
            .O(N__38226),
            .I(N__38223));
    LocalMux I__8369 (
            .O(N__38223),
            .I(N__38220));
    Span4Mux_h I__8368 (
            .O(N__38220),
            .I(N__38217));
    Odrv4 I__8367 (
            .O(N__38217),
            .I(\ppm_encoder_1.throttle_RNIJII96Z0Z_7 ));
    InMux I__8366 (
            .O(N__38214),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_6 ));
    InMux I__8365 (
            .O(N__38211),
            .I(N__38208));
    LocalMux I__8364 (
            .O(N__38208),
            .I(N__38205));
    Odrv4 I__8363 (
            .O(N__38205),
            .I(\ppm_encoder_1.throttle_RNIONI96Z0Z_8 ));
    InMux I__8362 (
            .O(N__38202),
            .I(bfn_17_15_0_));
    InMux I__8361 (
            .O(N__38199),
            .I(N__38196));
    LocalMux I__8360 (
            .O(N__38196),
            .I(N__38193));
    Odrv4 I__8359 (
            .O(N__38193),
            .I(\ppm_encoder_1.throttle_RNITSI96Z0Z_9 ));
    InMux I__8358 (
            .O(N__38190),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_8 ));
    InMux I__8357 (
            .O(N__38187),
            .I(N__38184));
    LocalMux I__8356 (
            .O(N__38184),
            .I(N__38181));
    Span4Mux_h I__8355 (
            .O(N__38181),
            .I(N__38178));
    Odrv4 I__8354 (
            .O(N__38178),
            .I(\ppm_encoder_1.elevator_RNI5GRT5Z0Z_10 ));
    InMux I__8353 (
            .O(N__38175),
            .I(N__38172));
    LocalMux I__8352 (
            .O(N__38172),
            .I(N__38169));
    Odrv4 I__8351 (
            .O(N__38169),
            .I(\ppm_encoder_1.un1_init_pulses_10_10 ));
    InMux I__8350 (
            .O(N__38166),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_9 ));
    InMux I__8349 (
            .O(N__38163),
            .I(N__38160));
    LocalMux I__8348 (
            .O(N__38160),
            .I(N__38157));
    Span4Mux_h I__8347 (
            .O(N__38157),
            .I(N__38154));
    Odrv4 I__8346 (
            .O(N__38154),
            .I(\ppm_encoder_1.elevator_RNIALRT5Z0Z_11 ));
    CascadeMux I__8345 (
            .O(N__38151),
            .I(N__38148));
    InMux I__8344 (
            .O(N__38148),
            .I(N__38145));
    LocalMux I__8343 (
            .O(N__38145),
            .I(N__38141));
    InMux I__8342 (
            .O(N__38144),
            .I(N__38138));
    Span4Mux_h I__8341 (
            .O(N__38141),
            .I(N__38135));
    LocalMux I__8340 (
            .O(N__38138),
            .I(N__38132));
    Span4Mux_v I__8339 (
            .O(N__38135),
            .I(N__38129));
    Odrv4 I__8338 (
            .O(N__38132),
            .I(\ppm_encoder_1.un1_init_pulses_0_11 ));
    Odrv4 I__8337 (
            .O(N__38129),
            .I(\ppm_encoder_1.un1_init_pulses_0_11 ));
    InMux I__8336 (
            .O(N__38124),
            .I(N__38121));
    LocalMux I__8335 (
            .O(N__38121),
            .I(N__38118));
    Odrv4 I__8334 (
            .O(N__38118),
            .I(\ppm_encoder_1.un1_init_pulses_10_11 ));
    InMux I__8333 (
            .O(N__38115),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_10 ));
    InMux I__8332 (
            .O(N__38112),
            .I(N__38109));
    LocalMux I__8331 (
            .O(N__38109),
            .I(N__38106));
    Span4Mux_v I__8330 (
            .O(N__38106),
            .I(N__38103));
    Odrv4 I__8329 (
            .O(N__38103),
            .I(\ppm_encoder_1.elevator_RNIFQRT5Z0Z_12 ));
    CascadeMux I__8328 (
            .O(N__38100),
            .I(N__38097));
    InMux I__8327 (
            .O(N__38097),
            .I(N__38093));
    InMux I__8326 (
            .O(N__38096),
            .I(N__38090));
    LocalMux I__8325 (
            .O(N__38093),
            .I(N__38087));
    LocalMux I__8324 (
            .O(N__38090),
            .I(N__38084));
    Span12Mux_v I__8323 (
            .O(N__38087),
            .I(N__38081));
    Odrv12 I__8322 (
            .O(N__38084),
            .I(\ppm_encoder_1.un1_init_pulses_0_12 ));
    Odrv12 I__8321 (
            .O(N__38081),
            .I(\ppm_encoder_1.un1_init_pulses_0_12 ));
    InMux I__8320 (
            .O(N__38076),
            .I(N__38073));
    LocalMux I__8319 (
            .O(N__38073),
            .I(N__38070));
    Odrv4 I__8318 (
            .O(N__38070),
            .I(\ppm_encoder_1.un1_init_pulses_10_12 ));
    InMux I__8317 (
            .O(N__38067),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_11 ));
    InMux I__8316 (
            .O(N__38064),
            .I(N__38061));
    LocalMux I__8315 (
            .O(N__38061),
            .I(N__38058));
    Span4Mux_v I__8314 (
            .O(N__38058),
            .I(N__38055));
    Odrv4 I__8313 (
            .O(N__38055),
            .I(\ppm_encoder_1.elevator_RNIKVRT5Z0Z_13 ));
    CascadeMux I__8312 (
            .O(N__38052),
            .I(N__38049));
    InMux I__8311 (
            .O(N__38049),
            .I(N__38046));
    LocalMux I__8310 (
            .O(N__38046),
            .I(N__38042));
    InMux I__8309 (
            .O(N__38045),
            .I(N__38039));
    Span4Mux_h I__8308 (
            .O(N__38042),
            .I(N__38036));
    LocalMux I__8307 (
            .O(N__38039),
            .I(\ppm_encoder_1.un1_init_pulses_0_13 ));
    Odrv4 I__8306 (
            .O(N__38036),
            .I(\ppm_encoder_1.un1_init_pulses_0_13 ));
    InMux I__8305 (
            .O(N__38031),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_12 ));
    CascadeMux I__8304 (
            .O(N__38028),
            .I(N__38025));
    InMux I__8303 (
            .O(N__38025),
            .I(N__38022));
    LocalMux I__8302 (
            .O(N__38022),
            .I(\ppm_encoder_1.aileron_esr_RNITH3L6Z0Z_14 ));
    InMux I__8301 (
            .O(N__38019),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_13 ));
    InMux I__8300 (
            .O(N__38016),
            .I(N__38013));
    LocalMux I__8299 (
            .O(N__38013),
            .I(N__38010));
    Span4Mux_v I__8298 (
            .O(N__38010),
            .I(N__38007));
    Odrv4 I__8297 (
            .O(N__38007),
            .I(\ppm_encoder_1.throttle_RNIN3352Z0Z_0 ));
    CascadeMux I__8296 (
            .O(N__38004),
            .I(N__38001));
    InMux I__8295 (
            .O(N__38001),
            .I(N__37997));
    InMux I__8294 (
            .O(N__38000),
            .I(N__37994));
    LocalMux I__8293 (
            .O(N__37997),
            .I(N__37991));
    LocalMux I__8292 (
            .O(N__37994),
            .I(\ppm_encoder_1.un1_init_pulses_0 ));
    Odrv12 I__8291 (
            .O(N__37991),
            .I(\ppm_encoder_1.un1_init_pulses_0 ));
    InMux I__8290 (
            .O(N__37986),
            .I(N__37983));
    LocalMux I__8289 (
            .O(N__37983),
            .I(N__37980));
    Span4Mux_h I__8288 (
            .O(N__37980),
            .I(N__37977));
    Odrv4 I__8287 (
            .O(N__37977),
            .I(\ppm_encoder_1.throttle_RNIALN65Z0Z_1 ));
    CascadeMux I__8286 (
            .O(N__37974),
            .I(N__37970));
    InMux I__8285 (
            .O(N__37973),
            .I(N__37967));
    InMux I__8284 (
            .O(N__37970),
            .I(N__37964));
    LocalMux I__8283 (
            .O(N__37967),
            .I(N__37961));
    LocalMux I__8282 (
            .O(N__37964),
            .I(N__37958));
    Odrv4 I__8281 (
            .O(N__37961),
            .I(\ppm_encoder_1.un1_init_pulses_0_1 ));
    Odrv4 I__8280 (
            .O(N__37958),
            .I(\ppm_encoder_1.un1_init_pulses_0_1 ));
    CascadeMux I__8279 (
            .O(N__37953),
            .I(N__37950));
    InMux I__8278 (
            .O(N__37950),
            .I(N__37947));
    LocalMux I__8277 (
            .O(N__37947),
            .I(N__37944));
    Odrv4 I__8276 (
            .O(N__37944),
            .I(\ppm_encoder_1.un1_init_pulses_10_1 ));
    InMux I__8275 (
            .O(N__37941),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_0 ));
    InMux I__8274 (
            .O(N__37938),
            .I(N__37935));
    LocalMux I__8273 (
            .O(N__37935),
            .I(\ppm_encoder_1.throttle_RNI5V123Z0Z_2 ));
    CascadeMux I__8272 (
            .O(N__37932),
            .I(N__37929));
    InMux I__8271 (
            .O(N__37929),
            .I(N__37925));
    InMux I__8270 (
            .O(N__37928),
            .I(N__37922));
    LocalMux I__8269 (
            .O(N__37925),
            .I(\ppm_encoder_1.un1_init_pulses_0_2 ));
    LocalMux I__8268 (
            .O(N__37922),
            .I(\ppm_encoder_1.un1_init_pulses_0_2 ));
    InMux I__8267 (
            .O(N__37917),
            .I(N__37914));
    LocalMux I__8266 (
            .O(N__37914),
            .I(\ppm_encoder_1.un1_init_pulses_10_2 ));
    InMux I__8265 (
            .O(N__37911),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_1 ));
    InMux I__8264 (
            .O(N__37908),
            .I(N__37905));
    LocalMux I__8263 (
            .O(N__37905),
            .I(\ppm_encoder_1.throttle_RNI82223Z0Z_3 ));
    CascadeMux I__8262 (
            .O(N__37902),
            .I(N__37899));
    InMux I__8261 (
            .O(N__37899),
            .I(N__37895));
    InMux I__8260 (
            .O(N__37898),
            .I(N__37892));
    LocalMux I__8259 (
            .O(N__37895),
            .I(\ppm_encoder_1.un1_init_pulses_0_3 ));
    LocalMux I__8258 (
            .O(N__37892),
            .I(\ppm_encoder_1.un1_init_pulses_0_3 ));
    InMux I__8257 (
            .O(N__37887),
            .I(N__37884));
    LocalMux I__8256 (
            .O(N__37884),
            .I(\ppm_encoder_1.un1_init_pulses_10_3 ));
    InMux I__8255 (
            .O(N__37881),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_2 ));
    InMux I__8254 (
            .O(N__37878),
            .I(N__37875));
    LocalMux I__8253 (
            .O(N__37875),
            .I(N__37872));
    Odrv4 I__8252 (
            .O(N__37872),
            .I(\ppm_encoder_1.aileron_esr_RNIV9IN5Z0Z_4 ));
    CascadeMux I__8251 (
            .O(N__37869),
            .I(N__37866));
    InMux I__8250 (
            .O(N__37866),
            .I(N__37862));
    InMux I__8249 (
            .O(N__37865),
            .I(N__37859));
    LocalMux I__8248 (
            .O(N__37862),
            .I(N__37856));
    LocalMux I__8247 (
            .O(N__37859),
            .I(\ppm_encoder_1.un1_init_pulses_0_4 ));
    Odrv12 I__8246 (
            .O(N__37856),
            .I(\ppm_encoder_1.un1_init_pulses_0_4 ));
    InMux I__8245 (
            .O(N__37851),
            .I(N__37848));
    LocalMux I__8244 (
            .O(N__37848),
            .I(N__37845));
    Odrv4 I__8243 (
            .O(N__37845),
            .I(\ppm_encoder_1.un1_init_pulses_10_4 ));
    InMux I__8242 (
            .O(N__37842),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_3 ));
    InMux I__8241 (
            .O(N__37839),
            .I(N__37836));
    LocalMux I__8240 (
            .O(N__37836),
            .I(\ppm_encoder_1.aileron_esr_RNI4FIN5Z0Z_5 ));
    InMux I__8239 (
            .O(N__37833),
            .I(N__37829));
    CascadeMux I__8238 (
            .O(N__37832),
            .I(N__37826));
    LocalMux I__8237 (
            .O(N__37829),
            .I(N__37823));
    InMux I__8236 (
            .O(N__37826),
            .I(N__37820));
    Span4Mux_h I__8235 (
            .O(N__37823),
            .I(N__37817));
    LocalMux I__8234 (
            .O(N__37820),
            .I(N__37814));
    Odrv4 I__8233 (
            .O(N__37817),
            .I(\ppm_encoder_1.un1_init_pulses_0_5 ));
    Odrv12 I__8232 (
            .O(N__37814),
            .I(\ppm_encoder_1.un1_init_pulses_0_5 ));
    InMux I__8231 (
            .O(N__37809),
            .I(N__37806));
    LocalMux I__8230 (
            .O(N__37806),
            .I(N__37803));
    Odrv4 I__8229 (
            .O(N__37803),
            .I(\ppm_encoder_1.un1_init_pulses_10_5 ));
    InMux I__8228 (
            .O(N__37800),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_4 ));
    InMux I__8227 (
            .O(N__37797),
            .I(N__37794));
    LocalMux I__8226 (
            .O(N__37794),
            .I(N__37791));
    Odrv4 I__8225 (
            .O(N__37791),
            .I(\ppm_encoder_1.throttle_RNIEDI96Z0Z_6 ));
    CascadeMux I__8224 (
            .O(N__37788),
            .I(N__37784));
    InMux I__8223 (
            .O(N__37787),
            .I(N__37781));
    InMux I__8222 (
            .O(N__37784),
            .I(N__37778));
    LocalMux I__8221 (
            .O(N__37781),
            .I(\ppm_encoder_1.un1_init_pulses_0_6 ));
    LocalMux I__8220 (
            .O(N__37778),
            .I(\ppm_encoder_1.un1_init_pulses_0_6 ));
    InMux I__8219 (
            .O(N__37773),
            .I(N__37770));
    LocalMux I__8218 (
            .O(N__37770),
            .I(\ppm_encoder_1.un1_init_pulses_10_6 ));
    InMux I__8217 (
            .O(N__37767),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_5 ));
    InMux I__8216 (
            .O(N__37764),
            .I(N__37757));
    InMux I__8215 (
            .O(N__37763),
            .I(N__37757));
    InMux I__8214 (
            .O(N__37762),
            .I(N__37754));
    LocalMux I__8213 (
            .O(N__37757),
            .I(N__37751));
    LocalMux I__8212 (
            .O(N__37754),
            .I(N__37746));
    Sp12to4 I__8211 (
            .O(N__37751),
            .I(N__37746));
    Span12Mux_v I__8210 (
            .O(N__37746),
            .I(N__37743));
    Odrv12 I__8209 (
            .O(N__37743),
            .I(\ppm_encoder_1.init_pulsesZ0Z_11 ));
    InMux I__8208 (
            .O(N__37740),
            .I(N__37735));
    InMux I__8207 (
            .O(N__37739),
            .I(N__37730));
    InMux I__8206 (
            .O(N__37738),
            .I(N__37730));
    LocalMux I__8205 (
            .O(N__37735),
            .I(N__37725));
    LocalMux I__8204 (
            .O(N__37730),
            .I(N__37725));
    Span12Mux_v I__8203 (
            .O(N__37725),
            .I(N__37722));
    Odrv12 I__8202 (
            .O(N__37722),
            .I(\ppm_encoder_1.init_pulsesZ0Z_12 ));
    CascadeMux I__8201 (
            .O(N__37719),
            .I(N__37714));
    InMux I__8200 (
            .O(N__37718),
            .I(N__37705));
    InMux I__8199 (
            .O(N__37717),
            .I(N__37705));
    InMux I__8198 (
            .O(N__37714),
            .I(N__37705));
    InMux I__8197 (
            .O(N__37713),
            .I(N__37700));
    InMux I__8196 (
            .O(N__37712),
            .I(N__37697));
    LocalMux I__8195 (
            .O(N__37705),
            .I(N__37694));
    InMux I__8194 (
            .O(N__37704),
            .I(N__37691));
    CascadeMux I__8193 (
            .O(N__37703),
            .I(N__37688));
    LocalMux I__8192 (
            .O(N__37700),
            .I(N__37683));
    LocalMux I__8191 (
            .O(N__37697),
            .I(N__37680));
    Span4Mux_h I__8190 (
            .O(N__37694),
            .I(N__37675));
    LocalMux I__8189 (
            .O(N__37691),
            .I(N__37675));
    InMux I__8188 (
            .O(N__37688),
            .I(N__37670));
    InMux I__8187 (
            .O(N__37687),
            .I(N__37670));
    InMux I__8186 (
            .O(N__37686),
            .I(N__37667));
    Span12Mux_s10_h I__8185 (
            .O(N__37683),
            .I(N__37662));
    Sp12to4 I__8184 (
            .O(N__37680),
            .I(N__37662));
    Odrv4 I__8183 (
            .O(N__37675),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1Z0Z_0 ));
    LocalMux I__8182 (
            .O(N__37670),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1Z0Z_0 ));
    LocalMux I__8181 (
            .O(N__37667),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1Z0Z_0 ));
    Odrv12 I__8180 (
            .O(N__37662),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1Z0Z_0 ));
    InMux I__8179 (
            .O(N__37653),
            .I(N__37647));
    InMux I__8178 (
            .O(N__37652),
            .I(N__37642));
    InMux I__8177 (
            .O(N__37651),
            .I(N__37642));
    InMux I__8176 (
            .O(N__37650),
            .I(N__37639));
    LocalMux I__8175 (
            .O(N__37647),
            .I(\ppm_encoder_1.init_pulsesZ0Z_2 ));
    LocalMux I__8174 (
            .O(N__37642),
            .I(\ppm_encoder_1.init_pulsesZ0Z_2 ));
    LocalMux I__8173 (
            .O(N__37639),
            .I(\ppm_encoder_1.init_pulsesZ0Z_2 ));
    CascadeMux I__8172 (
            .O(N__37632),
            .I(N__37627));
    CascadeMux I__8171 (
            .O(N__37631),
            .I(N__37624));
    InMux I__8170 (
            .O(N__37630),
            .I(N__37621));
    InMux I__8169 (
            .O(N__37627),
            .I(N__37618));
    InMux I__8168 (
            .O(N__37624),
            .I(N__37615));
    LocalMux I__8167 (
            .O(N__37621),
            .I(N__37612));
    LocalMux I__8166 (
            .O(N__37618),
            .I(N__37609));
    LocalMux I__8165 (
            .O(N__37615),
            .I(N__37604));
    Span4Mux_v I__8164 (
            .O(N__37612),
            .I(N__37604));
    Span4Mux_h I__8163 (
            .O(N__37609),
            .I(N__37601));
    Odrv4 I__8162 (
            .O(N__37604),
            .I(\ppm_encoder_1.throttleZ0Z_2 ));
    Odrv4 I__8161 (
            .O(N__37601),
            .I(\ppm_encoder_1.throttleZ0Z_2 ));
    InMux I__8160 (
            .O(N__37596),
            .I(N__37593));
    LocalMux I__8159 (
            .O(N__37593),
            .I(N__37587));
    InMux I__8158 (
            .O(N__37592),
            .I(N__37584));
    InMux I__8157 (
            .O(N__37591),
            .I(N__37578));
    InMux I__8156 (
            .O(N__37590),
            .I(N__37575));
    Span4Mux_h I__8155 (
            .O(N__37587),
            .I(N__37569));
    LocalMux I__8154 (
            .O(N__37584),
            .I(N__37569));
    InMux I__8153 (
            .O(N__37583),
            .I(N__37565));
    InMux I__8152 (
            .O(N__37582),
            .I(N__37562));
    InMux I__8151 (
            .O(N__37581),
            .I(N__37559));
    LocalMux I__8150 (
            .O(N__37578),
            .I(N__37554));
    LocalMux I__8149 (
            .O(N__37575),
            .I(N__37554));
    InMux I__8148 (
            .O(N__37574),
            .I(N__37545));
    Span4Mux_v I__8147 (
            .O(N__37569),
            .I(N__37542));
    InMux I__8146 (
            .O(N__37568),
            .I(N__37539));
    LocalMux I__8145 (
            .O(N__37565),
            .I(N__37530));
    LocalMux I__8144 (
            .O(N__37562),
            .I(N__37530));
    LocalMux I__8143 (
            .O(N__37559),
            .I(N__37530));
    Span4Mux_v I__8142 (
            .O(N__37554),
            .I(N__37530));
    InMux I__8141 (
            .O(N__37553),
            .I(N__37525));
    InMux I__8140 (
            .O(N__37552),
            .I(N__37525));
    InMux I__8139 (
            .O(N__37551),
            .I(N__37518));
    InMux I__8138 (
            .O(N__37550),
            .I(N__37518));
    InMux I__8137 (
            .O(N__37549),
            .I(N__37518));
    InMux I__8136 (
            .O(N__37548),
            .I(N__37515));
    LocalMux I__8135 (
            .O(N__37545),
            .I(N__37512));
    Odrv4 I__8134 (
            .O(N__37542),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_0 ));
    LocalMux I__8133 (
            .O(N__37539),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_0 ));
    Odrv4 I__8132 (
            .O(N__37530),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_0 ));
    LocalMux I__8131 (
            .O(N__37525),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_0 ));
    LocalMux I__8130 (
            .O(N__37518),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_0 ));
    LocalMux I__8129 (
            .O(N__37515),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_0 ));
    Odrv4 I__8128 (
            .O(N__37512),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_0 ));
    CascadeMux I__8127 (
            .O(N__37497),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_2_cascade_ ));
    InMux I__8126 (
            .O(N__37494),
            .I(N__37491));
    LocalMux I__8125 (
            .O(N__37491),
            .I(N__37488));
    Span4Mux_v I__8124 (
            .O(N__37488),
            .I(N__37483));
    InMux I__8123 (
            .O(N__37487),
            .I(N__37480));
    InMux I__8122 (
            .O(N__37486),
            .I(N__37477));
    Odrv4 I__8121 (
            .O(N__37483),
            .I(\ppm_encoder_1.init_pulsesZ0Z_6 ));
    LocalMux I__8120 (
            .O(N__37480),
            .I(\ppm_encoder_1.init_pulsesZ0Z_6 ));
    LocalMux I__8119 (
            .O(N__37477),
            .I(\ppm_encoder_1.init_pulsesZ0Z_6 ));
    InMux I__8118 (
            .O(N__37470),
            .I(N__37461));
    InMux I__8117 (
            .O(N__37469),
            .I(N__37461));
    InMux I__8116 (
            .O(N__37468),
            .I(N__37461));
    LocalMux I__8115 (
            .O(N__37461),
            .I(\ppm_encoder_1.init_pulsesZ0Z_4 ));
    InMux I__8114 (
            .O(N__37458),
            .I(N__37455));
    LocalMux I__8113 (
            .O(N__37455),
            .I(N__37451));
    InMux I__8112 (
            .O(N__37454),
            .I(N__37448));
    Span4Mux_v I__8111 (
            .O(N__37451),
            .I(N__37443));
    LocalMux I__8110 (
            .O(N__37448),
            .I(N__37443));
    Odrv4 I__8109 (
            .O(N__37443),
            .I(\ppm_encoder_1.rudderZ0Z_4 ));
    InMux I__8108 (
            .O(N__37440),
            .I(N__37437));
    LocalMux I__8107 (
            .O(N__37437),
            .I(N__37434));
    Span4Mux_v I__8106 (
            .O(N__37434),
            .I(N__37431));
    Odrv4 I__8105 (
            .O(N__37431),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_4 ));
    InMux I__8104 (
            .O(N__37428),
            .I(N__37419));
    InMux I__8103 (
            .O(N__37427),
            .I(N__37419));
    InMux I__8102 (
            .O(N__37426),
            .I(N__37419));
    LocalMux I__8101 (
            .O(N__37419),
            .I(\ppm_encoder_1.init_pulsesZ0Z_5 ));
    InMux I__8100 (
            .O(N__37416),
            .I(N__37413));
    LocalMux I__8099 (
            .O(N__37413),
            .I(N__37409));
    InMux I__8098 (
            .O(N__37412),
            .I(N__37406));
    Span4Mux_v I__8097 (
            .O(N__37409),
            .I(N__37401));
    LocalMux I__8096 (
            .O(N__37406),
            .I(N__37401));
    Odrv4 I__8095 (
            .O(N__37401),
            .I(\ppm_encoder_1.rudderZ0Z_5 ));
    InMux I__8094 (
            .O(N__37398),
            .I(N__37395));
    LocalMux I__8093 (
            .O(N__37395),
            .I(N__37392));
    Span4Mux_v I__8092 (
            .O(N__37392),
            .I(N__37389));
    Odrv4 I__8091 (
            .O(N__37389),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_5 ));
    InMux I__8090 (
            .O(N__37386),
            .I(N__37381));
    InMux I__8089 (
            .O(N__37385),
            .I(N__37376));
    InMux I__8088 (
            .O(N__37384),
            .I(N__37376));
    LocalMux I__8087 (
            .O(N__37381),
            .I(\ppm_encoder_1.init_pulsesZ0Z_1 ));
    LocalMux I__8086 (
            .O(N__37376),
            .I(\ppm_encoder_1.init_pulsesZ0Z_1 ));
    InMux I__8085 (
            .O(N__37371),
            .I(N__37367));
    InMux I__8084 (
            .O(N__37370),
            .I(N__37364));
    LocalMux I__8083 (
            .O(N__37367),
            .I(\reset_module_System.countZ0Z_11 ));
    LocalMux I__8082 (
            .O(N__37364),
            .I(\reset_module_System.countZ0Z_11 ));
    InMux I__8081 (
            .O(N__37359),
            .I(N__37355));
    InMux I__8080 (
            .O(N__37358),
            .I(N__37352));
    LocalMux I__8079 (
            .O(N__37355),
            .I(\reset_module_System.countZ0Z_14 ));
    LocalMux I__8078 (
            .O(N__37352),
            .I(\reset_module_System.countZ0Z_14 ));
    CascadeMux I__8077 (
            .O(N__37347),
            .I(N__37344));
    InMux I__8076 (
            .O(N__37344),
            .I(N__37340));
    InMux I__8075 (
            .O(N__37343),
            .I(N__37337));
    LocalMux I__8074 (
            .O(N__37340),
            .I(\reset_module_System.countZ0Z_17 ));
    LocalMux I__8073 (
            .O(N__37337),
            .I(\reset_module_System.countZ0Z_17 ));
    InMux I__8072 (
            .O(N__37332),
            .I(N__37328));
    InMux I__8071 (
            .O(N__37331),
            .I(N__37325));
    LocalMux I__8070 (
            .O(N__37328),
            .I(\reset_module_System.countZ0Z_10 ));
    LocalMux I__8069 (
            .O(N__37325),
            .I(\reset_module_System.countZ0Z_10 ));
    InMux I__8068 (
            .O(N__37320),
            .I(N__37314));
    InMux I__8067 (
            .O(N__37319),
            .I(N__37311));
    InMux I__8066 (
            .O(N__37318),
            .I(N__37308));
    InMux I__8065 (
            .O(N__37317),
            .I(N__37305));
    LocalMux I__8064 (
            .O(N__37314),
            .I(N__37302));
    LocalMux I__8063 (
            .O(N__37311),
            .I(N__37299));
    LocalMux I__8062 (
            .O(N__37308),
            .I(N__37294));
    LocalMux I__8061 (
            .O(N__37305),
            .I(N__37294));
    Span4Mux_h I__8060 (
            .O(N__37302),
            .I(N__37291));
    Span4Mux_h I__8059 (
            .O(N__37299),
            .I(N__37288));
    Span4Mux_h I__8058 (
            .O(N__37294),
            .I(N__37285));
    Span4Mux_h I__8057 (
            .O(N__37291),
            .I(N__37282));
    Odrv4 I__8056 (
            .O(N__37288),
            .I(\reset_module_System.reset6_14 ));
    Odrv4 I__8055 (
            .O(N__37285),
            .I(\reset_module_System.reset6_14 ));
    Odrv4 I__8054 (
            .O(N__37282),
            .I(\reset_module_System.reset6_14 ));
    InMux I__8053 (
            .O(N__37275),
            .I(N__37272));
    LocalMux I__8052 (
            .O(N__37272),
            .I(\ppm_encoder_1.un1_init_pulses_10_0 ));
    CascadeMux I__8051 (
            .O(N__37269),
            .I(\ppm_encoder_1.un1_init_pulses_11_0_cascade_ ));
    CascadeMux I__8050 (
            .O(N__37266),
            .I(\ppm_encoder_1.un1_init_pulses_0_cascade_ ));
    CascadeMux I__8049 (
            .O(N__37263),
            .I(N__37251));
    CascadeMux I__8048 (
            .O(N__37262),
            .I(N__37247));
    CascadeMux I__8047 (
            .O(N__37261),
            .I(N__37244));
    CascadeMux I__8046 (
            .O(N__37260),
            .I(N__37237));
    CascadeMux I__8045 (
            .O(N__37259),
            .I(N__37234));
    CascadeMux I__8044 (
            .O(N__37258),
            .I(N__37228));
    CascadeMux I__8043 (
            .O(N__37257),
            .I(N__37221));
    CascadeMux I__8042 (
            .O(N__37256),
            .I(N__37218));
    CascadeMux I__8041 (
            .O(N__37255),
            .I(N__37215));
    InMux I__8040 (
            .O(N__37254),
            .I(N__37207));
    InMux I__8039 (
            .O(N__37251),
            .I(N__37207));
    InMux I__8038 (
            .O(N__37250),
            .I(N__37207));
    InMux I__8037 (
            .O(N__37247),
            .I(N__37204));
    InMux I__8036 (
            .O(N__37244),
            .I(N__37200));
    CascadeMux I__8035 (
            .O(N__37243),
            .I(N__37197));
    CascadeMux I__8034 (
            .O(N__37242),
            .I(N__37194));
    CascadeMux I__8033 (
            .O(N__37241),
            .I(N__37188));
    InMux I__8032 (
            .O(N__37240),
            .I(N__37181));
    InMux I__8031 (
            .O(N__37237),
            .I(N__37181));
    InMux I__8030 (
            .O(N__37234),
            .I(N__37181));
    InMux I__8029 (
            .O(N__37233),
            .I(N__37172));
    InMux I__8028 (
            .O(N__37232),
            .I(N__37172));
    InMux I__8027 (
            .O(N__37231),
            .I(N__37172));
    InMux I__8026 (
            .O(N__37228),
            .I(N__37172));
    CascadeMux I__8025 (
            .O(N__37227),
            .I(N__37169));
    CascadeMux I__8024 (
            .O(N__37226),
            .I(N__37166));
    InMux I__8023 (
            .O(N__37225),
            .I(N__37158));
    InMux I__8022 (
            .O(N__37224),
            .I(N__37158));
    InMux I__8021 (
            .O(N__37221),
            .I(N__37158));
    InMux I__8020 (
            .O(N__37218),
            .I(N__37151));
    InMux I__8019 (
            .O(N__37215),
            .I(N__37151));
    InMux I__8018 (
            .O(N__37214),
            .I(N__37151));
    LocalMux I__8017 (
            .O(N__37207),
            .I(N__37142));
    LocalMux I__8016 (
            .O(N__37204),
            .I(N__37142));
    InMux I__8015 (
            .O(N__37203),
            .I(N__37139));
    LocalMux I__8014 (
            .O(N__37200),
            .I(N__37136));
    InMux I__8013 (
            .O(N__37197),
            .I(N__37129));
    InMux I__8012 (
            .O(N__37194),
            .I(N__37129));
    InMux I__8011 (
            .O(N__37193),
            .I(N__37129));
    InMux I__8010 (
            .O(N__37192),
            .I(N__37122));
    InMux I__8009 (
            .O(N__37191),
            .I(N__37122));
    InMux I__8008 (
            .O(N__37188),
            .I(N__37122));
    LocalMux I__8007 (
            .O(N__37181),
            .I(N__37117));
    LocalMux I__8006 (
            .O(N__37172),
            .I(N__37117));
    InMux I__8005 (
            .O(N__37169),
            .I(N__37110));
    InMux I__8004 (
            .O(N__37166),
            .I(N__37110));
    InMux I__8003 (
            .O(N__37165),
            .I(N__37110));
    LocalMux I__8002 (
            .O(N__37158),
            .I(N__37105));
    LocalMux I__8001 (
            .O(N__37151),
            .I(N__37105));
    CascadeMux I__8000 (
            .O(N__37150),
            .I(N__37099));
    CascadeMux I__7999 (
            .O(N__37149),
            .I(N__37096));
    CascadeMux I__7998 (
            .O(N__37148),
            .I(N__37093));
    CascadeMux I__7997 (
            .O(N__37147),
            .I(N__37086));
    Span4Mux_v I__7996 (
            .O(N__37142),
            .I(N__37083));
    LocalMux I__7995 (
            .O(N__37139),
            .I(N__37080));
    Span4Mux_v I__7994 (
            .O(N__37136),
            .I(N__37071));
    LocalMux I__7993 (
            .O(N__37129),
            .I(N__37071));
    LocalMux I__7992 (
            .O(N__37122),
            .I(N__37071));
    Span4Mux_v I__7991 (
            .O(N__37117),
            .I(N__37071));
    LocalMux I__7990 (
            .O(N__37110),
            .I(N__37068));
    Span4Mux_v I__7989 (
            .O(N__37105),
            .I(N__37065));
    InMux I__7988 (
            .O(N__37104),
            .I(N__37054));
    InMux I__7987 (
            .O(N__37103),
            .I(N__37054));
    InMux I__7986 (
            .O(N__37102),
            .I(N__37054));
    InMux I__7985 (
            .O(N__37099),
            .I(N__37054));
    InMux I__7984 (
            .O(N__37096),
            .I(N__37054));
    InMux I__7983 (
            .O(N__37093),
            .I(N__37047));
    InMux I__7982 (
            .O(N__37092),
            .I(N__37047));
    InMux I__7981 (
            .O(N__37091),
            .I(N__37047));
    InMux I__7980 (
            .O(N__37090),
            .I(N__37040));
    InMux I__7979 (
            .O(N__37089),
            .I(N__37040));
    InMux I__7978 (
            .O(N__37086),
            .I(N__37040));
    Span4Mux_h I__7977 (
            .O(N__37083),
            .I(N__37037));
    Span4Mux_v I__7976 (
            .O(N__37080),
            .I(N__37032));
    Span4Mux_v I__7975 (
            .O(N__37071),
            .I(N__37032));
    Sp12to4 I__7974 (
            .O(N__37068),
            .I(N__37029));
    Span4Mux_h I__7973 (
            .O(N__37065),
            .I(N__37026));
    LocalMux I__7972 (
            .O(N__37054),
            .I(N__37021));
    LocalMux I__7971 (
            .O(N__37047),
            .I(N__37021));
    LocalMux I__7970 (
            .O(N__37040),
            .I(N__37012));
    Sp12to4 I__7969 (
            .O(N__37037),
            .I(N__37012));
    Sp12to4 I__7968 (
            .O(N__37032),
            .I(N__37012));
    Span12Mux_v I__7967 (
            .O(N__37029),
            .I(N__37012));
    Span4Mux_h I__7966 (
            .O(N__37026),
            .I(N__37009));
    Span12Mux_v I__7965 (
            .O(N__37021),
            .I(N__37006));
    Span12Mux_h I__7964 (
            .O(N__37012),
            .I(N__37003));
    Odrv4 I__7963 (
            .O(N__37009),
            .I(pid_altitude_dv));
    Odrv12 I__7962 (
            .O(N__37006),
            .I(pid_altitude_dv));
    Odrv12 I__7961 (
            .O(N__37003),
            .I(pid_altitude_dv));
    InMux I__7960 (
            .O(N__36996),
            .I(N__36993));
    LocalMux I__7959 (
            .O(N__36993),
            .I(N__36989));
    CascadeMux I__7958 (
            .O(N__36992),
            .I(N__36985));
    Span4Mux_v I__7957 (
            .O(N__36989),
            .I(N__36982));
    InMux I__7956 (
            .O(N__36988),
            .I(N__36979));
    InMux I__7955 (
            .O(N__36985),
            .I(N__36976));
    Span4Mux_h I__7954 (
            .O(N__36982),
            .I(N__36971));
    LocalMux I__7953 (
            .O(N__36979),
            .I(N__36971));
    LocalMux I__7952 (
            .O(N__36976),
            .I(throttle_command_0));
    Odrv4 I__7951 (
            .O(N__36971),
            .I(throttle_command_0));
    InMux I__7950 (
            .O(N__36966),
            .I(N__36960));
    InMux I__7949 (
            .O(N__36965),
            .I(N__36957));
    InMux I__7948 (
            .O(N__36964),
            .I(N__36952));
    InMux I__7947 (
            .O(N__36963),
            .I(N__36952));
    LocalMux I__7946 (
            .O(N__36960),
            .I(\ppm_encoder_1.throttleZ0Z_0 ));
    LocalMux I__7945 (
            .O(N__36957),
            .I(\ppm_encoder_1.throttleZ0Z_0 ));
    LocalMux I__7944 (
            .O(N__36952),
            .I(\ppm_encoder_1.throttleZ0Z_0 ));
    CascadeMux I__7943 (
            .O(N__36945),
            .I(N__36942));
    InMux I__7942 (
            .O(N__36942),
            .I(N__36936));
    InMux I__7941 (
            .O(N__36941),
            .I(N__36933));
    InMux I__7940 (
            .O(N__36940),
            .I(N__36928));
    InMux I__7939 (
            .O(N__36939),
            .I(N__36928));
    LocalMux I__7938 (
            .O(N__36936),
            .I(\ppm_encoder_1.init_pulsesZ0Z_0 ));
    LocalMux I__7937 (
            .O(N__36933),
            .I(\ppm_encoder_1.init_pulsesZ0Z_0 ));
    LocalMux I__7936 (
            .O(N__36928),
            .I(\ppm_encoder_1.init_pulsesZ0Z_0 ));
    InMux I__7935 (
            .O(N__36921),
            .I(N__36918));
    LocalMux I__7934 (
            .O(N__36918),
            .I(N__36915));
    Span4Mux_v I__7933 (
            .O(N__36915),
            .I(N__36912));
    Span4Mux_v I__7932 (
            .O(N__36912),
            .I(N__36909));
    Odrv4 I__7931 (
            .O(N__36909),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_0 ));
    InMux I__7930 (
            .O(N__36906),
            .I(\ppm_encoder_1.un1_counter_13_cry_17 ));
    SRMux I__7929 (
            .O(N__36903),
            .I(N__36894));
    SRMux I__7928 (
            .O(N__36902),
            .I(N__36894));
    SRMux I__7927 (
            .O(N__36901),
            .I(N__36894));
    GlobalMux I__7926 (
            .O(N__36894),
            .I(N__36891));
    gio2CtrlBuf I__7925 (
            .O(N__36891),
            .I(\ppm_encoder_1.N_322_g ));
    InMux I__7924 (
            .O(N__36888),
            .I(N__36884));
    InMux I__7923 (
            .O(N__36887),
            .I(N__36881));
    LocalMux I__7922 (
            .O(N__36884),
            .I(N__36877));
    LocalMux I__7921 (
            .O(N__36881),
            .I(N__36874));
    InMux I__7920 (
            .O(N__36880),
            .I(N__36868));
    Span4Mux_h I__7919 (
            .O(N__36877),
            .I(N__36861));
    Span4Mux_v I__7918 (
            .O(N__36874),
            .I(N__36858));
    InMux I__7917 (
            .O(N__36873),
            .I(N__36852));
    InMux I__7916 (
            .O(N__36872),
            .I(N__36849));
    InMux I__7915 (
            .O(N__36871),
            .I(N__36846));
    LocalMux I__7914 (
            .O(N__36868),
            .I(N__36843));
    CascadeMux I__7913 (
            .O(N__36867),
            .I(N__36840));
    CascadeMux I__7912 (
            .O(N__36866),
            .I(N__36835));
    InMux I__7911 (
            .O(N__36865),
            .I(N__36832));
    InMux I__7910 (
            .O(N__36864),
            .I(N__36829));
    Sp12to4 I__7909 (
            .O(N__36861),
            .I(N__36826));
    Sp12to4 I__7908 (
            .O(N__36858),
            .I(N__36823));
    InMux I__7907 (
            .O(N__36857),
            .I(N__36820));
    InMux I__7906 (
            .O(N__36856),
            .I(N__36816));
    InMux I__7905 (
            .O(N__36855),
            .I(N__36813));
    LocalMux I__7904 (
            .O(N__36852),
            .I(N__36810));
    LocalMux I__7903 (
            .O(N__36849),
            .I(N__36807));
    LocalMux I__7902 (
            .O(N__36846),
            .I(N__36802));
    Span12Mux_s10_v I__7901 (
            .O(N__36843),
            .I(N__36802));
    InMux I__7900 (
            .O(N__36840),
            .I(N__36799));
    InMux I__7899 (
            .O(N__36839),
            .I(N__36792));
    InMux I__7898 (
            .O(N__36838),
            .I(N__36792));
    InMux I__7897 (
            .O(N__36835),
            .I(N__36792));
    LocalMux I__7896 (
            .O(N__36832),
            .I(N__36781));
    LocalMux I__7895 (
            .O(N__36829),
            .I(N__36781));
    Span12Mux_s10_v I__7894 (
            .O(N__36826),
            .I(N__36781));
    Span12Mux_h I__7893 (
            .O(N__36823),
            .I(N__36781));
    LocalMux I__7892 (
            .O(N__36820),
            .I(N__36781));
    InMux I__7891 (
            .O(N__36819),
            .I(N__36778));
    LocalMux I__7890 (
            .O(N__36816),
            .I(N__36769));
    LocalMux I__7889 (
            .O(N__36813),
            .I(N__36769));
    Span4Mux_v I__7888 (
            .O(N__36810),
            .I(N__36769));
    Span4Mux_v I__7887 (
            .O(N__36807),
            .I(N__36769));
    Span12Mux_v I__7886 (
            .O(N__36802),
            .I(N__36766));
    LocalMux I__7885 (
            .O(N__36799),
            .I(N__36759));
    LocalMux I__7884 (
            .O(N__36792),
            .I(N__36759));
    Span12Mux_v I__7883 (
            .O(N__36781),
            .I(N__36759));
    LocalMux I__7882 (
            .O(N__36778),
            .I(uart_pc_data_2));
    Odrv4 I__7881 (
            .O(N__36769),
            .I(uart_pc_data_2));
    Odrv12 I__7880 (
            .O(N__36766),
            .I(uart_pc_data_2));
    Odrv12 I__7879 (
            .O(N__36759),
            .I(uart_pc_data_2));
    InMux I__7878 (
            .O(N__36750),
            .I(N__36747));
    LocalMux I__7877 (
            .O(N__36747),
            .I(N__36744));
    Span12Mux_s9_h I__7876 (
            .O(N__36744),
            .I(N__36741));
    Odrv12 I__7875 (
            .O(N__36741),
            .I(alt_ki_2));
    InMux I__7874 (
            .O(N__36738),
            .I(N__36735));
    LocalMux I__7873 (
            .O(N__36735),
            .I(N__36732));
    Odrv12 I__7872 (
            .O(N__36732),
            .I(\pid_alt.O_0_6 ));
    CascadeMux I__7871 (
            .O(N__36729),
            .I(N__36726));
    InMux I__7870 (
            .O(N__36726),
            .I(N__36723));
    LocalMux I__7869 (
            .O(N__36723),
            .I(N__36720));
    Span4Mux_h I__7868 (
            .O(N__36720),
            .I(N__36717));
    Odrv4 I__7867 (
            .O(N__36717),
            .I(\pid_alt.error_i_regZ0Z_2 ));
    CascadeMux I__7866 (
            .O(N__36714),
            .I(N__36711));
    InMux I__7865 (
            .O(N__36711),
            .I(N__36707));
    InMux I__7864 (
            .O(N__36710),
            .I(N__36704));
    LocalMux I__7863 (
            .O(N__36707),
            .I(N__36699));
    LocalMux I__7862 (
            .O(N__36704),
            .I(N__36699));
    Span4Mux_v I__7861 (
            .O(N__36699),
            .I(N__36696));
    Odrv4 I__7860 (
            .O(N__36696),
            .I(\uart_drone.N_144_1 ));
    CascadeMux I__7859 (
            .O(N__36693),
            .I(N__36688));
    InMux I__7858 (
            .O(N__36692),
            .I(N__36683));
    InMux I__7857 (
            .O(N__36691),
            .I(N__36680));
    InMux I__7856 (
            .O(N__36688),
            .I(N__36672));
    InMux I__7855 (
            .O(N__36687),
            .I(N__36672));
    CascadeMux I__7854 (
            .O(N__36686),
            .I(N__36668));
    LocalMux I__7853 (
            .O(N__36683),
            .I(N__36663));
    LocalMux I__7852 (
            .O(N__36680),
            .I(N__36663));
    InMux I__7851 (
            .O(N__36679),
            .I(N__36660));
    InMux I__7850 (
            .O(N__36678),
            .I(N__36655));
    InMux I__7849 (
            .O(N__36677),
            .I(N__36655));
    LocalMux I__7848 (
            .O(N__36672),
            .I(N__36652));
    InMux I__7847 (
            .O(N__36671),
            .I(N__36649));
    InMux I__7846 (
            .O(N__36668),
            .I(N__36646));
    Span4Mux_v I__7845 (
            .O(N__36663),
            .I(N__36641));
    LocalMux I__7844 (
            .O(N__36660),
            .I(N__36641));
    LocalMux I__7843 (
            .O(N__36655),
            .I(N__36638));
    Span4Mux_h I__7842 (
            .O(N__36652),
            .I(N__36633));
    LocalMux I__7841 (
            .O(N__36649),
            .I(N__36633));
    LocalMux I__7840 (
            .O(N__36646),
            .I(N__36626));
    Span4Mux_h I__7839 (
            .O(N__36641),
            .I(N__36626));
    Span4Mux_v I__7838 (
            .O(N__36638),
            .I(N__36626));
    Span4Mux_h I__7837 (
            .O(N__36633),
            .I(N__36623));
    Odrv4 I__7836 (
            .O(N__36626),
            .I(\uart_drone.bit_CountZ0Z_2 ));
    Odrv4 I__7835 (
            .O(N__36623),
            .I(\uart_drone.bit_CountZ0Z_2 ));
    InMux I__7834 (
            .O(N__36618),
            .I(N__36612));
    InMux I__7833 (
            .O(N__36617),
            .I(N__36609));
    InMux I__7832 (
            .O(N__36616),
            .I(N__36601));
    InMux I__7831 (
            .O(N__36615),
            .I(N__36598));
    LocalMux I__7830 (
            .O(N__36612),
            .I(N__36595));
    LocalMux I__7829 (
            .O(N__36609),
            .I(N__36592));
    CascadeMux I__7828 (
            .O(N__36608),
            .I(N__36589));
    InMux I__7827 (
            .O(N__36607),
            .I(N__36586));
    InMux I__7826 (
            .O(N__36606),
            .I(N__36583));
    InMux I__7825 (
            .O(N__36605),
            .I(N__36580));
    InMux I__7824 (
            .O(N__36604),
            .I(N__36577));
    LocalMux I__7823 (
            .O(N__36601),
            .I(N__36572));
    LocalMux I__7822 (
            .O(N__36598),
            .I(N__36572));
    Span4Mux_v I__7821 (
            .O(N__36595),
            .I(N__36567));
    Span4Mux_v I__7820 (
            .O(N__36592),
            .I(N__36567));
    InMux I__7819 (
            .O(N__36589),
            .I(N__36564));
    LocalMux I__7818 (
            .O(N__36586),
            .I(\uart_drone.timer_CountZ0Z_4 ));
    LocalMux I__7817 (
            .O(N__36583),
            .I(\uart_drone.timer_CountZ0Z_4 ));
    LocalMux I__7816 (
            .O(N__36580),
            .I(\uart_drone.timer_CountZ0Z_4 ));
    LocalMux I__7815 (
            .O(N__36577),
            .I(\uart_drone.timer_CountZ0Z_4 ));
    Odrv4 I__7814 (
            .O(N__36572),
            .I(\uart_drone.timer_CountZ0Z_4 ));
    Odrv4 I__7813 (
            .O(N__36567),
            .I(\uart_drone.timer_CountZ0Z_4 ));
    LocalMux I__7812 (
            .O(N__36564),
            .I(\uart_drone.timer_CountZ0Z_4 ));
    InMux I__7811 (
            .O(N__36549),
            .I(N__36546));
    LocalMux I__7810 (
            .O(N__36546),
            .I(N__36541));
    InMux I__7809 (
            .O(N__36545),
            .I(N__36538));
    InMux I__7808 (
            .O(N__36544),
            .I(N__36532));
    Span4Mux_v I__7807 (
            .O(N__36541),
            .I(N__36526));
    LocalMux I__7806 (
            .O(N__36538),
            .I(N__36526));
    InMux I__7805 (
            .O(N__36537),
            .I(N__36522));
    InMux I__7804 (
            .O(N__36536),
            .I(N__36519));
    InMux I__7803 (
            .O(N__36535),
            .I(N__36516));
    LocalMux I__7802 (
            .O(N__36532),
            .I(N__36513));
    InMux I__7801 (
            .O(N__36531),
            .I(N__36510));
    Span4Mux_h I__7800 (
            .O(N__36526),
            .I(N__36507));
    InMux I__7799 (
            .O(N__36525),
            .I(N__36504));
    LocalMux I__7798 (
            .O(N__36522),
            .I(\uart_drone.timer_CountZ1Z_3 ));
    LocalMux I__7797 (
            .O(N__36519),
            .I(\uart_drone.timer_CountZ1Z_3 ));
    LocalMux I__7796 (
            .O(N__36516),
            .I(\uart_drone.timer_CountZ1Z_3 ));
    Odrv4 I__7795 (
            .O(N__36513),
            .I(\uart_drone.timer_CountZ1Z_3 ));
    LocalMux I__7794 (
            .O(N__36510),
            .I(\uart_drone.timer_CountZ1Z_3 ));
    Odrv4 I__7793 (
            .O(N__36507),
            .I(\uart_drone.timer_CountZ1Z_3 ));
    LocalMux I__7792 (
            .O(N__36504),
            .I(\uart_drone.timer_CountZ1Z_3 ));
    InMux I__7791 (
            .O(N__36489),
            .I(N__36485));
    InMux I__7790 (
            .O(N__36488),
            .I(N__36480));
    LocalMux I__7789 (
            .O(N__36485),
            .I(N__36477));
    InMux I__7788 (
            .O(N__36484),
            .I(N__36472));
    InMux I__7787 (
            .O(N__36483),
            .I(N__36469));
    LocalMux I__7786 (
            .O(N__36480),
            .I(N__36464));
    Span4Mux_h I__7785 (
            .O(N__36477),
            .I(N__36464));
    InMux I__7784 (
            .O(N__36476),
            .I(N__36459));
    InMux I__7783 (
            .O(N__36475),
            .I(N__36459));
    LocalMux I__7782 (
            .O(N__36472),
            .I(\uart_drone.stateZ0Z_4 ));
    LocalMux I__7781 (
            .O(N__36469),
            .I(\uart_drone.stateZ0Z_4 ));
    Odrv4 I__7780 (
            .O(N__36464),
            .I(\uart_drone.stateZ0Z_4 ));
    LocalMux I__7779 (
            .O(N__36459),
            .I(\uart_drone.stateZ0Z_4 ));
    CascadeMux I__7778 (
            .O(N__36450),
            .I(\uart_drone.un1_state_4_0_cascade_ ));
    InMux I__7777 (
            .O(N__36447),
            .I(bfn_16_20_0_));
    InMux I__7776 (
            .O(N__36444),
            .I(\ppm_encoder_1.un1_counter_13_cry_8 ));
    InMux I__7775 (
            .O(N__36441),
            .I(\ppm_encoder_1.un1_counter_13_cry_9 ));
    InMux I__7774 (
            .O(N__36438),
            .I(\ppm_encoder_1.un1_counter_13_cry_10 ));
    InMux I__7773 (
            .O(N__36435),
            .I(\ppm_encoder_1.un1_counter_13_cry_11 ));
    InMux I__7772 (
            .O(N__36432),
            .I(\ppm_encoder_1.un1_counter_13_cry_12 ));
    InMux I__7771 (
            .O(N__36429),
            .I(\ppm_encoder_1.un1_counter_13_cry_13 ));
    InMux I__7770 (
            .O(N__36426),
            .I(\ppm_encoder_1.un1_counter_13_cry_14 ));
    InMux I__7769 (
            .O(N__36423),
            .I(bfn_16_21_0_));
    InMux I__7768 (
            .O(N__36420),
            .I(\ppm_encoder_1.un1_counter_13_cry_16 ));
    CascadeMux I__7767 (
            .O(N__36417),
            .I(N__36413));
    InMux I__7766 (
            .O(N__36416),
            .I(N__36410));
    InMux I__7765 (
            .O(N__36413),
            .I(N__36407));
    LocalMux I__7764 (
            .O(N__36410),
            .I(N__36404));
    LocalMux I__7763 (
            .O(N__36407),
            .I(N__36401));
    Span4Mux_v I__7762 (
            .O(N__36404),
            .I(N__36396));
    Span4Mux_v I__7761 (
            .O(N__36401),
            .I(N__36396));
    Odrv4 I__7760 (
            .O(N__36396),
            .I(\ppm_encoder_1.N_1330_i ));
    CascadeMux I__7759 (
            .O(N__36393),
            .I(N__36388));
    InMux I__7758 (
            .O(N__36392),
            .I(N__36385));
    InMux I__7757 (
            .O(N__36391),
            .I(N__36382));
    InMux I__7756 (
            .O(N__36388),
            .I(N__36379));
    LocalMux I__7755 (
            .O(N__36385),
            .I(\ppm_encoder_1.counterZ0Z_0 ));
    LocalMux I__7754 (
            .O(N__36382),
            .I(\ppm_encoder_1.counterZ0Z_0 ));
    LocalMux I__7753 (
            .O(N__36379),
            .I(\ppm_encoder_1.counterZ0Z_0 ));
    InMux I__7752 (
            .O(N__36372),
            .I(N__36366));
    InMux I__7751 (
            .O(N__36371),
            .I(N__36361));
    InMux I__7750 (
            .O(N__36370),
            .I(N__36361));
    InMux I__7749 (
            .O(N__36369),
            .I(N__36358));
    LocalMux I__7748 (
            .O(N__36366),
            .I(\ppm_encoder_1.counterZ0Z_1 ));
    LocalMux I__7747 (
            .O(N__36361),
            .I(\ppm_encoder_1.counterZ0Z_1 ));
    LocalMux I__7746 (
            .O(N__36358),
            .I(\ppm_encoder_1.counterZ0Z_1 ));
    InMux I__7745 (
            .O(N__36351),
            .I(\ppm_encoder_1.un1_counter_13_cry_0 ));
    InMux I__7744 (
            .O(N__36348),
            .I(\ppm_encoder_1.un1_counter_13_cry_1 ));
    InMux I__7743 (
            .O(N__36345),
            .I(\ppm_encoder_1.un1_counter_13_cry_2 ));
    InMux I__7742 (
            .O(N__36342),
            .I(N__36337));
    InMux I__7741 (
            .O(N__36341),
            .I(N__36334));
    InMux I__7740 (
            .O(N__36340),
            .I(N__36331));
    LocalMux I__7739 (
            .O(N__36337),
            .I(\ppm_encoder_1.counterZ0Z_4 ));
    LocalMux I__7738 (
            .O(N__36334),
            .I(\ppm_encoder_1.counterZ0Z_4 ));
    LocalMux I__7737 (
            .O(N__36331),
            .I(\ppm_encoder_1.counterZ0Z_4 ));
    InMux I__7736 (
            .O(N__36324),
            .I(\ppm_encoder_1.un1_counter_13_cry_3 ));
    InMux I__7735 (
            .O(N__36321),
            .I(N__36316));
    InMux I__7734 (
            .O(N__36320),
            .I(N__36313));
    InMux I__7733 (
            .O(N__36319),
            .I(N__36310));
    LocalMux I__7732 (
            .O(N__36316),
            .I(\ppm_encoder_1.counterZ0Z_5 ));
    LocalMux I__7731 (
            .O(N__36313),
            .I(\ppm_encoder_1.counterZ0Z_5 ));
    LocalMux I__7730 (
            .O(N__36310),
            .I(\ppm_encoder_1.counterZ0Z_5 ));
    InMux I__7729 (
            .O(N__36303),
            .I(\ppm_encoder_1.un1_counter_13_cry_4 ));
    InMux I__7728 (
            .O(N__36300),
            .I(\ppm_encoder_1.un1_counter_13_cry_5 ));
    InMux I__7727 (
            .O(N__36297),
            .I(\ppm_encoder_1.un1_counter_13_cry_6 ));
    InMux I__7726 (
            .O(N__36294),
            .I(N__36291));
    LocalMux I__7725 (
            .O(N__36291),
            .I(N__36287));
    InMux I__7724 (
            .O(N__36290),
            .I(N__36284));
    Odrv12 I__7723 (
            .O(N__36287),
            .I(scaler_4_data_13));
    LocalMux I__7722 (
            .O(N__36284),
            .I(scaler_4_data_13));
    InMux I__7721 (
            .O(N__36279),
            .I(N__36276));
    LocalMux I__7720 (
            .O(N__36276),
            .I(N__36273));
    Span4Mux_h I__7719 (
            .O(N__36273),
            .I(N__36270));
    Odrv4 I__7718 (
            .O(N__36270),
            .I(\ppm_encoder_1.un1_rudder_cry_12_THRU_CO ));
    CEMux I__7717 (
            .O(N__36267),
            .I(N__36263));
    CEMux I__7716 (
            .O(N__36266),
            .I(N__36259));
    LocalMux I__7715 (
            .O(N__36263),
            .I(N__36256));
    CEMux I__7714 (
            .O(N__36262),
            .I(N__36253));
    LocalMux I__7713 (
            .O(N__36259),
            .I(N__36250));
    Span4Mux_v I__7712 (
            .O(N__36256),
            .I(N__36245));
    LocalMux I__7711 (
            .O(N__36253),
            .I(N__36245));
    Span4Mux_v I__7710 (
            .O(N__36250),
            .I(N__36241));
    Span4Mux_h I__7709 (
            .O(N__36245),
            .I(N__36238));
    CEMux I__7708 (
            .O(N__36244),
            .I(N__36235));
    Span4Mux_v I__7707 (
            .O(N__36241),
            .I(N__36228));
    Span4Mux_v I__7706 (
            .O(N__36238),
            .I(N__36228));
    LocalMux I__7705 (
            .O(N__36235),
            .I(N__36228));
    Span4Mux_h I__7704 (
            .O(N__36228),
            .I(N__36224));
    CEMux I__7703 (
            .O(N__36227),
            .I(N__36221));
    Odrv4 I__7702 (
            .O(N__36224),
            .I(\ppm_encoder_1.pid_altitude_dv_0 ));
    LocalMux I__7701 (
            .O(N__36221),
            .I(\ppm_encoder_1.pid_altitude_dv_0 ));
    CascadeMux I__7700 (
            .O(N__36216),
            .I(N__36213));
    InMux I__7699 (
            .O(N__36213),
            .I(N__36209));
    InMux I__7698 (
            .O(N__36212),
            .I(N__36206));
    LocalMux I__7697 (
            .O(N__36209),
            .I(N__36202));
    LocalMux I__7696 (
            .O(N__36206),
            .I(N__36199));
    InMux I__7695 (
            .O(N__36205),
            .I(N__36196));
    Span4Mux_v I__7694 (
            .O(N__36202),
            .I(N__36191));
    Span4Mux_v I__7693 (
            .O(N__36199),
            .I(N__36191));
    LocalMux I__7692 (
            .O(N__36196),
            .I(\ppm_encoder_1.rudderZ0Z_6 ));
    Odrv4 I__7691 (
            .O(N__36191),
            .I(\ppm_encoder_1.rudderZ0Z_6 ));
    InMux I__7690 (
            .O(N__36186),
            .I(N__36182));
    InMux I__7689 (
            .O(N__36185),
            .I(N__36179));
    LocalMux I__7688 (
            .O(N__36182),
            .I(N__36176));
    LocalMux I__7687 (
            .O(N__36179),
            .I(N__36173));
    Span4Mux_v I__7686 (
            .O(N__36176),
            .I(N__36170));
    Span4Mux_h I__7685 (
            .O(N__36173),
            .I(N__36167));
    Odrv4 I__7684 (
            .O(N__36170),
            .I(scaler_2_data_11));
    Odrv4 I__7683 (
            .O(N__36167),
            .I(scaler_2_data_11));
    InMux I__7682 (
            .O(N__36162),
            .I(N__36159));
    LocalMux I__7681 (
            .O(N__36159),
            .I(N__36156));
    Odrv4 I__7680 (
            .O(N__36156),
            .I(\ppm_encoder_1.un1_aileron_cry_10_THRU_CO ));
    InMux I__7679 (
            .O(N__36153),
            .I(N__36150));
    LocalMux I__7678 (
            .O(N__36150),
            .I(N__36145));
    InMux I__7677 (
            .O(N__36149),
            .I(N__36142));
    InMux I__7676 (
            .O(N__36148),
            .I(N__36139));
    Span4Mux_h I__7675 (
            .O(N__36145),
            .I(N__36136));
    LocalMux I__7674 (
            .O(N__36142),
            .I(\ppm_encoder_1.aileronZ0Z_11 ));
    LocalMux I__7673 (
            .O(N__36139),
            .I(\ppm_encoder_1.aileronZ0Z_11 ));
    Odrv4 I__7672 (
            .O(N__36136),
            .I(\ppm_encoder_1.aileronZ0Z_11 ));
    InMux I__7671 (
            .O(N__36129),
            .I(N__36126));
    LocalMux I__7670 (
            .O(N__36126),
            .I(N__36123));
    Span4Mux_v I__7669 (
            .O(N__36123),
            .I(N__36120));
    Odrv4 I__7668 (
            .O(N__36120),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_4 ));
    InMux I__7667 (
            .O(N__36117),
            .I(N__36114));
    LocalMux I__7666 (
            .O(N__36114),
            .I(\ppm_encoder_1.pulses2countZ0Z_4 ));
    InMux I__7665 (
            .O(N__36111),
            .I(N__36108));
    LocalMux I__7664 (
            .O(N__36108),
            .I(N__36105));
    Span12Mux_v I__7663 (
            .O(N__36105),
            .I(N__36102));
    Odrv12 I__7662 (
            .O(N__36102),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_5 ));
    CascadeMux I__7661 (
            .O(N__36099),
            .I(N__36096));
    InMux I__7660 (
            .O(N__36096),
            .I(N__36093));
    LocalMux I__7659 (
            .O(N__36093),
            .I(\ppm_encoder_1.pulses2countZ0Z_5 ));
    InMux I__7658 (
            .O(N__36090),
            .I(N__36087));
    LocalMux I__7657 (
            .O(N__36087),
            .I(N__36084));
    Odrv12 I__7656 (
            .O(N__36084),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_0 ));
    InMux I__7655 (
            .O(N__36081),
            .I(N__36078));
    LocalMux I__7654 (
            .O(N__36078),
            .I(N__36075));
    Odrv4 I__7653 (
            .O(N__36075),
            .I(\ppm_encoder_1.pulses2countZ0Z_0 ));
    InMux I__7652 (
            .O(N__36072),
            .I(N__36069));
    LocalMux I__7651 (
            .O(N__36069),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_1 ));
    InMux I__7650 (
            .O(N__36066),
            .I(N__36063));
    LocalMux I__7649 (
            .O(N__36063),
            .I(N__36060));
    Odrv12 I__7648 (
            .O(N__36060),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_1 ));
    InMux I__7647 (
            .O(N__36057),
            .I(N__36054));
    LocalMux I__7646 (
            .O(N__36054),
            .I(N__36051));
    Odrv4 I__7645 (
            .O(N__36051),
            .I(\ppm_encoder_1.pulses2countZ0Z_1 ));
    InMux I__7644 (
            .O(N__36048),
            .I(N__36044));
    InMux I__7643 (
            .O(N__36047),
            .I(N__36041));
    LocalMux I__7642 (
            .O(N__36044),
            .I(N__36038));
    LocalMux I__7641 (
            .O(N__36041),
            .I(N__36035));
    Span4Mux_v I__7640 (
            .O(N__36038),
            .I(N__36032));
    Odrv4 I__7639 (
            .O(N__36035),
            .I(scaler_2_data_8));
    Odrv4 I__7638 (
            .O(N__36032),
            .I(scaler_2_data_8));
    CascadeMux I__7637 (
            .O(N__36027),
            .I(N__36024));
    InMux I__7636 (
            .O(N__36024),
            .I(N__36021));
    LocalMux I__7635 (
            .O(N__36021),
            .I(\ppm_encoder_1.un1_aileron_cry_7_THRU_CO ));
    InMux I__7634 (
            .O(N__36018),
            .I(\ppm_encoder_1.un1_aileron_cry_7 ));
    InMux I__7633 (
            .O(N__36015),
            .I(N__36011));
    InMux I__7632 (
            .O(N__36014),
            .I(N__36008));
    LocalMux I__7631 (
            .O(N__36011),
            .I(N__36005));
    LocalMux I__7630 (
            .O(N__36008),
            .I(N__36000));
    Span4Mux_h I__7629 (
            .O(N__36005),
            .I(N__36000));
    Odrv4 I__7628 (
            .O(N__36000),
            .I(scaler_2_data_9));
    InMux I__7627 (
            .O(N__35997),
            .I(N__35994));
    LocalMux I__7626 (
            .O(N__35994),
            .I(N__35991));
    Odrv4 I__7625 (
            .O(N__35991),
            .I(\ppm_encoder_1.un1_aileron_cry_8_THRU_CO ));
    InMux I__7624 (
            .O(N__35988),
            .I(\ppm_encoder_1.un1_aileron_cry_8 ));
    InMux I__7623 (
            .O(N__35985),
            .I(N__35981));
    InMux I__7622 (
            .O(N__35984),
            .I(N__35978));
    LocalMux I__7621 (
            .O(N__35981),
            .I(N__35975));
    LocalMux I__7620 (
            .O(N__35978),
            .I(N__35972));
    Span4Mux_v I__7619 (
            .O(N__35975),
            .I(N__35967));
    Span4Mux_h I__7618 (
            .O(N__35972),
            .I(N__35967));
    Odrv4 I__7617 (
            .O(N__35967),
            .I(scaler_2_data_10));
    InMux I__7616 (
            .O(N__35964),
            .I(N__35961));
    LocalMux I__7615 (
            .O(N__35961),
            .I(N__35958));
    Span4Mux_v I__7614 (
            .O(N__35958),
            .I(N__35955));
    Odrv4 I__7613 (
            .O(N__35955),
            .I(\ppm_encoder_1.un1_aileron_cry_9_THRU_CO ));
    InMux I__7612 (
            .O(N__35952),
            .I(\ppm_encoder_1.un1_aileron_cry_9 ));
    InMux I__7611 (
            .O(N__35949),
            .I(\ppm_encoder_1.un1_aileron_cry_10 ));
    InMux I__7610 (
            .O(N__35946),
            .I(N__35942));
    InMux I__7609 (
            .O(N__35945),
            .I(N__35939));
    LocalMux I__7608 (
            .O(N__35942),
            .I(N__35936));
    LocalMux I__7607 (
            .O(N__35939),
            .I(N__35933));
    Span4Mux_h I__7606 (
            .O(N__35936),
            .I(N__35930));
    Span4Mux_h I__7605 (
            .O(N__35933),
            .I(N__35927));
    Odrv4 I__7604 (
            .O(N__35930),
            .I(scaler_2_data_12));
    Odrv4 I__7603 (
            .O(N__35927),
            .I(scaler_2_data_12));
    InMux I__7602 (
            .O(N__35922),
            .I(N__35919));
    LocalMux I__7601 (
            .O(N__35919),
            .I(N__35916));
    Span4Mux_h I__7600 (
            .O(N__35916),
            .I(N__35913));
    Odrv4 I__7599 (
            .O(N__35913),
            .I(\ppm_encoder_1.un1_aileron_cry_11_THRU_CO ));
    InMux I__7598 (
            .O(N__35910),
            .I(\ppm_encoder_1.un1_aileron_cry_11 ));
    CascadeMux I__7597 (
            .O(N__35907),
            .I(N__35903));
    InMux I__7596 (
            .O(N__35906),
            .I(N__35900));
    InMux I__7595 (
            .O(N__35903),
            .I(N__35897));
    LocalMux I__7594 (
            .O(N__35900),
            .I(N__35894));
    LocalMux I__7593 (
            .O(N__35897),
            .I(N__35891));
    Span4Mux_h I__7592 (
            .O(N__35894),
            .I(N__35888));
    Odrv4 I__7591 (
            .O(N__35891),
            .I(scaler_2_data_13));
    Odrv4 I__7590 (
            .O(N__35888),
            .I(scaler_2_data_13));
    InMux I__7589 (
            .O(N__35883),
            .I(N__35880));
    LocalMux I__7588 (
            .O(N__35880),
            .I(\ppm_encoder_1.un1_aileron_cry_12_THRU_CO ));
    InMux I__7587 (
            .O(N__35877),
            .I(\ppm_encoder_1.un1_aileron_cry_12 ));
    InMux I__7586 (
            .O(N__35874),
            .I(N__35871));
    LocalMux I__7585 (
            .O(N__35871),
            .I(N__35868));
    Span4Mux_h I__7584 (
            .O(N__35868),
            .I(N__35865));
    Odrv4 I__7583 (
            .O(N__35865),
            .I(scaler_2_data_14));
    InMux I__7582 (
            .O(N__35862),
            .I(bfn_16_16_0_));
    InMux I__7581 (
            .O(N__35859),
            .I(N__35855));
    CascadeMux I__7580 (
            .O(N__35858),
            .I(N__35852));
    LocalMux I__7579 (
            .O(N__35855),
            .I(N__35849));
    InMux I__7578 (
            .O(N__35852),
            .I(N__35845));
    Span4Mux_h I__7577 (
            .O(N__35849),
            .I(N__35842));
    InMux I__7576 (
            .O(N__35848),
            .I(N__35839));
    LocalMux I__7575 (
            .O(N__35845),
            .I(\ppm_encoder_1.rudderZ0Z_10 ));
    Odrv4 I__7574 (
            .O(N__35842),
            .I(\ppm_encoder_1.rudderZ0Z_10 ));
    LocalMux I__7573 (
            .O(N__35839),
            .I(\ppm_encoder_1.rudderZ0Z_10 ));
    CascadeMux I__7572 (
            .O(N__35832),
            .I(\ppm_encoder_1.un2_throttle_iv_1_5_cascade_ ));
    InMux I__7571 (
            .O(N__35829),
            .I(N__35826));
    LocalMux I__7570 (
            .O(N__35826),
            .I(N__35823));
    Odrv4 I__7569 (
            .O(N__35823),
            .I(\ppm_encoder_1.un2_throttle_iv_0_5 ));
    InMux I__7568 (
            .O(N__35820),
            .I(N__35815));
    InMux I__7567 (
            .O(N__35819),
            .I(N__35811));
    InMux I__7566 (
            .O(N__35818),
            .I(N__35808));
    LocalMux I__7565 (
            .O(N__35815),
            .I(N__35805));
    InMux I__7564 (
            .O(N__35814),
            .I(N__35802));
    LocalMux I__7563 (
            .O(N__35811),
            .I(N__35791));
    LocalMux I__7562 (
            .O(N__35808),
            .I(N__35791));
    Span4Mux_v I__7561 (
            .O(N__35805),
            .I(N__35791));
    LocalMux I__7560 (
            .O(N__35802),
            .I(N__35791));
    InMux I__7559 (
            .O(N__35801),
            .I(N__35788));
    InMux I__7558 (
            .O(N__35800),
            .I(N__35785));
    Span4Mux_v I__7557 (
            .O(N__35791),
            .I(N__35772));
    LocalMux I__7556 (
            .O(N__35788),
            .I(N__35772));
    LocalMux I__7555 (
            .O(N__35785),
            .I(N__35772));
    InMux I__7554 (
            .O(N__35784),
            .I(N__35769));
    InMux I__7553 (
            .O(N__35783),
            .I(N__35766));
    InMux I__7552 (
            .O(N__35782),
            .I(N__35761));
    InMux I__7551 (
            .O(N__35781),
            .I(N__35761));
    InMux I__7550 (
            .O(N__35780),
            .I(N__35756));
    InMux I__7549 (
            .O(N__35779),
            .I(N__35756));
    Odrv4 I__7548 (
            .O(N__35772),
            .I(\ppm_encoder_1.init_pulses_2_sqmuxa_0 ));
    LocalMux I__7547 (
            .O(N__35769),
            .I(\ppm_encoder_1.init_pulses_2_sqmuxa_0 ));
    LocalMux I__7546 (
            .O(N__35766),
            .I(\ppm_encoder_1.init_pulses_2_sqmuxa_0 ));
    LocalMux I__7545 (
            .O(N__35761),
            .I(\ppm_encoder_1.init_pulses_2_sqmuxa_0 ));
    LocalMux I__7544 (
            .O(N__35756),
            .I(\ppm_encoder_1.init_pulses_2_sqmuxa_0 ));
    InMux I__7543 (
            .O(N__35745),
            .I(N__35741));
    InMux I__7542 (
            .O(N__35744),
            .I(N__35738));
    LocalMux I__7541 (
            .O(N__35741),
            .I(N__35735));
    LocalMux I__7540 (
            .O(N__35738),
            .I(N__35723));
    Span4Mux_v I__7539 (
            .O(N__35735),
            .I(N__35723));
    InMux I__7538 (
            .O(N__35734),
            .I(N__35720));
    InMux I__7537 (
            .O(N__35733),
            .I(N__35717));
    InMux I__7536 (
            .O(N__35732),
            .I(N__35714));
    InMux I__7535 (
            .O(N__35731),
            .I(N__35711));
    InMux I__7534 (
            .O(N__35730),
            .I(N__35708));
    InMux I__7533 (
            .O(N__35729),
            .I(N__35703));
    InMux I__7532 (
            .O(N__35728),
            .I(N__35703));
    Span4Mux_v I__7531 (
            .O(N__35723),
            .I(N__35698));
    LocalMux I__7530 (
            .O(N__35720),
            .I(N__35698));
    LocalMux I__7529 (
            .O(N__35717),
            .I(N__35690));
    LocalMux I__7528 (
            .O(N__35714),
            .I(N__35690));
    LocalMux I__7527 (
            .O(N__35711),
            .I(N__35690));
    LocalMux I__7526 (
            .O(N__35708),
            .I(N__35685));
    LocalMux I__7525 (
            .O(N__35703),
            .I(N__35685));
    Span4Mux_v I__7524 (
            .O(N__35698),
            .I(N__35680));
    InMux I__7523 (
            .O(N__35697),
            .I(N__35677));
    Span4Mux_v I__7522 (
            .O(N__35690),
            .I(N__35672));
    Span4Mux_h I__7521 (
            .O(N__35685),
            .I(N__35672));
    InMux I__7520 (
            .O(N__35684),
            .I(N__35667));
    InMux I__7519 (
            .O(N__35683),
            .I(N__35667));
    Odrv4 I__7518 (
            .O(N__35680),
            .I(\ppm_encoder_1.init_pulses_1_sqmuxa_0 ));
    LocalMux I__7517 (
            .O(N__35677),
            .I(\ppm_encoder_1.init_pulses_1_sqmuxa_0 ));
    Odrv4 I__7516 (
            .O(N__35672),
            .I(\ppm_encoder_1.init_pulses_1_sqmuxa_0 ));
    LocalMux I__7515 (
            .O(N__35667),
            .I(\ppm_encoder_1.init_pulses_1_sqmuxa_0 ));
    CascadeMux I__7514 (
            .O(N__35658),
            .I(\ppm_encoder_1.un2_throttle_iv_1_14_cascade_ ));
    InMux I__7513 (
            .O(N__35655),
            .I(N__35652));
    LocalMux I__7512 (
            .O(N__35652),
            .I(\ppm_encoder_1.un2_throttle_iv_0_14 ));
    CascadeMux I__7511 (
            .O(N__35649),
            .I(N__35646));
    InMux I__7510 (
            .O(N__35646),
            .I(N__35642));
    InMux I__7509 (
            .O(N__35645),
            .I(N__35639));
    LocalMux I__7508 (
            .O(N__35642),
            .I(N__35636));
    LocalMux I__7507 (
            .O(N__35639),
            .I(N__35633));
    Span4Mux_h I__7506 (
            .O(N__35636),
            .I(N__35630));
    Odrv12 I__7505 (
            .O(N__35633),
            .I(\ppm_encoder_1.throttleZ0Z_14 ));
    Odrv4 I__7504 (
            .O(N__35630),
            .I(\ppm_encoder_1.throttleZ0Z_14 ));
    CascadeMux I__7503 (
            .O(N__35625),
            .I(N__35621));
    InMux I__7502 (
            .O(N__35624),
            .I(N__35616));
    InMux I__7501 (
            .O(N__35621),
            .I(N__35616));
    LocalMux I__7500 (
            .O(N__35616),
            .I(N__35613));
    Span4Mux_h I__7499 (
            .O(N__35613),
            .I(N__35610));
    Span4Mux_v I__7498 (
            .O(N__35610),
            .I(N__35607));
    Odrv4 I__7497 (
            .O(N__35607),
            .I(\ppm_encoder_1.elevatorZ0Z_14 ));
    InMux I__7496 (
            .O(N__35604),
            .I(N__35601));
    LocalMux I__7495 (
            .O(N__35601),
            .I(N__35597));
    InMux I__7494 (
            .O(N__35600),
            .I(N__35594));
    Span4Mux_h I__7493 (
            .O(N__35597),
            .I(N__35591));
    LocalMux I__7492 (
            .O(N__35594),
            .I(scaler_2_data_6));
    Odrv4 I__7491 (
            .O(N__35591),
            .I(scaler_2_data_6));
    InMux I__7490 (
            .O(N__35586),
            .I(N__35583));
    LocalMux I__7489 (
            .O(N__35583),
            .I(N__35579));
    InMux I__7488 (
            .O(N__35582),
            .I(N__35576));
    Span12Mux_s11_h I__7487 (
            .O(N__35579),
            .I(N__35573));
    LocalMux I__7486 (
            .O(N__35576),
            .I(scaler_2_data_7));
    Odrv12 I__7485 (
            .O(N__35573),
            .I(scaler_2_data_7));
    InMux I__7484 (
            .O(N__35568),
            .I(N__35565));
    LocalMux I__7483 (
            .O(N__35565),
            .I(N__35562));
    Span12Mux_h I__7482 (
            .O(N__35562),
            .I(N__35559));
    Odrv12 I__7481 (
            .O(N__35559),
            .I(\ppm_encoder_1.un1_aileron_cry_6_THRU_CO ));
    InMux I__7480 (
            .O(N__35556),
            .I(\ppm_encoder_1.un1_aileron_cry_6 ));
    CascadeMux I__7479 (
            .O(N__35553),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_3_cascade_ ));
    InMux I__7478 (
            .O(N__35550),
            .I(N__35544));
    InMux I__7477 (
            .O(N__35549),
            .I(N__35537));
    InMux I__7476 (
            .O(N__35548),
            .I(N__35537));
    InMux I__7475 (
            .O(N__35547),
            .I(N__35537));
    LocalMux I__7474 (
            .O(N__35544),
            .I(\ppm_encoder_1.init_pulsesZ0Z_3 ));
    LocalMux I__7473 (
            .O(N__35537),
            .I(\ppm_encoder_1.init_pulsesZ0Z_3 ));
    InMux I__7472 (
            .O(N__35532),
            .I(N__35528));
    CascadeMux I__7471 (
            .O(N__35531),
            .I(N__35524));
    LocalMux I__7470 (
            .O(N__35528),
            .I(N__35520));
    InMux I__7469 (
            .O(N__35527),
            .I(N__35517));
    InMux I__7468 (
            .O(N__35524),
            .I(N__35512));
    InMux I__7467 (
            .O(N__35523),
            .I(N__35512));
    Span4Mux_h I__7466 (
            .O(N__35520),
            .I(N__35509));
    LocalMux I__7465 (
            .O(N__35517),
            .I(N__35506));
    LocalMux I__7464 (
            .O(N__35512),
            .I(N__35503));
    Span4Mux_v I__7463 (
            .O(N__35509),
            .I(N__35500));
    Span4Mux_v I__7462 (
            .O(N__35506),
            .I(N__35497));
    Odrv4 I__7461 (
            .O(N__35503),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_10_mux ));
    Odrv4 I__7460 (
            .O(N__35500),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_10_mux ));
    Odrv4 I__7459 (
            .O(N__35497),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_10_mux ));
    InMux I__7458 (
            .O(N__35490),
            .I(N__35487));
    LocalMux I__7457 (
            .O(N__35487),
            .I(N__35484));
    Span4Mux_h I__7456 (
            .O(N__35484),
            .I(N__35481));
    Odrv4 I__7455 (
            .O(N__35481),
            .I(\ppm_encoder_1.un1_throttle_cry_2_THRU_CO ));
    InMux I__7454 (
            .O(N__35478),
            .I(N__35474));
    CascadeMux I__7453 (
            .O(N__35477),
            .I(N__35470));
    LocalMux I__7452 (
            .O(N__35474),
            .I(N__35467));
    InMux I__7451 (
            .O(N__35473),
            .I(N__35464));
    InMux I__7450 (
            .O(N__35470),
            .I(N__35461));
    Span4Mux_h I__7449 (
            .O(N__35467),
            .I(N__35456));
    LocalMux I__7448 (
            .O(N__35464),
            .I(N__35456));
    LocalMux I__7447 (
            .O(N__35461),
            .I(throttle_command_3));
    Odrv4 I__7446 (
            .O(N__35456),
            .I(throttle_command_3));
    InMux I__7445 (
            .O(N__35451),
            .I(N__35447));
    CascadeMux I__7444 (
            .O(N__35450),
            .I(N__35443));
    LocalMux I__7443 (
            .O(N__35447),
            .I(N__35440));
    InMux I__7442 (
            .O(N__35446),
            .I(N__35435));
    InMux I__7441 (
            .O(N__35443),
            .I(N__35435));
    Odrv4 I__7440 (
            .O(N__35440),
            .I(\ppm_encoder_1.throttleZ0Z_3 ));
    LocalMux I__7439 (
            .O(N__35435),
            .I(\ppm_encoder_1.throttleZ0Z_3 ));
    InMux I__7438 (
            .O(N__35430),
            .I(N__35426));
    InMux I__7437 (
            .O(N__35429),
            .I(N__35423));
    LocalMux I__7436 (
            .O(N__35426),
            .I(N__35420));
    LocalMux I__7435 (
            .O(N__35423),
            .I(N__35417));
    Span4Mux_h I__7434 (
            .O(N__35420),
            .I(N__35412));
    Span4Mux_h I__7433 (
            .O(N__35417),
            .I(N__35412));
    Odrv4 I__7432 (
            .O(N__35412),
            .I(\ppm_encoder_1.aileronZ0Z_5 ));
    CascadeMux I__7431 (
            .O(N__35409),
            .I(N__35405));
    InMux I__7430 (
            .O(N__35408),
            .I(N__35402));
    InMux I__7429 (
            .O(N__35405),
            .I(N__35399));
    LocalMux I__7428 (
            .O(N__35402),
            .I(N__35396));
    LocalMux I__7427 (
            .O(N__35399),
            .I(N__35393));
    Span4Mux_v I__7426 (
            .O(N__35396),
            .I(N__35388));
    Span4Mux_v I__7425 (
            .O(N__35393),
            .I(N__35388));
    Odrv4 I__7424 (
            .O(N__35388),
            .I(\ppm_encoder_1.elevatorZ0Z_5 ));
    CascadeMux I__7423 (
            .O(N__35385),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_10_mux_cascade_ ));
    CascadeMux I__7422 (
            .O(N__35382),
            .I(N__35379));
    InMux I__7421 (
            .O(N__35379),
            .I(N__35375));
    InMux I__7420 (
            .O(N__35378),
            .I(N__35371));
    LocalMux I__7419 (
            .O(N__35375),
            .I(N__35368));
    CascadeMux I__7418 (
            .O(N__35374),
            .I(N__35365));
    LocalMux I__7417 (
            .O(N__35371),
            .I(N__35360));
    Span4Mux_h I__7416 (
            .O(N__35368),
            .I(N__35360));
    InMux I__7415 (
            .O(N__35365),
            .I(N__35357));
    Span4Mux_v I__7414 (
            .O(N__35360),
            .I(N__35354));
    LocalMux I__7413 (
            .O(N__35357),
            .I(\ppm_encoder_1.throttleZ0Z_4 ));
    Odrv4 I__7412 (
            .O(N__35354),
            .I(\ppm_encoder_1.throttleZ0Z_4 ));
    CascadeMux I__7411 (
            .O(N__35349),
            .I(\ppm_encoder_1.un2_throttle_iv_0_4_cascade_ ));
    InMux I__7410 (
            .O(N__35346),
            .I(N__35343));
    LocalMux I__7409 (
            .O(N__35343),
            .I(\ppm_encoder_1.un2_throttle_iv_1_4 ));
    CascadeMux I__7408 (
            .O(N__35340),
            .I(N__35335));
    InMux I__7407 (
            .O(N__35339),
            .I(N__35330));
    InMux I__7406 (
            .O(N__35338),
            .I(N__35330));
    InMux I__7405 (
            .O(N__35335),
            .I(N__35327));
    LocalMux I__7404 (
            .O(N__35330),
            .I(N__35322));
    LocalMux I__7403 (
            .O(N__35327),
            .I(N__35322));
    Odrv4 I__7402 (
            .O(N__35322),
            .I(\ppm_encoder_1.throttleZ0Z_7 ));
    InMux I__7401 (
            .O(N__35319),
            .I(N__35316));
    LocalMux I__7400 (
            .O(N__35316),
            .I(N__35313));
    Odrv4 I__7399 (
            .O(N__35313),
            .I(\ppm_encoder_1.un2_throttle_iv_0_7 ));
    InMux I__7398 (
            .O(N__35310),
            .I(N__35302));
    InMux I__7397 (
            .O(N__35309),
            .I(N__35302));
    InMux I__7396 (
            .O(N__35308),
            .I(N__35299));
    InMux I__7395 (
            .O(N__35307),
            .I(N__35296));
    LocalMux I__7394 (
            .O(N__35302),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2 ));
    LocalMux I__7393 (
            .O(N__35299),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2 ));
    LocalMux I__7392 (
            .O(N__35296),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2 ));
    InMux I__7391 (
            .O(N__35289),
            .I(N__35282));
    InMux I__7390 (
            .O(N__35288),
            .I(N__35279));
    InMux I__7389 (
            .O(N__35287),
            .I(N__35276));
    InMux I__7388 (
            .O(N__35286),
            .I(N__35273));
    InMux I__7387 (
            .O(N__35285),
            .I(N__35270));
    LocalMux I__7386 (
            .O(N__35282),
            .I(N__35256));
    LocalMux I__7385 (
            .O(N__35279),
            .I(N__35256));
    LocalMux I__7384 (
            .O(N__35276),
            .I(N__35256));
    LocalMux I__7383 (
            .O(N__35273),
            .I(N__35256));
    LocalMux I__7382 (
            .O(N__35270),
            .I(N__35256));
    InMux I__7381 (
            .O(N__35269),
            .I(N__35251));
    InMux I__7380 (
            .O(N__35268),
            .I(N__35251));
    InMux I__7379 (
            .O(N__35267),
            .I(N__35245));
    Span4Mux_v I__7378 (
            .O(N__35256),
            .I(N__35240));
    LocalMux I__7377 (
            .O(N__35251),
            .I(N__35240));
    InMux I__7376 (
            .O(N__35250),
            .I(N__35233));
    InMux I__7375 (
            .O(N__35249),
            .I(N__35233));
    InMux I__7374 (
            .O(N__35248),
            .I(N__35233));
    LocalMux I__7373 (
            .O(N__35245),
            .I(\ppm_encoder_1.init_pulses_3_sqmuxa_0 ));
    Odrv4 I__7372 (
            .O(N__35240),
            .I(\ppm_encoder_1.init_pulses_3_sqmuxa_0 ));
    LocalMux I__7371 (
            .O(N__35233),
            .I(\ppm_encoder_1.init_pulses_3_sqmuxa_0 ));
    CascadeMux I__7370 (
            .O(N__35226),
            .I(N__35223));
    InMux I__7369 (
            .O(N__35223),
            .I(N__35219));
    InMux I__7368 (
            .O(N__35222),
            .I(N__35215));
    LocalMux I__7367 (
            .O(N__35219),
            .I(N__35212));
    InMux I__7366 (
            .O(N__35218),
            .I(N__35209));
    LocalMux I__7365 (
            .O(N__35215),
            .I(N__35206));
    Span4Mux_h I__7364 (
            .O(N__35212),
            .I(N__35203));
    LocalMux I__7363 (
            .O(N__35209),
            .I(\ppm_encoder_1.throttleZ0Z_5 ));
    Odrv12 I__7362 (
            .O(N__35206),
            .I(\ppm_encoder_1.throttleZ0Z_5 ));
    Odrv4 I__7361 (
            .O(N__35203),
            .I(\ppm_encoder_1.throttleZ0Z_5 ));
    CascadeMux I__7360 (
            .O(N__35196),
            .I(N__35193));
    InMux I__7359 (
            .O(N__35193),
            .I(N__35189));
    InMux I__7358 (
            .O(N__35192),
            .I(N__35186));
    LocalMux I__7357 (
            .O(N__35189),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_ns_3 ));
    LocalMux I__7356 (
            .O(N__35186),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_ns_3 ));
    InMux I__7355 (
            .O(N__35181),
            .I(N__35177));
    InMux I__7354 (
            .O(N__35180),
            .I(N__35174));
    LocalMux I__7353 (
            .O(N__35177),
            .I(\reset_module_System.countZ0Z_15 ));
    LocalMux I__7352 (
            .O(N__35174),
            .I(\reset_module_System.countZ0Z_15 ));
    CascadeMux I__7351 (
            .O(N__35169),
            .I(N__35165));
    InMux I__7350 (
            .O(N__35168),
            .I(N__35160));
    InMux I__7349 (
            .O(N__35165),
            .I(N__35160));
    LocalMux I__7348 (
            .O(N__35160),
            .I(\reset_module_System.countZ0Z_21 ));
    InMux I__7347 (
            .O(N__35157),
            .I(N__35153));
    InMux I__7346 (
            .O(N__35156),
            .I(N__35150));
    LocalMux I__7345 (
            .O(N__35153),
            .I(\reset_module_System.countZ0Z_13 ));
    LocalMux I__7344 (
            .O(N__35150),
            .I(\reset_module_System.countZ0Z_13 ));
    CascadeMux I__7343 (
            .O(N__35145),
            .I(N__35142));
    InMux I__7342 (
            .O(N__35142),
            .I(N__35139));
    LocalMux I__7341 (
            .O(N__35139),
            .I(\reset_module_System.reset6_11 ));
    CascadeMux I__7340 (
            .O(N__35136),
            .I(\ppm_encoder_1.N_297_cascade_ ));
    CascadeMux I__7339 (
            .O(N__35133),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_159_d_cascade_ ));
    InMux I__7338 (
            .O(N__35130),
            .I(N__35125));
    InMux I__7337 (
            .O(N__35129),
            .I(N__35122));
    InMux I__7336 (
            .O(N__35128),
            .I(N__35119));
    LocalMux I__7335 (
            .O(N__35125),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_3 ));
    LocalMux I__7334 (
            .O(N__35122),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_3 ));
    LocalMux I__7333 (
            .O(N__35119),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_3 ));
    InMux I__7332 (
            .O(N__35112),
            .I(\reset_module_System.count_1_cry_13 ));
    InMux I__7331 (
            .O(N__35109),
            .I(\reset_module_System.count_1_cry_14 ));
    InMux I__7330 (
            .O(N__35106),
            .I(N__35102));
    InMux I__7329 (
            .O(N__35105),
            .I(N__35099));
    LocalMux I__7328 (
            .O(N__35102),
            .I(\reset_module_System.countZ0Z_16 ));
    LocalMux I__7327 (
            .O(N__35099),
            .I(\reset_module_System.countZ0Z_16 ));
    InMux I__7326 (
            .O(N__35094),
            .I(\reset_module_System.count_1_cry_15 ));
    InMux I__7325 (
            .O(N__35091),
            .I(bfn_16_9_0_));
    InMux I__7324 (
            .O(N__35088),
            .I(N__35084));
    InMux I__7323 (
            .O(N__35087),
            .I(N__35081));
    LocalMux I__7322 (
            .O(N__35084),
            .I(N__35078));
    LocalMux I__7321 (
            .O(N__35081),
            .I(\reset_module_System.countZ0Z_18 ));
    Odrv4 I__7320 (
            .O(N__35078),
            .I(\reset_module_System.countZ0Z_18 ));
    InMux I__7319 (
            .O(N__35073),
            .I(\reset_module_System.count_1_cry_17 ));
    InMux I__7318 (
            .O(N__35070),
            .I(\reset_module_System.count_1_cry_18 ));
    CascadeMux I__7317 (
            .O(N__35067),
            .I(N__35063));
    InMux I__7316 (
            .O(N__35066),
            .I(N__35060));
    InMux I__7315 (
            .O(N__35063),
            .I(N__35057));
    LocalMux I__7314 (
            .O(N__35060),
            .I(\reset_module_System.countZ0Z_20 ));
    LocalMux I__7313 (
            .O(N__35057),
            .I(\reset_module_System.countZ0Z_20 ));
    InMux I__7312 (
            .O(N__35052),
            .I(\reset_module_System.count_1_cry_19 ));
    InMux I__7311 (
            .O(N__35049),
            .I(\reset_module_System.count_1_cry_20 ));
    CascadeMux I__7310 (
            .O(N__35046),
            .I(N__35043));
    InMux I__7309 (
            .O(N__35043),
            .I(N__35037));
    InMux I__7308 (
            .O(N__35042),
            .I(N__35037));
    LocalMux I__7307 (
            .O(N__35037),
            .I(\reset_module_System.countZ0Z_19 ));
    InMux I__7306 (
            .O(N__35034),
            .I(N__35030));
    InMux I__7305 (
            .O(N__35033),
            .I(N__35027));
    LocalMux I__7304 (
            .O(N__35030),
            .I(\reset_module_System.countZ0Z_5 ));
    LocalMux I__7303 (
            .O(N__35027),
            .I(\reset_module_System.countZ0Z_5 ));
    InMux I__7302 (
            .O(N__35022),
            .I(\reset_module_System.count_1_cry_4 ));
    InMux I__7301 (
            .O(N__35019),
            .I(N__35015));
    InMux I__7300 (
            .O(N__35018),
            .I(N__35012));
    LocalMux I__7299 (
            .O(N__35015),
            .I(\reset_module_System.countZ0Z_6 ));
    LocalMux I__7298 (
            .O(N__35012),
            .I(\reset_module_System.countZ0Z_6 ));
    InMux I__7297 (
            .O(N__35007),
            .I(\reset_module_System.count_1_cry_5 ));
    InMux I__7296 (
            .O(N__35004),
            .I(N__35000));
    InMux I__7295 (
            .O(N__35003),
            .I(N__34997));
    LocalMux I__7294 (
            .O(N__35000),
            .I(\reset_module_System.countZ0Z_7 ));
    LocalMux I__7293 (
            .O(N__34997),
            .I(\reset_module_System.countZ0Z_7 ));
    InMux I__7292 (
            .O(N__34992),
            .I(\reset_module_System.count_1_cry_6 ));
    InMux I__7291 (
            .O(N__34989),
            .I(N__34985));
    InMux I__7290 (
            .O(N__34988),
            .I(N__34982));
    LocalMux I__7289 (
            .O(N__34985),
            .I(\reset_module_System.countZ0Z_8 ));
    LocalMux I__7288 (
            .O(N__34982),
            .I(\reset_module_System.countZ0Z_8 ));
    InMux I__7287 (
            .O(N__34977),
            .I(\reset_module_System.count_1_cry_7 ));
    CascadeMux I__7286 (
            .O(N__34974),
            .I(N__34971));
    InMux I__7285 (
            .O(N__34971),
            .I(N__34967));
    InMux I__7284 (
            .O(N__34970),
            .I(N__34964));
    LocalMux I__7283 (
            .O(N__34967),
            .I(N__34961));
    LocalMux I__7282 (
            .O(N__34964),
            .I(\reset_module_System.countZ0Z_9 ));
    Odrv4 I__7281 (
            .O(N__34961),
            .I(\reset_module_System.countZ0Z_9 ));
    InMux I__7280 (
            .O(N__34956),
            .I(bfn_16_8_0_));
    InMux I__7279 (
            .O(N__34953),
            .I(\reset_module_System.count_1_cry_9 ));
    InMux I__7278 (
            .O(N__34950),
            .I(\reset_module_System.count_1_cry_10 ));
    InMux I__7277 (
            .O(N__34947),
            .I(N__34943));
    InMux I__7276 (
            .O(N__34946),
            .I(N__34940));
    LocalMux I__7275 (
            .O(N__34943),
            .I(\reset_module_System.countZ0Z_12 ));
    LocalMux I__7274 (
            .O(N__34940),
            .I(\reset_module_System.countZ0Z_12 ));
    InMux I__7273 (
            .O(N__34935),
            .I(\reset_module_System.count_1_cry_11 ));
    InMux I__7272 (
            .O(N__34932),
            .I(\reset_module_System.count_1_cry_12 ));
    CascadeMux I__7271 (
            .O(N__34929),
            .I(N__34925));
    CascadeMux I__7270 (
            .O(N__34928),
            .I(N__34922));
    InMux I__7269 (
            .O(N__34925),
            .I(N__34918));
    InMux I__7268 (
            .O(N__34922),
            .I(N__34915));
    InMux I__7267 (
            .O(N__34921),
            .I(N__34912));
    LocalMux I__7266 (
            .O(N__34918),
            .I(N__34909));
    LocalMux I__7265 (
            .O(N__34915),
            .I(\ppm_encoder_1.elevatorZ0Z_11 ));
    LocalMux I__7264 (
            .O(N__34912),
            .I(\ppm_encoder_1.elevatorZ0Z_11 ));
    Odrv4 I__7263 (
            .O(N__34909),
            .I(\ppm_encoder_1.elevatorZ0Z_11 ));
    InMux I__7262 (
            .O(N__34902),
            .I(N__34899));
    LocalMux I__7261 (
            .O(N__34899),
            .I(N__34896));
    Odrv4 I__7260 (
            .O(N__34896),
            .I(\ppm_encoder_1.un2_throttle_iv_1_11 ));
    InMux I__7259 (
            .O(N__34893),
            .I(N__34889));
    InMux I__7258 (
            .O(N__34892),
            .I(N__34886));
    LocalMux I__7257 (
            .O(N__34889),
            .I(\ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_5_0 ));
    LocalMux I__7256 (
            .O(N__34886),
            .I(\ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_5_0 ));
    InMux I__7255 (
            .O(N__34881),
            .I(N__34878));
    LocalMux I__7254 (
            .O(N__34878),
            .I(N__34875));
    Span4Mux_v I__7253 (
            .O(N__34875),
            .I(N__34872));
    Sp12to4 I__7252 (
            .O(N__34872),
            .I(N__34869));
    Odrv12 I__7251 (
            .O(N__34869),
            .I(\pid_alt.O_0_5 ));
    CascadeMux I__7250 (
            .O(N__34866),
            .I(N__34863));
    InMux I__7249 (
            .O(N__34863),
            .I(N__34860));
    LocalMux I__7248 (
            .O(N__34860),
            .I(N__34857));
    Odrv4 I__7247 (
            .O(N__34857),
            .I(\pid_alt.error_i_regZ0Z_1 ));
    InMux I__7246 (
            .O(N__34854),
            .I(N__34850));
    InMux I__7245 (
            .O(N__34853),
            .I(N__34846));
    LocalMux I__7244 (
            .O(N__34850),
            .I(N__34843));
    InMux I__7243 (
            .O(N__34849),
            .I(N__34840));
    LocalMux I__7242 (
            .O(N__34846),
            .I(\reset_module_System.countZ0Z_1 ));
    Odrv12 I__7241 (
            .O(N__34843),
            .I(\reset_module_System.countZ0Z_1 ));
    LocalMux I__7240 (
            .O(N__34840),
            .I(\reset_module_System.countZ0Z_1 ));
    CascadeMux I__7239 (
            .O(N__34833),
            .I(N__34828));
    InMux I__7238 (
            .O(N__34832),
            .I(N__34825));
    InMux I__7237 (
            .O(N__34831),
            .I(N__34822));
    InMux I__7236 (
            .O(N__34828),
            .I(N__34819));
    LocalMux I__7235 (
            .O(N__34825),
            .I(N__34815));
    LocalMux I__7234 (
            .O(N__34822),
            .I(N__34812));
    LocalMux I__7233 (
            .O(N__34819),
            .I(N__34809));
    InMux I__7232 (
            .O(N__34818),
            .I(N__34806));
    Span4Mux_v I__7231 (
            .O(N__34815),
            .I(N__34803));
    Sp12to4 I__7230 (
            .O(N__34812),
            .I(N__34798));
    Span12Mux_s8_v I__7229 (
            .O(N__34809),
            .I(N__34798));
    LocalMux I__7228 (
            .O(N__34806),
            .I(\reset_module_System.countZ0Z_0 ));
    Odrv4 I__7227 (
            .O(N__34803),
            .I(\reset_module_System.countZ0Z_0 ));
    Odrv12 I__7226 (
            .O(N__34798),
            .I(\reset_module_System.countZ0Z_0 ));
    InMux I__7225 (
            .O(N__34791),
            .I(N__34787));
    InMux I__7224 (
            .O(N__34790),
            .I(N__34784));
    LocalMux I__7223 (
            .O(N__34787),
            .I(\reset_module_System.countZ0Z_2 ));
    LocalMux I__7222 (
            .O(N__34784),
            .I(\reset_module_System.countZ0Z_2 ));
    InMux I__7221 (
            .O(N__34779),
            .I(N__34776));
    LocalMux I__7220 (
            .O(N__34776),
            .I(\reset_module_System.count_1_2 ));
    InMux I__7219 (
            .O(N__34773),
            .I(\reset_module_System.count_1_cry_1 ));
    InMux I__7218 (
            .O(N__34770),
            .I(N__34766));
    InMux I__7217 (
            .O(N__34769),
            .I(N__34763));
    LocalMux I__7216 (
            .O(N__34766),
            .I(\reset_module_System.countZ0Z_3 ));
    LocalMux I__7215 (
            .O(N__34763),
            .I(\reset_module_System.countZ0Z_3 ));
    InMux I__7214 (
            .O(N__34758),
            .I(\reset_module_System.count_1_cry_2 ));
    InMux I__7213 (
            .O(N__34755),
            .I(N__34751));
    InMux I__7212 (
            .O(N__34754),
            .I(N__34748));
    LocalMux I__7211 (
            .O(N__34751),
            .I(N__34745));
    LocalMux I__7210 (
            .O(N__34748),
            .I(\reset_module_System.countZ0Z_4 ));
    Odrv4 I__7209 (
            .O(N__34745),
            .I(\reset_module_System.countZ0Z_4 ));
    InMux I__7208 (
            .O(N__34740),
            .I(\reset_module_System.count_1_cry_3 ));
    InMux I__7207 (
            .O(N__34737),
            .I(N__34732));
    InMux I__7206 (
            .O(N__34736),
            .I(N__34727));
    InMux I__7205 (
            .O(N__34735),
            .I(N__34727));
    LocalMux I__7204 (
            .O(N__34732),
            .I(\ppm_encoder_1.aileronZ0Z_10 ));
    LocalMux I__7203 (
            .O(N__34727),
            .I(\ppm_encoder_1.aileronZ0Z_10 ));
    InMux I__7202 (
            .O(N__34722),
            .I(N__34719));
    LocalMux I__7201 (
            .O(N__34719),
            .I(\ppm_encoder_1.N_145_17 ));
    CascadeMux I__7200 (
            .O(N__34716),
            .I(\ppm_encoder_1.N_145_17_cascade_ ));
    InMux I__7199 (
            .O(N__34713),
            .I(N__34704));
    InMux I__7198 (
            .O(N__34712),
            .I(N__34704));
    InMux I__7197 (
            .O(N__34711),
            .I(N__34704));
    LocalMux I__7196 (
            .O(N__34704),
            .I(\ppm_encoder_1.N_238 ));
    CascadeMux I__7195 (
            .O(N__34701),
            .I(N__34698));
    InMux I__7194 (
            .O(N__34698),
            .I(N__34695));
    LocalMux I__7193 (
            .O(N__34695),
            .I(\ppm_encoder_1.un1_PPM_STATE_1_sqmuxa_i_a3_0_1 ));
    InMux I__7192 (
            .O(N__34692),
            .I(N__34689));
    LocalMux I__7191 (
            .O(N__34689),
            .I(\ppm_encoder_1.un2_throttle_iv_1_10 ));
    InMux I__7190 (
            .O(N__34686),
            .I(N__34683));
    LocalMux I__7189 (
            .O(N__34683),
            .I(\ppm_encoder_1.un2_throttle_iv_0_10 ));
    InMux I__7188 (
            .O(N__34680),
            .I(N__34676));
    CascadeMux I__7187 (
            .O(N__34679),
            .I(N__34672));
    LocalMux I__7186 (
            .O(N__34676),
            .I(N__34668));
    InMux I__7185 (
            .O(N__34675),
            .I(N__34665));
    InMux I__7184 (
            .O(N__34672),
            .I(N__34660));
    InMux I__7183 (
            .O(N__34671),
            .I(N__34660));
    Odrv4 I__7182 (
            .O(N__34668),
            .I(\ppm_encoder_1.PPM_STATEZ0Z_1 ));
    LocalMux I__7181 (
            .O(N__34665),
            .I(\ppm_encoder_1.PPM_STATEZ0Z_1 ));
    LocalMux I__7180 (
            .O(N__34660),
            .I(\ppm_encoder_1.PPM_STATEZ0Z_1 ));
    InMux I__7179 (
            .O(N__34653),
            .I(N__34650));
    LocalMux I__7178 (
            .O(N__34650),
            .I(\ppm_encoder_1.PPM_STATE_ns_0_a3_0_1_0 ));
    CascadeMux I__7177 (
            .O(N__34647),
            .I(N__34644));
    InMux I__7176 (
            .O(N__34644),
            .I(N__34641));
    LocalMux I__7175 (
            .O(N__34641),
            .I(\ppm_encoder_1.PPM_STATE_ns_0_a3_0_17_4_0 ));
    InMux I__7174 (
            .O(N__34638),
            .I(N__34635));
    LocalMux I__7173 (
            .O(N__34635),
            .I(\ppm_encoder_1.PPM_STATE_ns_0_a3_0_17_3_0 ));
    CascadeMux I__7172 (
            .O(N__34632),
            .I(N__34627));
    InMux I__7171 (
            .O(N__34631),
            .I(N__34624));
    InMux I__7170 (
            .O(N__34630),
            .I(N__34619));
    InMux I__7169 (
            .O(N__34627),
            .I(N__34619));
    LocalMux I__7168 (
            .O(N__34624),
            .I(\ppm_encoder_1.throttleZ0Z_11 ));
    LocalMux I__7167 (
            .O(N__34619),
            .I(\ppm_encoder_1.throttleZ0Z_11 ));
    CascadeMux I__7166 (
            .O(N__34614),
            .I(\ppm_encoder_1.N_303_cascade_ ));
    InMux I__7165 (
            .O(N__34611),
            .I(N__34608));
    LocalMux I__7164 (
            .O(N__34608),
            .I(\ppm_encoder_1.un2_throttle_iv_0_11 ));
    CascadeMux I__7163 (
            .O(N__34605),
            .I(N__34602));
    InMux I__7162 (
            .O(N__34602),
            .I(N__34597));
    InMux I__7161 (
            .O(N__34601),
            .I(N__34594));
    InMux I__7160 (
            .O(N__34600),
            .I(N__34591));
    LocalMux I__7159 (
            .O(N__34597),
            .I(\ppm_encoder_1.rudderZ0Z_11 ));
    LocalMux I__7158 (
            .O(N__34594),
            .I(\ppm_encoder_1.rudderZ0Z_11 ));
    LocalMux I__7157 (
            .O(N__34591),
            .I(\ppm_encoder_1.rudderZ0Z_11 ));
    CascadeMux I__7156 (
            .O(N__34584),
            .I(\ppm_encoder_1.N_319_cascade_ ));
    InMux I__7155 (
            .O(N__34581),
            .I(N__34578));
    LocalMux I__7154 (
            .O(N__34578),
            .I(N__34574));
    InMux I__7153 (
            .O(N__34577),
            .I(N__34571));
    Span4Mux_h I__7152 (
            .O(N__34574),
            .I(N__34567));
    LocalMux I__7151 (
            .O(N__34571),
            .I(N__34564));
    InMux I__7150 (
            .O(N__34570),
            .I(N__34561));
    Span4Mux_v I__7149 (
            .O(N__34567),
            .I(N__34558));
    Span4Mux_h I__7148 (
            .O(N__34564),
            .I(N__34555));
    LocalMux I__7147 (
            .O(N__34561),
            .I(\ppm_encoder_1.throttleZ0Z_1 ));
    Odrv4 I__7146 (
            .O(N__34558),
            .I(\ppm_encoder_1.throttleZ0Z_1 ));
    Odrv4 I__7145 (
            .O(N__34555),
            .I(\ppm_encoder_1.throttleZ0Z_1 ));
    InMux I__7144 (
            .O(N__34548),
            .I(N__34545));
    LocalMux I__7143 (
            .O(N__34545),
            .I(\ppm_encoder_1.N_302 ));
    InMux I__7142 (
            .O(N__34542),
            .I(N__34539));
    LocalMux I__7141 (
            .O(N__34539),
            .I(N__34536));
    Span4Mux_v I__7140 (
            .O(N__34536),
            .I(N__34533));
    Span4Mux_v I__7139 (
            .O(N__34533),
            .I(N__34530));
    Odrv4 I__7138 (
            .O(N__34530),
            .I(\ppm_encoder_1.un1_rudder_cry_7_THRU_CO ));
    InMux I__7137 (
            .O(N__34527),
            .I(N__34524));
    LocalMux I__7136 (
            .O(N__34524),
            .I(N__34521));
    Span4Mux_h I__7135 (
            .O(N__34521),
            .I(N__34517));
    InMux I__7134 (
            .O(N__34520),
            .I(N__34514));
    Odrv4 I__7133 (
            .O(N__34517),
            .I(scaler_4_data_8));
    LocalMux I__7132 (
            .O(N__34514),
            .I(scaler_4_data_8));
    CascadeMux I__7131 (
            .O(N__34509),
            .I(\ppm_encoder_1.un2_throttle_iv_0_13_cascade_ ));
    InMux I__7130 (
            .O(N__34506),
            .I(N__34503));
    LocalMux I__7129 (
            .O(N__34503),
            .I(\ppm_encoder_1.un2_throttle_iv_1_13 ));
    InMux I__7128 (
            .O(N__34500),
            .I(N__34496));
    InMux I__7127 (
            .O(N__34499),
            .I(N__34493));
    LocalMux I__7126 (
            .O(N__34496),
            .I(N__34490));
    LocalMux I__7125 (
            .O(N__34493),
            .I(N__34487));
    Span4Mux_v I__7124 (
            .O(N__34490),
            .I(N__34484));
    Span4Mux_v I__7123 (
            .O(N__34487),
            .I(N__34481));
    Odrv4 I__7122 (
            .O(N__34484),
            .I(scaler_3_data_13));
    Odrv4 I__7121 (
            .O(N__34481),
            .I(scaler_3_data_13));
    InMux I__7120 (
            .O(N__34476),
            .I(N__34473));
    LocalMux I__7119 (
            .O(N__34473),
            .I(N__34470));
    Span4Mux_h I__7118 (
            .O(N__34470),
            .I(N__34467));
    Odrv4 I__7117 (
            .O(N__34467),
            .I(\ppm_encoder_1.un1_elevator_cry_12_THRU_CO ));
    InMux I__7116 (
            .O(N__34464),
            .I(N__34461));
    LocalMux I__7115 (
            .O(N__34461),
            .I(N__34457));
    InMux I__7114 (
            .O(N__34460),
            .I(N__34454));
    Span4Mux_v I__7113 (
            .O(N__34457),
            .I(N__34449));
    LocalMux I__7112 (
            .O(N__34454),
            .I(N__34449));
    Span4Mux_h I__7111 (
            .O(N__34449),
            .I(N__34446));
    Span4Mux_h I__7110 (
            .O(N__34446),
            .I(N__34443));
    Odrv4 I__7109 (
            .O(N__34443),
            .I(throttle_command_13));
    CascadeMux I__7108 (
            .O(N__34440),
            .I(N__34437));
    InMux I__7107 (
            .O(N__34437),
            .I(N__34434));
    LocalMux I__7106 (
            .O(N__34434),
            .I(N__34431));
    Span4Mux_h I__7105 (
            .O(N__34431),
            .I(N__34428));
    Odrv4 I__7104 (
            .O(N__34428),
            .I(\ppm_encoder_1.un1_throttle_cry_12_THRU_CO ));
    CascadeMux I__7103 (
            .O(N__34425),
            .I(N__34420));
    InMux I__7102 (
            .O(N__34424),
            .I(N__34417));
    InMux I__7101 (
            .O(N__34423),
            .I(N__34412));
    InMux I__7100 (
            .O(N__34420),
            .I(N__34412));
    LocalMux I__7099 (
            .O(N__34417),
            .I(\ppm_encoder_1.throttleZ0Z_13 ));
    LocalMux I__7098 (
            .O(N__34412),
            .I(\ppm_encoder_1.throttleZ0Z_13 ));
    CascadeMux I__7097 (
            .O(N__34407),
            .I(N__34402));
    InMux I__7096 (
            .O(N__34406),
            .I(N__34399));
    InMux I__7095 (
            .O(N__34405),
            .I(N__34394));
    InMux I__7094 (
            .O(N__34402),
            .I(N__34394));
    LocalMux I__7093 (
            .O(N__34399),
            .I(\ppm_encoder_1.elevatorZ0Z_13 ));
    LocalMux I__7092 (
            .O(N__34394),
            .I(\ppm_encoder_1.elevatorZ0Z_13 ));
    CascadeMux I__7091 (
            .O(N__34389),
            .I(\ppm_encoder_1.N_305_cascade_ ));
    InMux I__7090 (
            .O(N__34386),
            .I(N__34381));
    InMux I__7089 (
            .O(N__34385),
            .I(N__34376));
    InMux I__7088 (
            .O(N__34384),
            .I(N__34376));
    LocalMux I__7087 (
            .O(N__34381),
            .I(\ppm_encoder_1.aileronZ0Z_13 ));
    LocalMux I__7086 (
            .O(N__34376),
            .I(\ppm_encoder_1.aileronZ0Z_13 ));
    CascadeMux I__7085 (
            .O(N__34371),
            .I(\ppm_encoder_1.N_298_cascade_ ));
    InMux I__7084 (
            .O(N__34368),
            .I(N__34359));
    InMux I__7083 (
            .O(N__34367),
            .I(N__34359));
    InMux I__7082 (
            .O(N__34366),
            .I(N__34359));
    LocalMux I__7081 (
            .O(N__34359),
            .I(\ppm_encoder_1.aileronZ0Z_6 ));
    InMux I__7080 (
            .O(N__34356),
            .I(N__34352));
    InMux I__7079 (
            .O(N__34355),
            .I(N__34349));
    LocalMux I__7078 (
            .O(N__34352),
            .I(N__34346));
    LocalMux I__7077 (
            .O(N__34349),
            .I(N__34343));
    Span4Mux_v I__7076 (
            .O(N__34346),
            .I(N__34340));
    Odrv12 I__7075 (
            .O(N__34343),
            .I(scaler_3_data_6));
    Odrv4 I__7074 (
            .O(N__34340),
            .I(scaler_3_data_6));
    CascadeMux I__7073 (
            .O(N__34335),
            .I(N__34330));
    InMux I__7072 (
            .O(N__34334),
            .I(N__34323));
    InMux I__7071 (
            .O(N__34333),
            .I(N__34323));
    InMux I__7070 (
            .O(N__34330),
            .I(N__34323));
    LocalMux I__7069 (
            .O(N__34323),
            .I(\ppm_encoder_1.elevatorZ0Z_6 ));
    InMux I__7068 (
            .O(N__34320),
            .I(N__34317));
    LocalMux I__7067 (
            .O(N__34317),
            .I(N__34314));
    Span4Mux_h I__7066 (
            .O(N__34314),
            .I(N__34311));
    Odrv4 I__7065 (
            .O(N__34311),
            .I(\ppm_encoder_1.un1_throttle_cry_5_THRU_CO ));
    InMux I__7064 (
            .O(N__34308),
            .I(N__34304));
    CascadeMux I__7063 (
            .O(N__34307),
            .I(N__34301));
    LocalMux I__7062 (
            .O(N__34304),
            .I(N__34298));
    InMux I__7061 (
            .O(N__34301),
            .I(N__34295));
    Span4Mux_h I__7060 (
            .O(N__34298),
            .I(N__34292));
    LocalMux I__7059 (
            .O(N__34295),
            .I(N__34289));
    Span4Mux_h I__7058 (
            .O(N__34292),
            .I(N__34286));
    Span4Mux_h I__7057 (
            .O(N__34289),
            .I(N__34283));
    Odrv4 I__7056 (
            .O(N__34286),
            .I(throttle_command_6));
    Odrv4 I__7055 (
            .O(N__34283),
            .I(throttle_command_6));
    InMux I__7054 (
            .O(N__34278),
            .I(N__34271));
    InMux I__7053 (
            .O(N__34277),
            .I(N__34271));
    InMux I__7052 (
            .O(N__34276),
            .I(N__34268));
    LocalMux I__7051 (
            .O(N__34271),
            .I(\ppm_encoder_1.throttleZ0Z_6 ));
    LocalMux I__7050 (
            .O(N__34268),
            .I(\ppm_encoder_1.throttleZ0Z_6 ));
    CascadeMux I__7049 (
            .O(N__34263),
            .I(\ppm_encoder_1.un2_throttle_iv_1_8_cascade_ ));
    InMux I__7048 (
            .O(N__34260),
            .I(N__34257));
    LocalMux I__7047 (
            .O(N__34257),
            .I(N__34254));
    Odrv12 I__7046 (
            .O(N__34254),
            .I(\ppm_encoder_1.un2_throttle_iv_0_8 ));
    CascadeMux I__7045 (
            .O(N__34251),
            .I(N__34247));
    InMux I__7044 (
            .O(N__34250),
            .I(N__34242));
    InMux I__7043 (
            .O(N__34247),
            .I(N__34242));
    LocalMux I__7042 (
            .O(N__34242),
            .I(N__34238));
    InMux I__7041 (
            .O(N__34241),
            .I(N__34235));
    Span4Mux_h I__7040 (
            .O(N__34238),
            .I(N__34232));
    LocalMux I__7039 (
            .O(N__34235),
            .I(\ppm_encoder_1.elevatorZ0Z_8 ));
    Odrv4 I__7038 (
            .O(N__34232),
            .I(\ppm_encoder_1.elevatorZ0Z_8 ));
    InMux I__7037 (
            .O(N__34227),
            .I(N__34224));
    LocalMux I__7036 (
            .O(N__34224),
            .I(N__34220));
    InMux I__7035 (
            .O(N__34223),
            .I(N__34217));
    Span4Mux_h I__7034 (
            .O(N__34220),
            .I(N__34214));
    LocalMux I__7033 (
            .O(N__34217),
            .I(N__34211));
    Span4Mux_h I__7032 (
            .O(N__34214),
            .I(N__34208));
    Span4Mux_h I__7031 (
            .O(N__34211),
            .I(N__34205));
    Odrv4 I__7030 (
            .O(N__34208),
            .I(throttle_command_8));
    Odrv4 I__7029 (
            .O(N__34205),
            .I(throttle_command_8));
    InMux I__7028 (
            .O(N__34200),
            .I(N__34197));
    LocalMux I__7027 (
            .O(N__34197),
            .I(N__34194));
    Span4Mux_h I__7026 (
            .O(N__34194),
            .I(N__34191));
    Odrv4 I__7025 (
            .O(N__34191),
            .I(\ppm_encoder_1.un1_throttle_cry_7_THRU_CO ));
    CascadeMux I__7024 (
            .O(N__34188),
            .I(N__34185));
    InMux I__7023 (
            .O(N__34185),
            .I(N__34180));
    InMux I__7022 (
            .O(N__34184),
            .I(N__34175));
    InMux I__7021 (
            .O(N__34183),
            .I(N__34175));
    LocalMux I__7020 (
            .O(N__34180),
            .I(N__34172));
    LocalMux I__7019 (
            .O(N__34175),
            .I(\ppm_encoder_1.throttleZ0Z_8 ));
    Odrv12 I__7018 (
            .O(N__34172),
            .I(\ppm_encoder_1.throttleZ0Z_8 ));
    InMux I__7017 (
            .O(N__34167),
            .I(N__34163));
    CascadeMux I__7016 (
            .O(N__34166),
            .I(N__34160));
    LocalMux I__7015 (
            .O(N__34163),
            .I(N__34157));
    InMux I__7014 (
            .O(N__34160),
            .I(N__34154));
    Span4Mux_v I__7013 (
            .O(N__34157),
            .I(N__34149));
    LocalMux I__7012 (
            .O(N__34154),
            .I(N__34149));
    Odrv4 I__7011 (
            .O(N__34149),
            .I(\ppm_encoder_1.elevatorZ0Z_4 ));
    CascadeMux I__7010 (
            .O(N__34146),
            .I(\ppm_encoder_1.N_296_cascade_ ));
    InMux I__7009 (
            .O(N__34143),
            .I(N__34140));
    LocalMux I__7008 (
            .O(N__34140),
            .I(N__34136));
    InMux I__7007 (
            .O(N__34139),
            .I(N__34133));
    Span4Mux_v I__7006 (
            .O(N__34136),
            .I(N__34128));
    LocalMux I__7005 (
            .O(N__34133),
            .I(N__34128));
    Odrv4 I__7004 (
            .O(N__34128),
            .I(\ppm_encoder_1.aileronZ0Z_4 ));
    CascadeMux I__7003 (
            .O(N__34125),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_0_cascade_ ));
    CascadeMux I__7002 (
            .O(N__34122),
            .I(\ppm_encoder_1.un2_throttle_iv_1_6_cascade_ ));
    InMux I__7001 (
            .O(N__34119),
            .I(N__34116));
    LocalMux I__7000 (
            .O(N__34116),
            .I(\ppm_encoder_1.un2_throttle_iv_0_6 ));
    CascadeMux I__6999 (
            .O(N__34113),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_d_4_cascade_ ));
    CascadeMux I__6998 (
            .O(N__34110),
            .I(\ppm_encoder_1.N_227_cascade_ ));
    CascadeMux I__6997 (
            .O(N__34107),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1Z0Z_0_cascade_ ));
    CascadeMux I__6996 (
            .O(N__34104),
            .I(N__34101));
    InMux I__6995 (
            .O(N__34101),
            .I(N__34095));
    InMux I__6994 (
            .O(N__34100),
            .I(N__34095));
    LocalMux I__6993 (
            .O(N__34095),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_d_4 ));
    CascadeMux I__6992 (
            .O(N__34092),
            .I(\ppm_encoder_1.un2_throttle_iv_1_1_cascade_ ));
    InMux I__6991 (
            .O(N__34089),
            .I(N__34086));
    LocalMux I__6990 (
            .O(N__34086),
            .I(N__34083));
    Span4Mux_h I__6989 (
            .O(N__34083),
            .I(N__34080));
    Odrv4 I__6988 (
            .O(N__34080),
            .I(\uart_drone.data_Auxce_0_0_2 ));
    InMux I__6987 (
            .O(N__34077),
            .I(N__34074));
    LocalMux I__6986 (
            .O(N__34074),
            .I(N__34071));
    Odrv12 I__6985 (
            .O(N__34071),
            .I(\uart_drone.data_Auxce_0_6 ));
    InMux I__6984 (
            .O(N__34068),
            .I(N__34065));
    LocalMux I__6983 (
            .O(N__34065),
            .I(N__34061));
    CascadeMux I__6982 (
            .O(N__34064),
            .I(N__34057));
    Span4Mux_v I__6981 (
            .O(N__34061),
            .I(N__34054));
    InMux I__6980 (
            .O(N__34060),
            .I(N__34049));
    InMux I__6979 (
            .O(N__34057),
            .I(N__34049));
    Odrv4 I__6978 (
            .O(N__34054),
            .I(\ppm_encoder_1.throttleZ0Z_12 ));
    LocalMux I__6977 (
            .O(N__34049),
            .I(\ppm_encoder_1.throttleZ0Z_12 ));
    InMux I__6976 (
            .O(N__34044),
            .I(N__34041));
    LocalMux I__6975 (
            .O(N__34041),
            .I(N__34037));
    CascadeMux I__6974 (
            .O(N__34040),
            .I(N__34033));
    Span4Mux_v I__6973 (
            .O(N__34037),
            .I(N__34030));
    InMux I__6972 (
            .O(N__34036),
            .I(N__34025));
    InMux I__6971 (
            .O(N__34033),
            .I(N__34025));
    Odrv4 I__6970 (
            .O(N__34030),
            .I(\ppm_encoder_1.elevatorZ0Z_12 ));
    LocalMux I__6969 (
            .O(N__34025),
            .I(\ppm_encoder_1.elevatorZ0Z_12 ));
    InMux I__6968 (
            .O(N__34020),
            .I(N__34017));
    LocalMux I__6967 (
            .O(N__34017),
            .I(N__34014));
    Span4Mux_v I__6966 (
            .O(N__34014),
            .I(N__34011));
    Odrv4 I__6965 (
            .O(N__34011),
            .I(\ppm_encoder_1.N_304 ));
    InMux I__6964 (
            .O(N__34008),
            .I(N__34005));
    LocalMux I__6963 (
            .O(N__34005),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_ns_2 ));
    CascadeMux I__6962 (
            .O(N__34002),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_ns_2_cascade_ ));
    InMux I__6961 (
            .O(N__33999),
            .I(N__33994));
    InMux I__6960 (
            .O(N__33998),
            .I(N__33991));
    InMux I__6959 (
            .O(N__33997),
            .I(N__33988));
    LocalMux I__6958 (
            .O(N__33994),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0 ));
    LocalMux I__6957 (
            .O(N__33991),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0 ));
    LocalMux I__6956 (
            .O(N__33988),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0 ));
    CascadeMux I__6955 (
            .O(N__33981),
            .I(N__33976));
    CascadeMux I__6954 (
            .O(N__33980),
            .I(N__33973));
    CascadeMux I__6953 (
            .O(N__33979),
            .I(N__33970));
    InMux I__6952 (
            .O(N__33976),
            .I(N__33967));
    InMux I__6951 (
            .O(N__33973),
            .I(N__33962));
    InMux I__6950 (
            .O(N__33970),
            .I(N__33962));
    LocalMux I__6949 (
            .O(N__33967),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_1 ));
    LocalMux I__6948 (
            .O(N__33962),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_1 ));
    CascadeMux I__6947 (
            .O(N__33957),
            .I(N__33951));
    InMux I__6946 (
            .O(N__33956),
            .I(N__33948));
    InMux I__6945 (
            .O(N__33955),
            .I(N__33945));
    InMux I__6944 (
            .O(N__33954),
            .I(N__33940));
    InMux I__6943 (
            .O(N__33951),
            .I(N__33940));
    LocalMux I__6942 (
            .O(N__33948),
            .I(\uart_drone.timer_CountZ0Z_0 ));
    LocalMux I__6941 (
            .O(N__33945),
            .I(\uart_drone.timer_CountZ0Z_0 ));
    LocalMux I__6940 (
            .O(N__33940),
            .I(\uart_drone.timer_CountZ0Z_0 ));
    CascadeMux I__6939 (
            .O(N__33933),
            .I(\uart_drone.timer_Count_RNO_0_0_1_cascade_ ));
    InMux I__6938 (
            .O(N__33930),
            .I(N__33926));
    InMux I__6937 (
            .O(N__33929),
            .I(N__33923));
    LocalMux I__6936 (
            .O(N__33926),
            .I(\uart_drone.timer_CountZ1Z_1 ));
    LocalMux I__6935 (
            .O(N__33923),
            .I(\uart_drone.timer_CountZ1Z_1 ));
    InMux I__6934 (
            .O(N__33918),
            .I(N__33908));
    InMux I__6933 (
            .O(N__33917),
            .I(N__33908));
    InMux I__6932 (
            .O(N__33916),
            .I(N__33905));
    InMux I__6931 (
            .O(N__33915),
            .I(N__33902));
    InMux I__6930 (
            .O(N__33914),
            .I(N__33899));
    InMux I__6929 (
            .O(N__33913),
            .I(N__33896));
    LocalMux I__6928 (
            .O(N__33908),
            .I(\uart_drone.N_143 ));
    LocalMux I__6927 (
            .O(N__33905),
            .I(\uart_drone.N_143 ));
    LocalMux I__6926 (
            .O(N__33902),
            .I(\uart_drone.N_143 ));
    LocalMux I__6925 (
            .O(N__33899),
            .I(\uart_drone.N_143 ));
    LocalMux I__6924 (
            .O(N__33896),
            .I(\uart_drone.N_143 ));
    CascadeMux I__6923 (
            .O(N__33885),
            .I(N__33881));
    CascadeMux I__6922 (
            .O(N__33884),
            .I(N__33878));
    InMux I__6921 (
            .O(N__33881),
            .I(N__33875));
    InMux I__6920 (
            .O(N__33878),
            .I(N__33872));
    LocalMux I__6919 (
            .O(N__33875),
            .I(N__33864));
    LocalMux I__6918 (
            .O(N__33872),
            .I(N__33864));
    InMux I__6917 (
            .O(N__33871),
            .I(N__33859));
    InMux I__6916 (
            .O(N__33870),
            .I(N__33859));
    InMux I__6915 (
            .O(N__33869),
            .I(N__33856));
    Odrv4 I__6914 (
            .O(N__33864),
            .I(\uart_drone.timer_Count_0_sqmuxa ));
    LocalMux I__6913 (
            .O(N__33859),
            .I(\uart_drone.timer_Count_0_sqmuxa ));
    LocalMux I__6912 (
            .O(N__33856),
            .I(\uart_drone.timer_Count_0_sqmuxa ));
    CascadeMux I__6911 (
            .O(N__33849),
            .I(N__33846));
    InMux I__6910 (
            .O(N__33846),
            .I(N__33843));
    LocalMux I__6909 (
            .O(N__33843),
            .I(N__33837));
    InMux I__6908 (
            .O(N__33842),
            .I(N__33834));
    CascadeMux I__6907 (
            .O(N__33841),
            .I(N__33831));
    InMux I__6906 (
            .O(N__33840),
            .I(N__33828));
    Span4Mux_v I__6905 (
            .O(N__33837),
            .I(N__33823));
    LocalMux I__6904 (
            .O(N__33834),
            .I(N__33823));
    InMux I__6903 (
            .O(N__33831),
            .I(N__33820));
    LocalMux I__6902 (
            .O(N__33828),
            .I(N__33817));
    Span4Mux_h I__6901 (
            .O(N__33823),
            .I(N__33814));
    LocalMux I__6900 (
            .O(N__33820),
            .I(N__33811));
    Span4Mux_h I__6899 (
            .O(N__33817),
            .I(N__33808));
    Odrv4 I__6898 (
            .O(N__33814),
            .I(\reset_module_System.reset6_15 ));
    Odrv4 I__6897 (
            .O(N__33811),
            .I(\reset_module_System.reset6_15 ));
    Odrv4 I__6896 (
            .O(N__33808),
            .I(\reset_module_System.reset6_15 ));
    InMux I__6895 (
            .O(N__33801),
            .I(N__33798));
    LocalMux I__6894 (
            .O(N__33798),
            .I(N__33795));
    Odrv4 I__6893 (
            .O(N__33795),
            .I(\reset_module_System.reset6_17 ));
    InMux I__6892 (
            .O(N__33792),
            .I(N__33788));
    InMux I__6891 (
            .O(N__33791),
            .I(N__33783));
    LocalMux I__6890 (
            .O(N__33788),
            .I(N__33780));
    InMux I__6889 (
            .O(N__33787),
            .I(N__33777));
    InMux I__6888 (
            .O(N__33786),
            .I(N__33774));
    LocalMux I__6887 (
            .O(N__33783),
            .I(N__33771));
    Span4Mux_h I__6886 (
            .O(N__33780),
            .I(N__33768));
    LocalMux I__6885 (
            .O(N__33777),
            .I(N__33765));
    LocalMux I__6884 (
            .O(N__33774),
            .I(N__33760));
    Span12Mux_s8_v I__6883 (
            .O(N__33771),
            .I(N__33760));
    Odrv4 I__6882 (
            .O(N__33768),
            .I(\reset_module_System.reset6_19 ));
    Odrv4 I__6881 (
            .O(N__33765),
            .I(\reset_module_System.reset6_19 ));
    Odrv12 I__6880 (
            .O(N__33760),
            .I(\reset_module_System.reset6_19 ));
    CascadeMux I__6879 (
            .O(N__33753),
            .I(N__33747));
    CascadeMux I__6878 (
            .O(N__33752),
            .I(N__33744));
    InMux I__6877 (
            .O(N__33751),
            .I(N__33741));
    InMux I__6876 (
            .O(N__33750),
            .I(N__33738));
    InMux I__6875 (
            .O(N__33747),
            .I(N__33735));
    InMux I__6874 (
            .O(N__33744),
            .I(N__33732));
    LocalMux I__6873 (
            .O(N__33741),
            .I(\uart_drone.stateZ0Z_2 ));
    LocalMux I__6872 (
            .O(N__33738),
            .I(\uart_drone.stateZ0Z_2 ));
    LocalMux I__6871 (
            .O(N__33735),
            .I(\uart_drone.stateZ0Z_2 ));
    LocalMux I__6870 (
            .O(N__33732),
            .I(\uart_drone.stateZ0Z_2 ));
    CascadeMux I__6869 (
            .O(N__33723),
            .I(\uart_drone.N_145_cascade_ ));
    SRMux I__6868 (
            .O(N__33720),
            .I(N__33715));
    SRMux I__6867 (
            .O(N__33719),
            .I(N__33712));
    SRMux I__6866 (
            .O(N__33718),
            .I(N__33709));
    LocalMux I__6865 (
            .O(N__33715),
            .I(N__33704));
    LocalMux I__6864 (
            .O(N__33712),
            .I(N__33704));
    LocalMux I__6863 (
            .O(N__33709),
            .I(N__33700));
    Span4Mux_v I__6862 (
            .O(N__33704),
            .I(N__33697));
    SRMux I__6861 (
            .O(N__33703),
            .I(N__33694));
    Span4Mux_v I__6860 (
            .O(N__33700),
            .I(N__33690));
    Span4Mux_h I__6859 (
            .O(N__33697),
            .I(N__33687));
    LocalMux I__6858 (
            .O(N__33694),
            .I(N__33684));
    SRMux I__6857 (
            .O(N__33693),
            .I(N__33681));
    Odrv4 I__6856 (
            .O(N__33690),
            .I(\pid_alt.un1_reset_1_0_i ));
    Odrv4 I__6855 (
            .O(N__33687),
            .I(\pid_alt.un1_reset_1_0_i ));
    Odrv12 I__6854 (
            .O(N__33684),
            .I(\pid_alt.un1_reset_1_0_i ));
    LocalMux I__6853 (
            .O(N__33681),
            .I(\pid_alt.un1_reset_1_0_i ));
    InMux I__6852 (
            .O(N__33672),
            .I(N__33669));
    LocalMux I__6851 (
            .O(N__33669),
            .I(N__33666));
    Span4Mux_v I__6850 (
            .O(N__33666),
            .I(N__33662));
    InMux I__6849 (
            .O(N__33665),
            .I(N__33659));
    Odrv4 I__6848 (
            .O(N__33662),
            .I(\pid_alt.error_i_acummZ0Z_0 ));
    LocalMux I__6847 (
            .O(N__33659),
            .I(\pid_alt.error_i_acummZ0Z_0 ));
    InMux I__6846 (
            .O(N__33654),
            .I(N__33650));
    InMux I__6845 (
            .O(N__33653),
            .I(N__33647));
    LocalMux I__6844 (
            .O(N__33650),
            .I(N__33644));
    LocalMux I__6843 (
            .O(N__33647),
            .I(N__33641));
    Span4Mux_v I__6842 (
            .O(N__33644),
            .I(N__33638));
    Span4Mux_h I__6841 (
            .O(N__33641),
            .I(N__33635));
    Odrv4 I__6840 (
            .O(N__33638),
            .I(\pid_alt.error_i_acumm_preregZ0Z_0 ));
    Odrv4 I__6839 (
            .O(N__33635),
            .I(\pid_alt.error_i_acumm_preregZ0Z_0 ));
    CEMux I__6838 (
            .O(N__33630),
            .I(N__33531));
    CEMux I__6837 (
            .O(N__33629),
            .I(N__33531));
    CEMux I__6836 (
            .O(N__33628),
            .I(N__33531));
    CEMux I__6835 (
            .O(N__33627),
            .I(N__33531));
    CEMux I__6834 (
            .O(N__33626),
            .I(N__33531));
    CEMux I__6833 (
            .O(N__33625),
            .I(N__33531));
    CEMux I__6832 (
            .O(N__33624),
            .I(N__33531));
    CEMux I__6831 (
            .O(N__33623),
            .I(N__33531));
    CEMux I__6830 (
            .O(N__33622),
            .I(N__33531));
    CEMux I__6829 (
            .O(N__33621),
            .I(N__33531));
    CEMux I__6828 (
            .O(N__33620),
            .I(N__33531));
    CEMux I__6827 (
            .O(N__33619),
            .I(N__33531));
    CEMux I__6826 (
            .O(N__33618),
            .I(N__33531));
    CEMux I__6825 (
            .O(N__33617),
            .I(N__33531));
    CEMux I__6824 (
            .O(N__33616),
            .I(N__33531));
    CEMux I__6823 (
            .O(N__33615),
            .I(N__33531));
    CEMux I__6822 (
            .O(N__33614),
            .I(N__33531));
    CEMux I__6821 (
            .O(N__33613),
            .I(N__33531));
    CEMux I__6820 (
            .O(N__33612),
            .I(N__33531));
    CEMux I__6819 (
            .O(N__33611),
            .I(N__33531));
    CEMux I__6818 (
            .O(N__33610),
            .I(N__33531));
    CEMux I__6817 (
            .O(N__33609),
            .I(N__33531));
    CEMux I__6816 (
            .O(N__33608),
            .I(N__33531));
    CEMux I__6815 (
            .O(N__33607),
            .I(N__33531));
    CEMux I__6814 (
            .O(N__33606),
            .I(N__33531));
    CEMux I__6813 (
            .O(N__33605),
            .I(N__33531));
    CEMux I__6812 (
            .O(N__33604),
            .I(N__33531));
    CEMux I__6811 (
            .O(N__33603),
            .I(N__33531));
    CEMux I__6810 (
            .O(N__33602),
            .I(N__33531));
    CEMux I__6809 (
            .O(N__33601),
            .I(N__33531));
    CEMux I__6808 (
            .O(N__33600),
            .I(N__33531));
    CEMux I__6807 (
            .O(N__33599),
            .I(N__33531));
    CEMux I__6806 (
            .O(N__33598),
            .I(N__33531));
    GlobalMux I__6805 (
            .O(N__33531),
            .I(N__33528));
    gio2CtrlBuf I__6804 (
            .O(N__33528),
            .I(\pid_alt.state_0_g_0 ));
    CascadeMux I__6803 (
            .O(N__33525),
            .I(N__33522));
    InMux I__6802 (
            .O(N__33522),
            .I(N__33519));
    LocalMux I__6801 (
            .O(N__33519),
            .I(N__33516));
    Span4Mux_h I__6800 (
            .O(N__33516),
            .I(N__33513));
    Odrv4 I__6799 (
            .O(N__33513),
            .I(\uart_drone.un1_state_2_0_a3_0 ));
    InMux I__6798 (
            .O(N__33510),
            .I(N__33505));
    InMux I__6797 (
            .O(N__33509),
            .I(N__33502));
    InMux I__6796 (
            .O(N__33508),
            .I(N__33499));
    LocalMux I__6795 (
            .O(N__33505),
            .I(N__33496));
    LocalMux I__6794 (
            .O(N__33502),
            .I(\uart_drone.timer_CountZ1Z_2 ));
    LocalMux I__6793 (
            .O(N__33499),
            .I(\uart_drone.timer_CountZ1Z_2 ));
    Odrv4 I__6792 (
            .O(N__33496),
            .I(\uart_drone.timer_CountZ1Z_2 ));
    InMux I__6791 (
            .O(N__33489),
            .I(N__33486));
    LocalMux I__6790 (
            .O(N__33486),
            .I(\uart_drone.timer_Count_RNO_0_0_2 ));
    InMux I__6789 (
            .O(N__33483),
            .I(\uart_drone.un4_timer_Count_1_cry_1 ));
    InMux I__6788 (
            .O(N__33480),
            .I(N__33477));
    LocalMux I__6787 (
            .O(N__33477),
            .I(N__33474));
    Span4Mux_v I__6786 (
            .O(N__33474),
            .I(N__33471));
    Odrv4 I__6785 (
            .O(N__33471),
            .I(\uart_drone.timer_Count_RNO_0_0_3 ));
    InMux I__6784 (
            .O(N__33468),
            .I(\uart_drone.un4_timer_Count_1_cry_2 ));
    InMux I__6783 (
            .O(N__33465),
            .I(\uart_drone.un4_timer_Count_1_cry_3 ));
    InMux I__6782 (
            .O(N__33462),
            .I(N__33459));
    LocalMux I__6781 (
            .O(N__33459),
            .I(N__33456));
    Span4Mux_v I__6780 (
            .O(N__33456),
            .I(N__33453));
    Odrv4 I__6779 (
            .O(N__33453),
            .I(\uart_drone.timer_Count_RNO_0_0_4 ));
    CascadeMux I__6778 (
            .O(N__33450),
            .I(\reset_module_System.reset6_13_cascade_ ));
    InMux I__6777 (
            .O(N__33447),
            .I(N__33444));
    LocalMux I__6776 (
            .O(N__33444),
            .I(\reset_module_System.reset6_3 ));
    InMux I__6775 (
            .O(N__33441),
            .I(N__33436));
    InMux I__6774 (
            .O(N__33440),
            .I(N__33432));
    InMux I__6773 (
            .O(N__33439),
            .I(N__33429));
    LocalMux I__6772 (
            .O(N__33436),
            .I(N__33426));
    InMux I__6771 (
            .O(N__33435),
            .I(N__33423));
    LocalMux I__6770 (
            .O(N__33432),
            .I(N__33420));
    LocalMux I__6769 (
            .O(N__33429),
            .I(N__33417));
    Span4Mux_v I__6768 (
            .O(N__33426),
            .I(N__33414));
    LocalMux I__6767 (
            .O(N__33423),
            .I(N__33410));
    Span4Mux_v I__6766 (
            .O(N__33420),
            .I(N__33406));
    Span4Mux_v I__6765 (
            .O(N__33417),
            .I(N__33401));
    Span4Mux_h I__6764 (
            .O(N__33414),
            .I(N__33398));
    InMux I__6763 (
            .O(N__33413),
            .I(N__33395));
    Span4Mux_v I__6762 (
            .O(N__33410),
            .I(N__33390));
    InMux I__6761 (
            .O(N__33409),
            .I(N__33386));
    Span4Mux_h I__6760 (
            .O(N__33406),
            .I(N__33383));
    InMux I__6759 (
            .O(N__33405),
            .I(N__33380));
    CascadeMux I__6758 (
            .O(N__33404),
            .I(N__33377));
    Span4Mux_h I__6757 (
            .O(N__33401),
            .I(N__33374));
    Span4Mux_v I__6756 (
            .O(N__33398),
            .I(N__33369));
    LocalMux I__6755 (
            .O(N__33395),
            .I(N__33369));
    InMux I__6754 (
            .O(N__33394),
            .I(N__33366));
    InMux I__6753 (
            .O(N__33393),
            .I(N__33363));
    Span4Mux_v I__6752 (
            .O(N__33390),
            .I(N__33359));
    InMux I__6751 (
            .O(N__33389),
            .I(N__33356));
    LocalMux I__6750 (
            .O(N__33386),
            .I(N__33349));
    Span4Mux_v I__6749 (
            .O(N__33383),
            .I(N__33349));
    LocalMux I__6748 (
            .O(N__33380),
            .I(N__33349));
    InMux I__6747 (
            .O(N__33377),
            .I(N__33346));
    Span4Mux_h I__6746 (
            .O(N__33374),
            .I(N__33336));
    Span4Mux_v I__6745 (
            .O(N__33369),
            .I(N__33336));
    LocalMux I__6744 (
            .O(N__33366),
            .I(N__33336));
    LocalMux I__6743 (
            .O(N__33363),
            .I(N__33336));
    InMux I__6742 (
            .O(N__33362),
            .I(N__33333));
    Sp12to4 I__6741 (
            .O(N__33359),
            .I(N__33330));
    LocalMux I__6740 (
            .O(N__33356),
            .I(N__33325));
    Span4Mux_v I__6739 (
            .O(N__33349),
            .I(N__33325));
    LocalMux I__6738 (
            .O(N__33346),
            .I(N__33322));
    InMux I__6737 (
            .O(N__33345),
            .I(N__33319));
    Sp12to4 I__6736 (
            .O(N__33336),
            .I(N__33312));
    LocalMux I__6735 (
            .O(N__33333),
            .I(N__33312));
    Span12Mux_h I__6734 (
            .O(N__33330),
            .I(N__33312));
    Span4Mux_v I__6733 (
            .O(N__33325),
            .I(N__33307));
    Span4Mux_v I__6732 (
            .O(N__33322),
            .I(N__33307));
    LocalMux I__6731 (
            .O(N__33319),
            .I(uart_pc_data_6));
    Odrv12 I__6730 (
            .O(N__33312),
            .I(uart_pc_data_6));
    Odrv4 I__6729 (
            .O(N__33307),
            .I(uart_pc_data_6));
    InMux I__6728 (
            .O(N__33300),
            .I(N__33297));
    LocalMux I__6727 (
            .O(N__33297),
            .I(N__33294));
    Span4Mux_s2_h I__6726 (
            .O(N__33294),
            .I(N__33291));
    Span4Mux_h I__6725 (
            .O(N__33291),
            .I(N__33288));
    Span4Mux_h I__6724 (
            .O(N__33288),
            .I(N__33285));
    Odrv4 I__6723 (
            .O(N__33285),
            .I(alt_ki_6));
    InMux I__6722 (
            .O(N__33282),
            .I(N__33279));
    LocalMux I__6721 (
            .O(N__33279),
            .I(N__33276));
    Span4Mux_h I__6720 (
            .O(N__33276),
            .I(N__33271));
    InMux I__6719 (
            .O(N__33275),
            .I(N__33266));
    InMux I__6718 (
            .O(N__33274),
            .I(N__33266));
    Odrv4 I__6717 (
            .O(N__33271),
            .I(\pid_alt.error_i_acumm_preregZ0Z_6 ));
    LocalMux I__6716 (
            .O(N__33266),
            .I(\pid_alt.error_i_acumm_preregZ0Z_6 ));
    CascadeMux I__6715 (
            .O(N__33261),
            .I(N__33257));
    InMux I__6714 (
            .O(N__33260),
            .I(N__33254));
    InMux I__6713 (
            .O(N__33257),
            .I(N__33251));
    LocalMux I__6712 (
            .O(N__33254),
            .I(\pid_alt.error_i_acummZ0Z_6 ));
    LocalMux I__6711 (
            .O(N__33251),
            .I(\pid_alt.error_i_acummZ0Z_6 ));
    CascadeMux I__6710 (
            .O(N__33246),
            .I(N__33241));
    CascadeMux I__6709 (
            .O(N__33245),
            .I(N__33237));
    CascadeMux I__6708 (
            .O(N__33244),
            .I(N__33232));
    InMux I__6707 (
            .O(N__33241),
            .I(N__33224));
    InMux I__6706 (
            .O(N__33240),
            .I(N__33224));
    InMux I__6705 (
            .O(N__33237),
            .I(N__33219));
    InMux I__6704 (
            .O(N__33236),
            .I(N__33219));
    InMux I__6703 (
            .O(N__33235),
            .I(N__33210));
    InMux I__6702 (
            .O(N__33232),
            .I(N__33210));
    InMux I__6701 (
            .O(N__33231),
            .I(N__33210));
    InMux I__6700 (
            .O(N__33230),
            .I(N__33210));
    InMux I__6699 (
            .O(N__33229),
            .I(N__33205));
    LocalMux I__6698 (
            .O(N__33224),
            .I(N__33201));
    LocalMux I__6697 (
            .O(N__33219),
            .I(N__33196));
    LocalMux I__6696 (
            .O(N__33210),
            .I(N__33196));
    InMux I__6695 (
            .O(N__33209),
            .I(N__33191));
    InMux I__6694 (
            .O(N__33208),
            .I(N__33191));
    LocalMux I__6693 (
            .O(N__33205),
            .I(N__33188));
    InMux I__6692 (
            .O(N__33204),
            .I(N__33185));
    Span4Mux_v I__6691 (
            .O(N__33201),
            .I(N__33182));
    Span4Mux_v I__6690 (
            .O(N__33196),
            .I(N__33178));
    LocalMux I__6689 (
            .O(N__33191),
            .I(N__33175));
    Span4Mux_v I__6688 (
            .O(N__33188),
            .I(N__33167));
    LocalMux I__6687 (
            .O(N__33185),
            .I(N__33167));
    Span4Mux_h I__6686 (
            .O(N__33182),
            .I(N__33160));
    InMux I__6685 (
            .O(N__33181),
            .I(N__33157));
    Span4Mux_v I__6684 (
            .O(N__33178),
            .I(N__33152));
    Span4Mux_v I__6683 (
            .O(N__33175),
            .I(N__33152));
    InMux I__6682 (
            .O(N__33174),
            .I(N__33147));
    InMux I__6681 (
            .O(N__33173),
            .I(N__33147));
    CascadeMux I__6680 (
            .O(N__33172),
            .I(N__33143));
    Span4Mux_h I__6679 (
            .O(N__33167),
            .I(N__33140));
    InMux I__6678 (
            .O(N__33166),
            .I(N__33131));
    InMux I__6677 (
            .O(N__33165),
            .I(N__33131));
    InMux I__6676 (
            .O(N__33164),
            .I(N__33131));
    InMux I__6675 (
            .O(N__33163),
            .I(N__33131));
    Span4Mux_v I__6674 (
            .O(N__33160),
            .I(N__33126));
    LocalMux I__6673 (
            .O(N__33157),
            .I(N__33126));
    Span4Mux_h I__6672 (
            .O(N__33152),
            .I(N__33121));
    LocalMux I__6671 (
            .O(N__33147),
            .I(N__33121));
    InMux I__6670 (
            .O(N__33146),
            .I(N__33116));
    InMux I__6669 (
            .O(N__33143),
            .I(N__33116));
    Odrv4 I__6668 (
            .O(N__33140),
            .I(\pid_alt.N_96_i ));
    LocalMux I__6667 (
            .O(N__33131),
            .I(\pid_alt.N_96_i ));
    Odrv4 I__6666 (
            .O(N__33126),
            .I(\pid_alt.N_96_i ));
    Odrv4 I__6665 (
            .O(N__33121),
            .I(\pid_alt.N_96_i ));
    LocalMux I__6664 (
            .O(N__33116),
            .I(\pid_alt.N_96_i ));
    CascadeMux I__6663 (
            .O(N__33105),
            .I(N__33102));
    InMux I__6662 (
            .O(N__33102),
            .I(N__33099));
    LocalMux I__6661 (
            .O(N__33099),
            .I(N__33094));
    InMux I__6660 (
            .O(N__33098),
            .I(N__33091));
    InMux I__6659 (
            .O(N__33097),
            .I(N__33088));
    Span4Mux_h I__6658 (
            .O(N__33094),
            .I(N__33081));
    LocalMux I__6657 (
            .O(N__33091),
            .I(N__33081));
    LocalMux I__6656 (
            .O(N__33088),
            .I(N__33081));
    Odrv4 I__6655 (
            .O(N__33081),
            .I(\pid_alt.error_i_acumm_preregZ0Z_11 ));
    InMux I__6654 (
            .O(N__33078),
            .I(N__33071));
    InMux I__6653 (
            .O(N__33077),
            .I(N__33071));
    InMux I__6652 (
            .O(N__33076),
            .I(N__33064));
    LocalMux I__6651 (
            .O(N__33071),
            .I(N__33061));
    InMux I__6650 (
            .O(N__33070),
            .I(N__33058));
    InMux I__6649 (
            .O(N__33069),
            .I(N__33051));
    InMux I__6648 (
            .O(N__33068),
            .I(N__33051));
    InMux I__6647 (
            .O(N__33067),
            .I(N__33051));
    LocalMux I__6646 (
            .O(N__33064),
            .I(N__33044));
    Span4Mux_v I__6645 (
            .O(N__33061),
            .I(N__33044));
    LocalMux I__6644 (
            .O(N__33058),
            .I(N__33039));
    LocalMux I__6643 (
            .O(N__33051),
            .I(N__33039));
    InMux I__6642 (
            .O(N__33050),
            .I(N__33034));
    InMux I__6641 (
            .O(N__33049),
            .I(N__33034));
    Odrv4 I__6640 (
            .O(N__33044),
            .I(\pid_alt.N_128 ));
    Odrv4 I__6639 (
            .O(N__33039),
            .I(\pid_alt.N_128 ));
    LocalMux I__6638 (
            .O(N__33034),
            .I(\pid_alt.N_128 ));
    InMux I__6637 (
            .O(N__33027),
            .I(N__33023));
    InMux I__6636 (
            .O(N__33026),
            .I(N__33020));
    LocalMux I__6635 (
            .O(N__33023),
            .I(\pid_alt.error_i_acummZ0Z_11 ));
    LocalMux I__6634 (
            .O(N__33020),
            .I(\pid_alt.error_i_acummZ0Z_11 ));
    InMux I__6633 (
            .O(N__33015),
            .I(N__33012));
    LocalMux I__6632 (
            .O(N__33012),
            .I(N__33008));
    InMux I__6631 (
            .O(N__33011),
            .I(N__33005));
    Span4Mux_h I__6630 (
            .O(N__33008),
            .I(N__33002));
    LocalMux I__6629 (
            .O(N__33005),
            .I(N__32999));
    Span4Mux_v I__6628 (
            .O(N__33002),
            .I(N__32996));
    Span4Mux_v I__6627 (
            .O(N__32999),
            .I(N__32993));
    Odrv4 I__6626 (
            .O(N__32996),
            .I(scaler_3_data_10));
    Odrv4 I__6625 (
            .O(N__32993),
            .I(scaler_3_data_10));
    InMux I__6624 (
            .O(N__32988),
            .I(N__32985));
    LocalMux I__6623 (
            .O(N__32985),
            .I(\ppm_encoder_1.un1_elevator_cry_9_THRU_CO ));
    CascadeMux I__6622 (
            .O(N__32982),
            .I(N__32977));
    InMux I__6621 (
            .O(N__32981),
            .I(N__32970));
    InMux I__6620 (
            .O(N__32980),
            .I(N__32970));
    InMux I__6619 (
            .O(N__32977),
            .I(N__32970));
    LocalMux I__6618 (
            .O(N__32970),
            .I(\ppm_encoder_1.elevatorZ0Z_10 ));
    InMux I__6617 (
            .O(N__32967),
            .I(N__32964));
    LocalMux I__6616 (
            .O(N__32964),
            .I(N__32961));
    Span4Mux_h I__6615 (
            .O(N__32961),
            .I(N__32957));
    InMux I__6614 (
            .O(N__32960),
            .I(N__32954));
    Odrv4 I__6613 (
            .O(N__32957),
            .I(scaler_4_data_10));
    LocalMux I__6612 (
            .O(N__32954),
            .I(scaler_4_data_10));
    InMux I__6611 (
            .O(N__32949),
            .I(N__32946));
    LocalMux I__6610 (
            .O(N__32946),
            .I(\ppm_encoder_1.un1_rudder_cry_9_THRU_CO ));
    CascadeMux I__6609 (
            .O(N__32943),
            .I(N__32939));
    InMux I__6608 (
            .O(N__32942),
            .I(N__32935));
    InMux I__6607 (
            .O(N__32939),
            .I(N__32932));
    IoInMux I__6606 (
            .O(N__32938),
            .I(N__32929));
    LocalMux I__6605 (
            .O(N__32935),
            .I(N__32923));
    LocalMux I__6604 (
            .O(N__32932),
            .I(N__32923));
    LocalMux I__6603 (
            .O(N__32929),
            .I(N__32920));
    InMux I__6602 (
            .O(N__32928),
            .I(N__32917));
    Span4Mux_h I__6601 (
            .O(N__32923),
            .I(N__32914));
    IoSpan4Mux I__6600 (
            .O(N__32920),
            .I(N__32911));
    LocalMux I__6599 (
            .O(N__32917),
            .I(N__32908));
    Span4Mux_v I__6598 (
            .O(N__32914),
            .I(N__32905));
    Span4Mux_s3_v I__6597 (
            .O(N__32911),
            .I(N__32902));
    Span4Mux_v I__6596 (
            .O(N__32908),
            .I(N__32899));
    Span4Mux_v I__6595 (
            .O(N__32905),
            .I(N__32896));
    Span4Mux_v I__6594 (
            .O(N__32902),
            .I(N__32893));
    Odrv4 I__6593 (
            .O(N__32899),
            .I(reset_system));
    Odrv4 I__6592 (
            .O(N__32896),
            .I(reset_system));
    Odrv4 I__6591 (
            .O(N__32893),
            .I(reset_system));
    IoInMux I__6590 (
            .O(N__32886),
            .I(N__32883));
    LocalMux I__6589 (
            .O(N__32883),
            .I(N__32880));
    Span4Mux_s3_v I__6588 (
            .O(N__32880),
            .I(N__32877));
    Span4Mux_v I__6587 (
            .O(N__32877),
            .I(N__32874));
    Span4Mux_v I__6586 (
            .O(N__32874),
            .I(N__32871));
    Odrv4 I__6585 (
            .O(N__32871),
            .I(\ppm_encoder_1.counter24_0_I_57_c_RNIGCOZ0Z83 ));
    InMux I__6584 (
            .O(N__32868),
            .I(N__32865));
    LocalMux I__6583 (
            .O(N__32865),
            .I(N__32862));
    Span4Mux_h I__6582 (
            .O(N__32862),
            .I(N__32859));
    Odrv4 I__6581 (
            .O(N__32859),
            .I(\ppm_encoder_1.N_145 ));
    InMux I__6580 (
            .O(N__32856),
            .I(N__32853));
    LocalMux I__6579 (
            .O(N__32853),
            .I(N__32849));
    InMux I__6578 (
            .O(N__32852),
            .I(N__32846));
    Span4Mux_v I__6577 (
            .O(N__32849),
            .I(N__32839));
    LocalMux I__6576 (
            .O(N__32846),
            .I(N__32839));
    InMux I__6575 (
            .O(N__32845),
            .I(N__32836));
    InMux I__6574 (
            .O(N__32844),
            .I(N__32833));
    Odrv4 I__6573 (
            .O(N__32839),
            .I(\pid_alt.error_i_acumm_preregZ0Z_21 ));
    LocalMux I__6572 (
            .O(N__32836),
            .I(\pid_alt.error_i_acumm_preregZ0Z_21 ));
    LocalMux I__6571 (
            .O(N__32833),
            .I(\pid_alt.error_i_acumm_preregZ0Z_21 ));
    InMux I__6570 (
            .O(N__32826),
            .I(N__32823));
    LocalMux I__6569 (
            .O(N__32823),
            .I(N__32818));
    InMux I__6568 (
            .O(N__32822),
            .I(N__32815));
    InMux I__6567 (
            .O(N__32821),
            .I(N__32812));
    Span4Mux_h I__6566 (
            .O(N__32818),
            .I(N__32805));
    LocalMux I__6565 (
            .O(N__32815),
            .I(N__32805));
    LocalMux I__6564 (
            .O(N__32812),
            .I(N__32805));
    Span4Mux_h I__6563 (
            .O(N__32805),
            .I(N__32802));
    Odrv4 I__6562 (
            .O(N__32802),
            .I(\pid_alt.error_i_acumm7lto13 ));
    InMux I__6561 (
            .O(N__32799),
            .I(N__32796));
    LocalMux I__6560 (
            .O(N__32796),
            .I(N__32792));
    InMux I__6559 (
            .O(N__32795),
            .I(N__32789));
    Odrv4 I__6558 (
            .O(N__32792),
            .I(\pid_alt.N_238 ));
    LocalMux I__6557 (
            .O(N__32789),
            .I(\pid_alt.N_238 ));
    InMux I__6556 (
            .O(N__32784),
            .I(N__32781));
    LocalMux I__6555 (
            .O(N__32781),
            .I(N__32778));
    Odrv4 I__6554 (
            .O(N__32778),
            .I(\pid_alt.error_i_acummZ0Z_13 ));
    CEMux I__6553 (
            .O(N__32775),
            .I(N__32772));
    LocalMux I__6552 (
            .O(N__32772),
            .I(N__32768));
    CEMux I__6551 (
            .O(N__32771),
            .I(N__32765));
    Span4Mux_h I__6550 (
            .O(N__32768),
            .I(N__32762));
    LocalMux I__6549 (
            .O(N__32765),
            .I(N__32759));
    Odrv4 I__6548 (
            .O(N__32762),
            .I(\pid_alt.N_96_i_0 ));
    Odrv12 I__6547 (
            .O(N__32759),
            .I(\pid_alt.N_96_i_0 ));
    InMux I__6546 (
            .O(N__32754),
            .I(N__32751));
    LocalMux I__6545 (
            .O(N__32751),
            .I(\ppm_encoder_1.un1_rudder_cry_10_THRU_CO ));
    InMux I__6544 (
            .O(N__32748),
            .I(N__32745));
    LocalMux I__6543 (
            .O(N__32745),
            .I(N__32742));
    Span4Mux_h I__6542 (
            .O(N__32742),
            .I(N__32738));
    InMux I__6541 (
            .O(N__32741),
            .I(N__32735));
    Odrv4 I__6540 (
            .O(N__32738),
            .I(scaler_4_data_11));
    LocalMux I__6539 (
            .O(N__32735),
            .I(scaler_4_data_11));
    CascadeMux I__6538 (
            .O(N__32730),
            .I(N__32727));
    InMux I__6537 (
            .O(N__32727),
            .I(N__32724));
    LocalMux I__6536 (
            .O(N__32724),
            .I(N__32720));
    InMux I__6535 (
            .O(N__32723),
            .I(N__32717));
    Span4Mux_h I__6534 (
            .O(N__32720),
            .I(N__32712));
    LocalMux I__6533 (
            .O(N__32717),
            .I(N__32712));
    Span4Mux_v I__6532 (
            .O(N__32712),
            .I(N__32709));
    Odrv4 I__6531 (
            .O(N__32709),
            .I(throttle_command_11));
    InMux I__6530 (
            .O(N__32706),
            .I(N__32703));
    LocalMux I__6529 (
            .O(N__32703),
            .I(N__32700));
    Odrv4 I__6528 (
            .O(N__32700),
            .I(\ppm_encoder_1.un1_throttle_cry_10_THRU_CO ));
    InMux I__6527 (
            .O(N__32697),
            .I(N__32693));
    InMux I__6526 (
            .O(N__32696),
            .I(N__32690));
    LocalMux I__6525 (
            .O(N__32693),
            .I(N__32687));
    LocalMux I__6524 (
            .O(N__32690),
            .I(N__32684));
    Span4Mux_v I__6523 (
            .O(N__32687),
            .I(N__32681));
    Span4Mux_v I__6522 (
            .O(N__32684),
            .I(N__32678));
    Odrv4 I__6521 (
            .O(N__32681),
            .I(scaler_3_data_11));
    Odrv4 I__6520 (
            .O(N__32678),
            .I(scaler_3_data_11));
    InMux I__6519 (
            .O(N__32673),
            .I(N__32670));
    LocalMux I__6518 (
            .O(N__32670),
            .I(N__32667));
    Span4Mux_h I__6517 (
            .O(N__32667),
            .I(N__32664));
    Odrv4 I__6516 (
            .O(N__32664),
            .I(\ppm_encoder_1.un1_elevator_cry_10_THRU_CO ));
    InMux I__6515 (
            .O(N__32661),
            .I(N__32658));
    LocalMux I__6514 (
            .O(N__32658),
            .I(N__32655));
    Span4Mux_v I__6513 (
            .O(N__32655),
            .I(N__32651));
    InMux I__6512 (
            .O(N__32654),
            .I(N__32648));
    Odrv4 I__6511 (
            .O(N__32651),
            .I(scaler_4_data_12));
    LocalMux I__6510 (
            .O(N__32648),
            .I(scaler_4_data_12));
    InMux I__6509 (
            .O(N__32643),
            .I(N__32640));
    LocalMux I__6508 (
            .O(N__32640),
            .I(\ppm_encoder_1.un1_rudder_cry_11_THRU_CO ));
    InMux I__6507 (
            .O(N__32637),
            .I(N__32630));
    InMux I__6506 (
            .O(N__32636),
            .I(N__32630));
    InMux I__6505 (
            .O(N__32635),
            .I(N__32627));
    LocalMux I__6504 (
            .O(N__32630),
            .I(\ppm_encoder_1.rudderZ0Z_12 ));
    LocalMux I__6503 (
            .O(N__32627),
            .I(\ppm_encoder_1.rudderZ0Z_12 ));
    CascadeMux I__6502 (
            .O(N__32622),
            .I(\ppm_encoder_1.N_320_cascade_ ));
    CascadeMux I__6501 (
            .O(N__32619),
            .I(N__32614));
    CascadeMux I__6500 (
            .O(N__32618),
            .I(N__32611));
    InMux I__6499 (
            .O(N__32617),
            .I(N__32606));
    InMux I__6498 (
            .O(N__32614),
            .I(N__32606));
    InMux I__6497 (
            .O(N__32611),
            .I(N__32603));
    LocalMux I__6496 (
            .O(N__32606),
            .I(N__32600));
    LocalMux I__6495 (
            .O(N__32603),
            .I(\ppm_encoder_1.throttleZ0Z_10 ));
    Odrv4 I__6494 (
            .O(N__32600),
            .I(\ppm_encoder_1.throttleZ0Z_10 ));
    InMux I__6493 (
            .O(N__32595),
            .I(N__32592));
    LocalMux I__6492 (
            .O(N__32592),
            .I(N__32589));
    Span4Mux_h I__6491 (
            .O(N__32589),
            .I(N__32585));
    InMux I__6490 (
            .O(N__32588),
            .I(N__32582));
    Odrv4 I__6489 (
            .O(N__32585),
            .I(throttle_command_9));
    LocalMux I__6488 (
            .O(N__32582),
            .I(throttle_command_9));
    InMux I__6487 (
            .O(N__32577),
            .I(N__32574));
    LocalMux I__6486 (
            .O(N__32574),
            .I(\ppm_encoder_1.un1_throttle_cry_8_THRU_CO ));
    CascadeMux I__6485 (
            .O(N__32571),
            .I(N__32566));
    InMux I__6484 (
            .O(N__32570),
            .I(N__32559));
    InMux I__6483 (
            .O(N__32569),
            .I(N__32559));
    InMux I__6482 (
            .O(N__32566),
            .I(N__32559));
    LocalMux I__6481 (
            .O(N__32559),
            .I(\ppm_encoder_1.throttleZ0Z_9 ));
    CascadeMux I__6480 (
            .O(N__32556),
            .I(\ppm_encoder_1.un2_throttle_iv_0_12_cascade_ ));
    InMux I__6479 (
            .O(N__32553),
            .I(N__32550));
    LocalMux I__6478 (
            .O(N__32550),
            .I(\ppm_encoder_1.un2_throttle_iv_1_12 ));
    CascadeMux I__6477 (
            .O(N__32547),
            .I(N__32544));
    InMux I__6476 (
            .O(N__32544),
            .I(N__32539));
    InMux I__6475 (
            .O(N__32543),
            .I(N__32534));
    InMux I__6474 (
            .O(N__32542),
            .I(N__32534));
    LocalMux I__6473 (
            .O(N__32539),
            .I(\ppm_encoder_1.aileronZ0Z_12 ));
    LocalMux I__6472 (
            .O(N__32534),
            .I(\ppm_encoder_1.aileronZ0Z_12 ));
    InMux I__6471 (
            .O(N__32529),
            .I(N__32525));
    InMux I__6470 (
            .O(N__32528),
            .I(N__32522));
    LocalMux I__6469 (
            .O(N__32525),
            .I(N__32519));
    LocalMux I__6468 (
            .O(N__32522),
            .I(N__32516));
    Span4Mux_h I__6467 (
            .O(N__32519),
            .I(N__32513));
    Span4Mux_v I__6466 (
            .O(N__32516),
            .I(N__32510));
    Odrv4 I__6465 (
            .O(N__32513),
            .I(scaler_3_data_12));
    Odrv4 I__6464 (
            .O(N__32510),
            .I(scaler_3_data_12));
    InMux I__6463 (
            .O(N__32505),
            .I(N__32502));
    LocalMux I__6462 (
            .O(N__32502),
            .I(N__32499));
    Span4Mux_h I__6461 (
            .O(N__32499),
            .I(N__32496));
    Odrv4 I__6460 (
            .O(N__32496),
            .I(\ppm_encoder_1.un1_elevator_cry_11_THRU_CO ));
    InMux I__6459 (
            .O(N__32493),
            .I(N__32489));
    InMux I__6458 (
            .O(N__32492),
            .I(N__32486));
    LocalMux I__6457 (
            .O(N__32489),
            .I(N__32483));
    LocalMux I__6456 (
            .O(N__32486),
            .I(N__32480));
    Span4Mux_h I__6455 (
            .O(N__32483),
            .I(N__32477));
    Span4Mux_h I__6454 (
            .O(N__32480),
            .I(N__32474));
    Span4Mux_h I__6453 (
            .O(N__32477),
            .I(N__32471));
    Span4Mux_h I__6452 (
            .O(N__32474),
            .I(N__32468));
    Odrv4 I__6451 (
            .O(N__32471),
            .I(throttle_command_12));
    Odrv4 I__6450 (
            .O(N__32468),
            .I(throttle_command_12));
    CascadeMux I__6449 (
            .O(N__32463),
            .I(N__32460));
    InMux I__6448 (
            .O(N__32460),
            .I(N__32457));
    LocalMux I__6447 (
            .O(N__32457),
            .I(N__32454));
    Odrv4 I__6446 (
            .O(N__32454),
            .I(\ppm_encoder_1.un1_throttle_cry_11_THRU_CO ));
    InMux I__6445 (
            .O(N__32451),
            .I(N__32447));
    InMux I__6444 (
            .O(N__32450),
            .I(N__32444));
    LocalMux I__6443 (
            .O(N__32447),
            .I(N__32441));
    LocalMux I__6442 (
            .O(N__32444),
            .I(N__32438));
    Span4Mux_h I__6441 (
            .O(N__32441),
            .I(N__32435));
    Span4Mux_h I__6440 (
            .O(N__32438),
            .I(N__32432));
    Odrv4 I__6439 (
            .O(N__32435),
            .I(\scaler_2.un3_source_data_0_cry_7_c_RNIJ0VM ));
    Odrv4 I__6438 (
            .O(N__32432),
            .I(\scaler_2.un3_source_data_0_cry_7_c_RNIJ0VM ));
    CascadeMux I__6437 (
            .O(N__32427),
            .I(N__32424));
    InMux I__6436 (
            .O(N__32424),
            .I(N__32421));
    LocalMux I__6435 (
            .O(N__32421),
            .I(N__32418));
    Span4Mux_h I__6434 (
            .O(N__32418),
            .I(N__32415));
    Odrv4 I__6433 (
            .O(N__32415),
            .I(\scaler_2.un3_source_data_0_cry_8_c_RNIQL42 ));
    InMux I__6432 (
            .O(N__32412),
            .I(bfn_14_14_0_));
    InMux I__6431 (
            .O(N__32409),
            .I(\scaler_2.un2_source_data_0_cry_9 ));
    CEMux I__6430 (
            .O(N__32406),
            .I(N__32385));
    CEMux I__6429 (
            .O(N__32405),
            .I(N__32385));
    CEMux I__6428 (
            .O(N__32404),
            .I(N__32385));
    CEMux I__6427 (
            .O(N__32403),
            .I(N__32385));
    CEMux I__6426 (
            .O(N__32402),
            .I(N__32385));
    CEMux I__6425 (
            .O(N__32401),
            .I(N__32385));
    CEMux I__6424 (
            .O(N__32400),
            .I(N__32385));
    GlobalMux I__6423 (
            .O(N__32385),
            .I(N__32382));
    gio2CtrlBuf I__6422 (
            .O(N__32382),
            .I(debug_CH3_20A_c_0_g));
    CascadeMux I__6421 (
            .O(N__32379),
            .I(\ppm_encoder_1.un2_throttle_iv_0_9_cascade_ ));
    InMux I__6420 (
            .O(N__32376),
            .I(N__32373));
    LocalMux I__6419 (
            .O(N__32373),
            .I(\ppm_encoder_1.un2_throttle_iv_1_9 ));
    CascadeMux I__6418 (
            .O(N__32370),
            .I(\ppm_encoder_1.N_301_cascade_ ));
    InMux I__6417 (
            .O(N__32367),
            .I(N__32358));
    InMux I__6416 (
            .O(N__32366),
            .I(N__32358));
    InMux I__6415 (
            .O(N__32365),
            .I(N__32358));
    LocalMux I__6414 (
            .O(N__32358),
            .I(\ppm_encoder_1.aileronZ0Z_9 ));
    CascadeMux I__6413 (
            .O(N__32355),
            .I(N__32352));
    InMux I__6412 (
            .O(N__32352),
            .I(N__32348));
    InMux I__6411 (
            .O(N__32351),
            .I(N__32345));
    LocalMux I__6410 (
            .O(N__32348),
            .I(N__32342));
    LocalMux I__6409 (
            .O(N__32345),
            .I(N__32339));
    Span4Mux_v I__6408 (
            .O(N__32342),
            .I(N__32336));
    Span4Mux_v I__6407 (
            .O(N__32339),
            .I(N__32333));
    Odrv4 I__6406 (
            .O(N__32336),
            .I(scaler_3_data_9));
    Odrv4 I__6405 (
            .O(N__32333),
            .I(scaler_3_data_9));
    InMux I__6404 (
            .O(N__32328),
            .I(N__32325));
    LocalMux I__6403 (
            .O(N__32325),
            .I(N__32322));
    Span4Mux_v I__6402 (
            .O(N__32322),
            .I(N__32319));
    Odrv4 I__6401 (
            .O(N__32319),
            .I(\ppm_encoder_1.un1_elevator_cry_8_THRU_CO ));
    CascadeMux I__6400 (
            .O(N__32316),
            .I(N__32311));
    InMux I__6399 (
            .O(N__32315),
            .I(N__32304));
    InMux I__6398 (
            .O(N__32314),
            .I(N__32304));
    InMux I__6397 (
            .O(N__32311),
            .I(N__32304));
    LocalMux I__6396 (
            .O(N__32304),
            .I(\ppm_encoder_1.elevatorZ0Z_9 ));
    CascadeMux I__6395 (
            .O(N__32301),
            .I(N__32298));
    InMux I__6394 (
            .O(N__32298),
            .I(N__32295));
    LocalMux I__6393 (
            .O(N__32295),
            .I(N__32292));
    Odrv4 I__6392 (
            .O(N__32292),
            .I(\scaler_2.un2_source_data_0_cry_1_c_RNOZ0 ));
    CascadeMux I__6391 (
            .O(N__32289),
            .I(N__32286));
    InMux I__6390 (
            .O(N__32286),
            .I(N__32279));
    InMux I__6389 (
            .O(N__32285),
            .I(N__32279));
    InMux I__6388 (
            .O(N__32284),
            .I(N__32275));
    LocalMux I__6387 (
            .O(N__32279),
            .I(N__32272));
    InMux I__6386 (
            .O(N__32278),
            .I(N__32269));
    LocalMux I__6385 (
            .O(N__32275),
            .I(N__32264));
    Span4Mux_h I__6384 (
            .O(N__32272),
            .I(N__32264));
    LocalMux I__6383 (
            .O(N__32269),
            .I(\scaler_2.un2_source_data_0 ));
    Odrv4 I__6382 (
            .O(N__32264),
            .I(\scaler_2.un2_source_data_0 ));
    InMux I__6381 (
            .O(N__32259),
            .I(\scaler_2.un2_source_data_0_cry_1 ));
    CascadeMux I__6380 (
            .O(N__32256),
            .I(N__32253));
    InMux I__6379 (
            .O(N__32253),
            .I(N__32247));
    InMux I__6378 (
            .O(N__32252),
            .I(N__32247));
    LocalMux I__6377 (
            .O(N__32247),
            .I(N__32244));
    Span4Mux_v I__6376 (
            .O(N__32244),
            .I(N__32241));
    Odrv4 I__6375 (
            .O(N__32241),
            .I(\scaler_2.un3_source_data_0_cry_1_c_RNI14IK ));
    InMux I__6374 (
            .O(N__32238),
            .I(\scaler_2.un2_source_data_0_cry_2 ));
    CascadeMux I__6373 (
            .O(N__32235),
            .I(N__32232));
    InMux I__6372 (
            .O(N__32232),
            .I(N__32226));
    InMux I__6371 (
            .O(N__32231),
            .I(N__32226));
    LocalMux I__6370 (
            .O(N__32226),
            .I(N__32223));
    Span4Mux_v I__6369 (
            .O(N__32223),
            .I(N__32220));
    Odrv4 I__6368 (
            .O(N__32220),
            .I(\scaler_2.un3_source_data_0_cry_2_c_RNI48JK ));
    InMux I__6367 (
            .O(N__32217),
            .I(\scaler_2.un2_source_data_0_cry_3 ));
    CascadeMux I__6366 (
            .O(N__32214),
            .I(N__32211));
    InMux I__6365 (
            .O(N__32211),
            .I(N__32205));
    InMux I__6364 (
            .O(N__32210),
            .I(N__32205));
    LocalMux I__6363 (
            .O(N__32205),
            .I(N__32202));
    Span4Mux_h I__6362 (
            .O(N__32202),
            .I(N__32199));
    Odrv4 I__6361 (
            .O(N__32199),
            .I(\scaler_2.un3_source_data_0_cry_3_c_RNI7CKK ));
    InMux I__6360 (
            .O(N__32196),
            .I(\scaler_2.un2_source_data_0_cry_4 ));
    CascadeMux I__6359 (
            .O(N__32193),
            .I(N__32190));
    InMux I__6358 (
            .O(N__32190),
            .I(N__32184));
    InMux I__6357 (
            .O(N__32189),
            .I(N__32184));
    LocalMux I__6356 (
            .O(N__32184),
            .I(N__32181));
    Span4Mux_h I__6355 (
            .O(N__32181),
            .I(N__32178));
    Odrv4 I__6354 (
            .O(N__32178),
            .I(\scaler_2.un3_source_data_0_cry_4_c_RNIAGLK ));
    InMux I__6353 (
            .O(N__32175),
            .I(\scaler_2.un2_source_data_0_cry_5 ));
    CascadeMux I__6352 (
            .O(N__32172),
            .I(N__32169));
    InMux I__6351 (
            .O(N__32169),
            .I(N__32163));
    InMux I__6350 (
            .O(N__32168),
            .I(N__32163));
    LocalMux I__6349 (
            .O(N__32163),
            .I(N__32160));
    Span4Mux_h I__6348 (
            .O(N__32160),
            .I(N__32157));
    Odrv4 I__6347 (
            .O(N__32157),
            .I(\scaler_2.un3_source_data_0_cry_5_c_RNIDKMK ));
    InMux I__6346 (
            .O(N__32154),
            .I(\scaler_2.un2_source_data_0_cry_6 ));
    CascadeMux I__6345 (
            .O(N__32151),
            .I(N__32148));
    InMux I__6344 (
            .O(N__32148),
            .I(N__32142));
    InMux I__6343 (
            .O(N__32147),
            .I(N__32142));
    LocalMux I__6342 (
            .O(N__32142),
            .I(N__32139));
    Span4Mux_h I__6341 (
            .O(N__32139),
            .I(N__32136));
    Odrv4 I__6340 (
            .O(N__32136),
            .I(\scaler_2.un3_source_data_0_cry_6_c_RNIIUTM ));
    InMux I__6339 (
            .O(N__32133),
            .I(\scaler_2.un2_source_data_0_cry_7 ));
    CascadeMux I__6338 (
            .O(N__32130),
            .I(N__32126));
    InMux I__6337 (
            .O(N__32129),
            .I(N__32110));
    InMux I__6336 (
            .O(N__32126),
            .I(N__32110));
    InMux I__6335 (
            .O(N__32125),
            .I(N__32110));
    InMux I__6334 (
            .O(N__32124),
            .I(N__32103));
    InMux I__6333 (
            .O(N__32123),
            .I(N__32103));
    InMux I__6332 (
            .O(N__32122),
            .I(N__32103));
    InMux I__6331 (
            .O(N__32121),
            .I(N__32096));
    InMux I__6330 (
            .O(N__32120),
            .I(N__32096));
    InMux I__6329 (
            .O(N__32119),
            .I(N__32096));
    InMux I__6328 (
            .O(N__32118),
            .I(N__32091));
    InMux I__6327 (
            .O(N__32117),
            .I(N__32091));
    LocalMux I__6326 (
            .O(N__32110),
            .I(\uart_pc.bit_CountZ0Z_0 ));
    LocalMux I__6325 (
            .O(N__32103),
            .I(\uart_pc.bit_CountZ0Z_0 ));
    LocalMux I__6324 (
            .O(N__32096),
            .I(\uart_pc.bit_CountZ0Z_0 ));
    LocalMux I__6323 (
            .O(N__32091),
            .I(\uart_pc.bit_CountZ0Z_0 ));
    CascadeMux I__6322 (
            .O(N__32082),
            .I(N__32077));
    CascadeMux I__6321 (
            .O(N__32081),
            .I(N__32068));
    InMux I__6320 (
            .O(N__32080),
            .I(N__32062));
    InMux I__6319 (
            .O(N__32077),
            .I(N__32062));
    InMux I__6318 (
            .O(N__32076),
            .I(N__32055));
    InMux I__6317 (
            .O(N__32075),
            .I(N__32055));
    InMux I__6316 (
            .O(N__32074),
            .I(N__32055));
    InMux I__6315 (
            .O(N__32073),
            .I(N__32048));
    InMux I__6314 (
            .O(N__32072),
            .I(N__32048));
    InMux I__6313 (
            .O(N__32071),
            .I(N__32048));
    InMux I__6312 (
            .O(N__32068),
            .I(N__32043));
    InMux I__6311 (
            .O(N__32067),
            .I(N__32043));
    LocalMux I__6310 (
            .O(N__32062),
            .I(\uart_pc.bit_CountZ0Z_1 ));
    LocalMux I__6309 (
            .O(N__32055),
            .I(\uart_pc.bit_CountZ0Z_1 ));
    LocalMux I__6308 (
            .O(N__32048),
            .I(\uart_pc.bit_CountZ0Z_1 ));
    LocalMux I__6307 (
            .O(N__32043),
            .I(\uart_pc.bit_CountZ0Z_1 ));
    CascadeMux I__6306 (
            .O(N__32034),
            .I(N__32026));
    InMux I__6305 (
            .O(N__32033),
            .I(N__32020));
    InMux I__6304 (
            .O(N__32032),
            .I(N__32013));
    InMux I__6303 (
            .O(N__32031),
            .I(N__32013));
    InMux I__6302 (
            .O(N__32030),
            .I(N__32013));
    InMux I__6301 (
            .O(N__32029),
            .I(N__32006));
    InMux I__6300 (
            .O(N__32026),
            .I(N__32006));
    InMux I__6299 (
            .O(N__32025),
            .I(N__32006));
    InMux I__6298 (
            .O(N__32024),
            .I(N__32001));
    InMux I__6297 (
            .O(N__32023),
            .I(N__32001));
    LocalMux I__6296 (
            .O(N__32020),
            .I(\uart_pc.bit_CountZ0Z_2 ));
    LocalMux I__6295 (
            .O(N__32013),
            .I(\uart_pc.bit_CountZ0Z_2 ));
    LocalMux I__6294 (
            .O(N__32006),
            .I(\uart_pc.bit_CountZ0Z_2 ));
    LocalMux I__6293 (
            .O(N__32001),
            .I(\uart_pc.bit_CountZ0Z_2 ));
    InMux I__6292 (
            .O(N__31992),
            .I(N__31989));
    LocalMux I__6291 (
            .O(N__31989),
            .I(N__31986));
    Span4Mux_h I__6290 (
            .O(N__31986),
            .I(N__31983));
    Odrv4 I__6289 (
            .O(N__31983),
            .I(\uart_pc.data_Auxce_0_6 ));
    CascadeMux I__6288 (
            .O(N__31980),
            .I(\ppm_encoder_1.un2_throttle_iv_1_7_cascade_ ));
    CascadeMux I__6287 (
            .O(N__31977),
            .I(\ppm_encoder_1.N_299_cascade_ ));
    CascadeMux I__6286 (
            .O(N__31974),
            .I(N__31971));
    InMux I__6285 (
            .O(N__31971),
            .I(N__31966));
    InMux I__6284 (
            .O(N__31970),
            .I(N__31961));
    InMux I__6283 (
            .O(N__31969),
            .I(N__31961));
    LocalMux I__6282 (
            .O(N__31966),
            .I(\ppm_encoder_1.aileronZ0Z_7 ));
    LocalMux I__6281 (
            .O(N__31961),
            .I(\ppm_encoder_1.aileronZ0Z_7 ));
    InMux I__6280 (
            .O(N__31956),
            .I(N__31953));
    LocalMux I__6279 (
            .O(N__31953),
            .I(N__31950));
    Span4Mux_v I__6278 (
            .O(N__31950),
            .I(N__31947));
    Odrv4 I__6277 (
            .O(N__31947),
            .I(\ppm_encoder_1.un1_elevator_cry_6_THRU_CO ));
    InMux I__6276 (
            .O(N__31944),
            .I(N__31940));
    InMux I__6275 (
            .O(N__31943),
            .I(N__31937));
    LocalMux I__6274 (
            .O(N__31940),
            .I(N__31934));
    LocalMux I__6273 (
            .O(N__31937),
            .I(N__31931));
    Span4Mux_v I__6272 (
            .O(N__31934),
            .I(N__31928));
    Span4Mux_v I__6271 (
            .O(N__31931),
            .I(N__31925));
    Odrv4 I__6270 (
            .O(N__31928),
            .I(scaler_3_data_7));
    Odrv4 I__6269 (
            .O(N__31925),
            .I(scaler_3_data_7));
    CascadeMux I__6268 (
            .O(N__31920),
            .I(N__31915));
    InMux I__6267 (
            .O(N__31919),
            .I(N__31908));
    InMux I__6266 (
            .O(N__31918),
            .I(N__31908));
    InMux I__6265 (
            .O(N__31915),
            .I(N__31908));
    LocalMux I__6264 (
            .O(N__31908),
            .I(\ppm_encoder_1.elevatorZ0Z_7 ));
    InMux I__6263 (
            .O(N__31905),
            .I(N__31902));
    LocalMux I__6262 (
            .O(N__31902),
            .I(\ppm_encoder_1.un1_throttle_cry_6_THRU_CO ));
    CascadeMux I__6261 (
            .O(N__31899),
            .I(N__31896));
    InMux I__6260 (
            .O(N__31896),
            .I(N__31893));
    LocalMux I__6259 (
            .O(N__31893),
            .I(N__31889));
    InMux I__6258 (
            .O(N__31892),
            .I(N__31886));
    Span4Mux_h I__6257 (
            .O(N__31889),
            .I(N__31883));
    LocalMux I__6256 (
            .O(N__31886),
            .I(N__31880));
    Span4Mux_h I__6255 (
            .O(N__31883),
            .I(N__31877));
    Sp12to4 I__6254 (
            .O(N__31880),
            .I(N__31874));
    Odrv4 I__6253 (
            .O(N__31877),
            .I(throttle_command_7));
    Odrv12 I__6252 (
            .O(N__31874),
            .I(throttle_command_7));
    SRMux I__6251 (
            .O(N__31869),
            .I(N__31866));
    LocalMux I__6250 (
            .O(N__31866),
            .I(N__31863));
    Span4Mux_v I__6249 (
            .O(N__31863),
            .I(N__31860));
    Span4Mux_h I__6248 (
            .O(N__31860),
            .I(N__31857));
    Odrv4 I__6247 (
            .O(N__31857),
            .I(\uart_drone.state_RNIOU0NZ0Z_4 ));
    CascadeMux I__6246 (
            .O(N__31854),
            .I(\uart_pc.CO0_cascade_ ));
    CascadeMux I__6245 (
            .O(N__31851),
            .I(N__31846));
    CascadeMux I__6244 (
            .O(N__31850),
            .I(N__31843));
    CascadeMux I__6243 (
            .O(N__31849),
            .I(N__31839));
    InMux I__6242 (
            .O(N__31846),
            .I(N__31836));
    InMux I__6241 (
            .O(N__31843),
            .I(N__31829));
    InMux I__6240 (
            .O(N__31842),
            .I(N__31829));
    InMux I__6239 (
            .O(N__31839),
            .I(N__31829));
    LocalMux I__6238 (
            .O(N__31836),
            .I(N__31825));
    LocalMux I__6237 (
            .O(N__31829),
            .I(N__31822));
    InMux I__6236 (
            .O(N__31828),
            .I(N__31819));
    Span4Mux_v I__6235 (
            .O(N__31825),
            .I(N__31814));
    Span4Mux_h I__6234 (
            .O(N__31822),
            .I(N__31814));
    LocalMux I__6233 (
            .O(N__31819),
            .I(N__31811));
    Span4Mux_v I__6232 (
            .O(N__31814),
            .I(N__31807));
    Span4Mux_h I__6231 (
            .O(N__31811),
            .I(N__31804));
    InMux I__6230 (
            .O(N__31810),
            .I(N__31801));
    Span4Mux_v I__6229 (
            .O(N__31807),
            .I(N__31796));
    Span4Mux_h I__6228 (
            .O(N__31804),
            .I(N__31796));
    LocalMux I__6227 (
            .O(N__31801),
            .I(\Commands_frame_decoder.un1_sink_data_valid_2_0 ));
    Odrv4 I__6226 (
            .O(N__31796),
            .I(\Commands_frame_decoder.un1_sink_data_valid_2_0 ));
    CEMux I__6225 (
            .O(N__31791),
            .I(N__31788));
    LocalMux I__6224 (
            .O(N__31788),
            .I(N__31785));
    Span4Mux_h I__6223 (
            .O(N__31785),
            .I(N__31782));
    Sp12to4 I__6222 (
            .O(N__31782),
            .I(N__31779));
    Span12Mux_v I__6221 (
            .O(N__31779),
            .I(N__31776));
    Odrv12 I__6220 (
            .O(N__31776),
            .I(\Commands_frame_decoder.un1_sink_data_valid_2_0_0 ));
    InMux I__6219 (
            .O(N__31773),
            .I(N__31769));
    InMux I__6218 (
            .O(N__31772),
            .I(N__31765));
    LocalMux I__6217 (
            .O(N__31769),
            .I(N__31762));
    InMux I__6216 (
            .O(N__31768),
            .I(N__31759));
    LocalMux I__6215 (
            .O(N__31765),
            .I(N__31754));
    Span4Mux_h I__6214 (
            .O(N__31762),
            .I(N__31754));
    LocalMux I__6213 (
            .O(N__31759),
            .I(\uart_pc.N_152 ));
    Odrv4 I__6212 (
            .O(N__31754),
            .I(\uart_pc.N_152 ));
    InMux I__6211 (
            .O(N__31749),
            .I(N__31739));
    InMux I__6210 (
            .O(N__31748),
            .I(N__31739));
    InMux I__6209 (
            .O(N__31747),
            .I(N__31739));
    InMux I__6208 (
            .O(N__31746),
            .I(N__31736));
    LocalMux I__6207 (
            .O(N__31739),
            .I(N__31731));
    LocalMux I__6206 (
            .O(N__31736),
            .I(N__31731));
    Odrv4 I__6205 (
            .O(N__31731),
            .I(\uart_pc.un1_state_4_0 ));
    CascadeMux I__6204 (
            .O(N__31728),
            .I(\uart_pc.N_152_cascade_ ));
    InMux I__6203 (
            .O(N__31725),
            .I(N__31718));
    InMux I__6202 (
            .O(N__31724),
            .I(N__31715));
    InMux I__6201 (
            .O(N__31723),
            .I(N__31712));
    InMux I__6200 (
            .O(N__31722),
            .I(N__31704));
    InMux I__6199 (
            .O(N__31721),
            .I(N__31704));
    LocalMux I__6198 (
            .O(N__31718),
            .I(N__31699));
    LocalMux I__6197 (
            .O(N__31715),
            .I(N__31699));
    LocalMux I__6196 (
            .O(N__31712),
            .I(N__31696));
    InMux I__6195 (
            .O(N__31711),
            .I(N__31693));
    InMux I__6194 (
            .O(N__31710),
            .I(N__31688));
    InMux I__6193 (
            .O(N__31709),
            .I(N__31688));
    LocalMux I__6192 (
            .O(N__31704),
            .I(N__31683));
    Span4Mux_v I__6191 (
            .O(N__31699),
            .I(N__31683));
    Span4Mux_h I__6190 (
            .O(N__31696),
            .I(N__31680));
    LocalMux I__6189 (
            .O(N__31693),
            .I(\uart_pc.stateZ0Z_3 ));
    LocalMux I__6188 (
            .O(N__31688),
            .I(\uart_pc.stateZ0Z_3 ));
    Odrv4 I__6187 (
            .O(N__31683),
            .I(\uart_pc.stateZ0Z_3 ));
    Odrv4 I__6186 (
            .O(N__31680),
            .I(\uart_pc.stateZ0Z_3 ));
    InMux I__6185 (
            .O(N__31671),
            .I(N__31665));
    InMux I__6184 (
            .O(N__31670),
            .I(N__31665));
    LocalMux I__6183 (
            .O(N__31665),
            .I(N__31662));
    Odrv4 I__6182 (
            .O(N__31662),
            .I(\uart_pc.un1_state_7_0 ));
    InMux I__6181 (
            .O(N__31659),
            .I(N__31655));
    InMux I__6180 (
            .O(N__31658),
            .I(N__31652));
    LocalMux I__6179 (
            .O(N__31655),
            .I(\uart_drone.stateZ0Z_0 ));
    LocalMux I__6178 (
            .O(N__31652),
            .I(\uart_drone.stateZ0Z_0 ));
    InMux I__6177 (
            .O(N__31647),
            .I(N__31644));
    LocalMux I__6176 (
            .O(N__31644),
            .I(N__31639));
    InMux I__6175 (
            .O(N__31643),
            .I(N__31634));
    InMux I__6174 (
            .O(N__31642),
            .I(N__31634));
    Span4Mux_v I__6173 (
            .O(N__31639),
            .I(N__31631));
    LocalMux I__6172 (
            .O(N__31634),
            .I(N__31628));
    Span4Mux_h I__6171 (
            .O(N__31631),
            .I(N__31623));
    Span4Mux_v I__6170 (
            .O(N__31628),
            .I(N__31623));
    Odrv4 I__6169 (
            .O(N__31623),
            .I(\uart_drone.data_rdyc_1 ));
    InMux I__6168 (
            .O(N__31620),
            .I(N__31616));
    InMux I__6167 (
            .O(N__31619),
            .I(N__31612));
    LocalMux I__6166 (
            .O(N__31616),
            .I(N__31608));
    CascadeMux I__6165 (
            .O(N__31615),
            .I(N__31602));
    LocalMux I__6164 (
            .O(N__31612),
            .I(N__31598));
    InMux I__6163 (
            .O(N__31611),
            .I(N__31595));
    Span4Mux_v I__6162 (
            .O(N__31608),
            .I(N__31592));
    InMux I__6161 (
            .O(N__31607),
            .I(N__31589));
    InMux I__6160 (
            .O(N__31606),
            .I(N__31584));
    InMux I__6159 (
            .O(N__31605),
            .I(N__31584));
    InMux I__6158 (
            .O(N__31602),
            .I(N__31579));
    InMux I__6157 (
            .O(N__31601),
            .I(N__31579));
    Span4Mux_h I__6156 (
            .O(N__31598),
            .I(N__31576));
    LocalMux I__6155 (
            .O(N__31595),
            .I(\uart_pc.timer_CountZ1Z_3 ));
    Odrv4 I__6154 (
            .O(N__31592),
            .I(\uart_pc.timer_CountZ1Z_3 ));
    LocalMux I__6153 (
            .O(N__31589),
            .I(\uart_pc.timer_CountZ1Z_3 ));
    LocalMux I__6152 (
            .O(N__31584),
            .I(\uart_pc.timer_CountZ1Z_3 ));
    LocalMux I__6151 (
            .O(N__31579),
            .I(\uart_pc.timer_CountZ1Z_3 ));
    Odrv4 I__6150 (
            .O(N__31576),
            .I(\uart_pc.timer_CountZ1Z_3 ));
    InMux I__6149 (
            .O(N__31563),
            .I(N__31559));
    InMux I__6148 (
            .O(N__31562),
            .I(N__31556));
    LocalMux I__6147 (
            .O(N__31559),
            .I(N__31551));
    LocalMux I__6146 (
            .O(N__31556),
            .I(N__31548));
    InMux I__6145 (
            .O(N__31555),
            .I(N__31543));
    InMux I__6144 (
            .O(N__31554),
            .I(N__31540));
    Span4Mux_h I__6143 (
            .O(N__31551),
            .I(N__31535));
    Span4Mux_h I__6142 (
            .O(N__31548),
            .I(N__31535));
    InMux I__6141 (
            .O(N__31547),
            .I(N__31530));
    InMux I__6140 (
            .O(N__31546),
            .I(N__31530));
    LocalMux I__6139 (
            .O(N__31543),
            .I(\uart_pc.stateZ0Z_4 ));
    LocalMux I__6138 (
            .O(N__31540),
            .I(\uart_pc.stateZ0Z_4 ));
    Odrv4 I__6137 (
            .O(N__31535),
            .I(\uart_pc.stateZ0Z_4 ));
    LocalMux I__6136 (
            .O(N__31530),
            .I(\uart_pc.stateZ0Z_4 ));
    CascadeMux I__6135 (
            .O(N__31521),
            .I(N__31516));
    InMux I__6134 (
            .O(N__31520),
            .I(N__31513));
    InMux I__6133 (
            .O(N__31519),
            .I(N__31510));
    InMux I__6132 (
            .O(N__31516),
            .I(N__31506));
    LocalMux I__6131 (
            .O(N__31513),
            .I(N__31500));
    LocalMux I__6130 (
            .O(N__31510),
            .I(N__31497));
    InMux I__6129 (
            .O(N__31509),
            .I(N__31494));
    LocalMux I__6128 (
            .O(N__31506),
            .I(N__31491));
    CascadeMux I__6127 (
            .O(N__31505),
            .I(N__31486));
    InMux I__6126 (
            .O(N__31504),
            .I(N__31483));
    InMux I__6125 (
            .O(N__31503),
            .I(N__31480));
    Span4Mux_v I__6124 (
            .O(N__31500),
            .I(N__31473));
    Span4Mux_h I__6123 (
            .O(N__31497),
            .I(N__31473));
    LocalMux I__6122 (
            .O(N__31494),
            .I(N__31473));
    Span4Mux_h I__6121 (
            .O(N__31491),
            .I(N__31470));
    InMux I__6120 (
            .O(N__31490),
            .I(N__31463));
    InMux I__6119 (
            .O(N__31489),
            .I(N__31463));
    InMux I__6118 (
            .O(N__31486),
            .I(N__31463));
    LocalMux I__6117 (
            .O(N__31483),
            .I(\uart_pc.timer_CountZ0Z_4 ));
    LocalMux I__6116 (
            .O(N__31480),
            .I(\uart_pc.timer_CountZ0Z_4 ));
    Odrv4 I__6115 (
            .O(N__31473),
            .I(\uart_pc.timer_CountZ0Z_4 ));
    Odrv4 I__6114 (
            .O(N__31470),
            .I(\uart_pc.timer_CountZ0Z_4 ));
    LocalMux I__6113 (
            .O(N__31463),
            .I(\uart_pc.timer_CountZ0Z_4 ));
    CascadeMux I__6112 (
            .O(N__31452),
            .I(N__31449));
    InMux I__6111 (
            .O(N__31449),
            .I(N__31445));
    InMux I__6110 (
            .O(N__31448),
            .I(N__31442));
    LocalMux I__6109 (
            .O(N__31445),
            .I(\uart_drone.N_126_li ));
    LocalMux I__6108 (
            .O(N__31442),
            .I(\uart_drone.N_126_li ));
    InMux I__6107 (
            .O(N__31437),
            .I(N__31413));
    InMux I__6106 (
            .O(N__31436),
            .I(N__31413));
    InMux I__6105 (
            .O(N__31435),
            .I(N__31413));
    InMux I__6104 (
            .O(N__31434),
            .I(N__31413));
    InMux I__6103 (
            .O(N__31433),
            .I(N__31413));
    InMux I__6102 (
            .O(N__31432),
            .I(N__31413));
    InMux I__6101 (
            .O(N__31431),
            .I(N__31413));
    InMux I__6100 (
            .O(N__31430),
            .I(N__31413));
    LocalMux I__6099 (
            .O(N__31413),
            .I(N__31410));
    Span4Mux_h I__6098 (
            .O(N__31410),
            .I(N__31407));
    Odrv4 I__6097 (
            .O(N__31407),
            .I(\uart_drone.un1_state_2_0 ));
    IoInMux I__6096 (
            .O(N__31404),
            .I(N__31401));
    LocalMux I__6095 (
            .O(N__31401),
            .I(N__31398));
    IoSpan4Mux I__6094 (
            .O(N__31398),
            .I(N__31394));
    CascadeMux I__6093 (
            .O(N__31397),
            .I(N__31385));
    Span4Mux_s1_v I__6092 (
            .O(N__31394),
            .I(N__31379));
    InMux I__6091 (
            .O(N__31393),
            .I(N__31376));
    InMux I__6090 (
            .O(N__31392),
            .I(N__31373));
    InMux I__6089 (
            .O(N__31391),
            .I(N__31359));
    InMux I__6088 (
            .O(N__31390),
            .I(N__31359));
    InMux I__6087 (
            .O(N__31389),
            .I(N__31359));
    InMux I__6086 (
            .O(N__31388),
            .I(N__31359));
    InMux I__6085 (
            .O(N__31385),
            .I(N__31359));
    InMux I__6084 (
            .O(N__31384),
            .I(N__31352));
    InMux I__6083 (
            .O(N__31383),
            .I(N__31352));
    InMux I__6082 (
            .O(N__31382),
            .I(N__31352));
    Span4Mux_v I__6081 (
            .O(N__31379),
            .I(N__31345));
    LocalMux I__6080 (
            .O(N__31376),
            .I(N__31345));
    LocalMux I__6079 (
            .O(N__31373),
            .I(N__31345));
    InMux I__6078 (
            .O(N__31372),
            .I(N__31342));
    InMux I__6077 (
            .O(N__31371),
            .I(N__31339));
    InMux I__6076 (
            .O(N__31370),
            .I(N__31336));
    LocalMux I__6075 (
            .O(N__31359),
            .I(N__31331));
    LocalMux I__6074 (
            .O(N__31352),
            .I(N__31331));
    Span4Mux_v I__6073 (
            .O(N__31345),
            .I(N__31326));
    LocalMux I__6072 (
            .O(N__31342),
            .I(N__31326));
    LocalMux I__6071 (
            .O(N__31339),
            .I(N__31323));
    LocalMux I__6070 (
            .O(N__31336),
            .I(N__31320));
    Span4Mux_v I__6069 (
            .O(N__31331),
            .I(N__31315));
    Span4Mux_h I__6068 (
            .O(N__31326),
            .I(N__31315));
    Span4Mux_v I__6067 (
            .O(N__31323),
            .I(N__31310));
    Span4Mux_h I__6066 (
            .O(N__31320),
            .I(N__31310));
    Odrv4 I__6065 (
            .O(N__31315),
            .I(debug_CH0_16A_c));
    Odrv4 I__6064 (
            .O(N__31310),
            .I(debug_CH0_16A_c));
    CascadeMux I__6063 (
            .O(N__31305),
            .I(\uart_drone.state_srsts_i_0_2_cascade_ ));
    CascadeMux I__6062 (
            .O(N__31302),
            .I(N__31297));
    CascadeMux I__6061 (
            .O(N__31301),
            .I(N__31294));
    InMux I__6060 (
            .O(N__31300),
            .I(N__31289));
    InMux I__6059 (
            .O(N__31297),
            .I(N__31289));
    InMux I__6058 (
            .O(N__31294),
            .I(N__31286));
    LocalMux I__6057 (
            .O(N__31289),
            .I(N__31283));
    LocalMux I__6056 (
            .O(N__31286),
            .I(\uart_drone.stateZ0Z_1 ));
    Odrv4 I__6055 (
            .O(N__31283),
            .I(\uart_drone.stateZ0Z_1 ));
    InMux I__6054 (
            .O(N__31278),
            .I(N__31275));
    LocalMux I__6053 (
            .O(N__31275),
            .I(N__31272));
    Span4Mux_h I__6052 (
            .O(N__31272),
            .I(N__31268));
    InMux I__6051 (
            .O(N__31271),
            .I(N__31265));
    Odrv4 I__6050 (
            .O(N__31268),
            .I(\uart_pc.N_126_li ));
    LocalMux I__6049 (
            .O(N__31265),
            .I(\uart_pc.N_126_li ));
    CascadeMux I__6048 (
            .O(N__31260),
            .I(\uart_pc.state_srsts_0_0_0_cascade_ ));
    InMux I__6047 (
            .O(N__31257),
            .I(N__31254));
    LocalMux I__6046 (
            .O(N__31254),
            .I(\uart_drone.state_srsts_0_0_0 ));
    CascadeMux I__6045 (
            .O(N__31251),
            .I(N__31248));
    InMux I__6044 (
            .O(N__31248),
            .I(N__31245));
    LocalMux I__6043 (
            .O(N__31245),
            .I(N__31241));
    InMux I__6042 (
            .O(N__31244),
            .I(N__31238));
    Odrv4 I__6041 (
            .O(N__31241),
            .I(\uart_pc.stateZ0Z_0 ));
    LocalMux I__6040 (
            .O(N__31238),
            .I(\uart_pc.stateZ0Z_0 ));
    CascadeMux I__6039 (
            .O(N__31233),
            .I(\uart_drone.N_126_li_cascade_ ));
    InMux I__6038 (
            .O(N__31230),
            .I(N__31217));
    IoInMux I__6037 (
            .O(N__31229),
            .I(N__31213));
    InMux I__6036 (
            .O(N__31228),
            .I(N__31209));
    InMux I__6035 (
            .O(N__31227),
            .I(N__31200));
    InMux I__6034 (
            .O(N__31226),
            .I(N__31200));
    InMux I__6033 (
            .O(N__31225),
            .I(N__31200));
    InMux I__6032 (
            .O(N__31224),
            .I(N__31200));
    InMux I__6031 (
            .O(N__31223),
            .I(N__31191));
    InMux I__6030 (
            .O(N__31222),
            .I(N__31191));
    InMux I__6029 (
            .O(N__31221),
            .I(N__31191));
    InMux I__6028 (
            .O(N__31220),
            .I(N__31191));
    LocalMux I__6027 (
            .O(N__31217),
            .I(N__31188));
    InMux I__6026 (
            .O(N__31216),
            .I(N__31185));
    LocalMux I__6025 (
            .O(N__31213),
            .I(N__31182));
    InMux I__6024 (
            .O(N__31212),
            .I(N__31179));
    LocalMux I__6023 (
            .O(N__31209),
            .I(N__31175));
    LocalMux I__6022 (
            .O(N__31200),
            .I(N__31170));
    LocalMux I__6021 (
            .O(N__31191),
            .I(N__31170));
    Span4Mux_v I__6020 (
            .O(N__31188),
            .I(N__31165));
    LocalMux I__6019 (
            .O(N__31185),
            .I(N__31165));
    Span4Mux_s2_v I__6018 (
            .O(N__31182),
            .I(N__31162));
    LocalMux I__6017 (
            .O(N__31179),
            .I(N__31159));
    InMux I__6016 (
            .O(N__31178),
            .I(N__31156));
    Span4Mux_v I__6015 (
            .O(N__31175),
            .I(N__31149));
    Span4Mux_h I__6014 (
            .O(N__31170),
            .I(N__31149));
    Span4Mux_h I__6013 (
            .O(N__31165),
            .I(N__31149));
    Span4Mux_h I__6012 (
            .O(N__31162),
            .I(N__31144));
    Span4Mux_h I__6011 (
            .O(N__31159),
            .I(N__31144));
    LocalMux I__6010 (
            .O(N__31156),
            .I(N__31141));
    Odrv4 I__6009 (
            .O(N__31149),
            .I(debug_CH2_18A_c));
    Odrv4 I__6008 (
            .O(N__31144),
            .I(debug_CH2_18A_c));
    Odrv12 I__6007 (
            .O(N__31141),
            .I(debug_CH2_18A_c));
    CascadeMux I__6006 (
            .O(N__31134),
            .I(\uart_pc.state_srsts_i_0_2_cascade_ ));
    CascadeMux I__6005 (
            .O(N__31131),
            .I(N__31126));
    InMux I__6004 (
            .O(N__31130),
            .I(N__31123));
    InMux I__6003 (
            .O(N__31129),
            .I(N__31118));
    InMux I__6002 (
            .O(N__31126),
            .I(N__31118));
    LocalMux I__6001 (
            .O(N__31123),
            .I(\uart_pc.stateZ0Z_1 ));
    LocalMux I__6000 (
            .O(N__31118),
            .I(\uart_pc.stateZ0Z_1 ));
    CascadeMux I__5999 (
            .O(N__31113),
            .I(N__31109));
    CascadeMux I__5998 (
            .O(N__31112),
            .I(N__31105));
    InMux I__5997 (
            .O(N__31109),
            .I(N__31102));
    InMux I__5996 (
            .O(N__31108),
            .I(N__31098));
    InMux I__5995 (
            .O(N__31105),
            .I(N__31095));
    LocalMux I__5994 (
            .O(N__31102),
            .I(N__31092));
    InMux I__5993 (
            .O(N__31101),
            .I(N__31089));
    LocalMux I__5992 (
            .O(N__31098),
            .I(N__31084));
    LocalMux I__5991 (
            .O(N__31095),
            .I(N__31084));
    Span4Mux_h I__5990 (
            .O(N__31092),
            .I(N__31081));
    LocalMux I__5989 (
            .O(N__31089),
            .I(\uart_pc.stateZ0Z_2 ));
    Odrv4 I__5988 (
            .O(N__31084),
            .I(\uart_pc.stateZ0Z_2 ));
    Odrv4 I__5987 (
            .O(N__31081),
            .I(\uart_pc.stateZ0Z_2 ));
    CascadeMux I__5986 (
            .O(N__31074),
            .I(N__31069));
    InMux I__5985 (
            .O(N__31073),
            .I(N__31064));
    InMux I__5984 (
            .O(N__31072),
            .I(N__31061));
    InMux I__5983 (
            .O(N__31069),
            .I(N__31053));
    InMux I__5982 (
            .O(N__31068),
            .I(N__31053));
    InMux I__5981 (
            .O(N__31067),
            .I(N__31053));
    LocalMux I__5980 (
            .O(N__31064),
            .I(N__31047));
    LocalMux I__5979 (
            .O(N__31061),
            .I(N__31047));
    InMux I__5978 (
            .O(N__31060),
            .I(N__31044));
    LocalMux I__5977 (
            .O(N__31053),
            .I(N__31040));
    InMux I__5976 (
            .O(N__31052),
            .I(N__31037));
    Span4Mux_h I__5975 (
            .O(N__31047),
            .I(N__31032));
    LocalMux I__5974 (
            .O(N__31044),
            .I(N__31032));
    InMux I__5973 (
            .O(N__31043),
            .I(N__31029));
    Odrv4 I__5972 (
            .O(N__31040),
            .I(\uart_pc.timer_Count_RNILR1B2Z0Z_2 ));
    LocalMux I__5971 (
            .O(N__31037),
            .I(\uart_pc.timer_Count_RNILR1B2Z0Z_2 ));
    Odrv4 I__5970 (
            .O(N__31032),
            .I(\uart_pc.timer_Count_RNILR1B2Z0Z_2 ));
    LocalMux I__5969 (
            .O(N__31029),
            .I(\uart_pc.timer_Count_RNILR1B2Z0Z_2 ));
    CascadeMux I__5968 (
            .O(N__31020),
            .I(N__31016));
    CascadeMux I__5967 (
            .O(N__31019),
            .I(N__31013));
    InMux I__5966 (
            .O(N__31016),
            .I(N__31010));
    InMux I__5965 (
            .O(N__31013),
            .I(N__31007));
    LocalMux I__5964 (
            .O(N__31010),
            .I(\uart_pc.data_AuxZ0Z_3 ));
    LocalMux I__5963 (
            .O(N__31007),
            .I(\uart_pc.data_AuxZ0Z_3 ));
    InMux I__5962 (
            .O(N__31002),
            .I(N__30996));
    CascadeMux I__5961 (
            .O(N__31001),
            .I(N__30993));
    InMux I__5960 (
            .O(N__31000),
            .I(N__30987));
    InMux I__5959 (
            .O(N__30999),
            .I(N__30984));
    LocalMux I__5958 (
            .O(N__30996),
            .I(N__30981));
    InMux I__5957 (
            .O(N__30993),
            .I(N__30978));
    InMux I__5956 (
            .O(N__30992),
            .I(N__30975));
    InMux I__5955 (
            .O(N__30991),
            .I(N__30970));
    InMux I__5954 (
            .O(N__30990),
            .I(N__30970));
    LocalMux I__5953 (
            .O(N__30987),
            .I(N__30967));
    LocalMux I__5952 (
            .O(N__30984),
            .I(N__30962));
    Span4Mux_h I__5951 (
            .O(N__30981),
            .I(N__30962));
    LocalMux I__5950 (
            .O(N__30978),
            .I(\uart_pc.timer_Count_RNIMQ8T1Z0Z_2 ));
    LocalMux I__5949 (
            .O(N__30975),
            .I(\uart_pc.timer_Count_RNIMQ8T1Z0Z_2 ));
    LocalMux I__5948 (
            .O(N__30970),
            .I(\uart_pc.timer_Count_RNIMQ8T1Z0Z_2 ));
    Odrv4 I__5947 (
            .O(N__30967),
            .I(\uart_pc.timer_Count_RNIMQ8T1Z0Z_2 ));
    Odrv4 I__5946 (
            .O(N__30962),
            .I(\uart_pc.timer_Count_RNIMQ8T1Z0Z_2 ));
    InMux I__5945 (
            .O(N__30951),
            .I(N__30945));
    InMux I__5944 (
            .O(N__30950),
            .I(N__30945));
    LocalMux I__5943 (
            .O(N__30945),
            .I(N__30941));
    InMux I__5942 (
            .O(N__30944),
            .I(N__30938));
    Span4Mux_h I__5941 (
            .O(N__30941),
            .I(N__30935));
    LocalMux I__5940 (
            .O(N__30938),
            .I(N__30932));
    Span4Mux_v I__5939 (
            .O(N__30935),
            .I(N__30929));
    Span4Mux_h I__5938 (
            .O(N__30932),
            .I(N__30926));
    Span4Mux_h I__5937 (
            .O(N__30929),
            .I(N__30923));
    Odrv4 I__5936 (
            .O(N__30926),
            .I(\pid_alt.error_i_reg_esr_RNI38LJZ0Z_15 ));
    Odrv4 I__5935 (
            .O(N__30923),
            .I(\pid_alt.error_i_reg_esr_RNI38LJZ0Z_15 ));
    InMux I__5934 (
            .O(N__30918),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_14 ));
    InMux I__5933 (
            .O(N__30915),
            .I(N__30908));
    InMux I__5932 (
            .O(N__30914),
            .I(N__30908));
    InMux I__5931 (
            .O(N__30913),
            .I(N__30905));
    LocalMux I__5930 (
            .O(N__30908),
            .I(N__30902));
    LocalMux I__5929 (
            .O(N__30905),
            .I(N__30899));
    Span4Mux_h I__5928 (
            .O(N__30902),
            .I(N__30896));
    Span4Mux_h I__5927 (
            .O(N__30899),
            .I(N__30891));
    Span4Mux_h I__5926 (
            .O(N__30896),
            .I(N__30891));
    Sp12to4 I__5925 (
            .O(N__30891),
            .I(N__30888));
    Odrv12 I__5924 (
            .O(N__30888),
            .I(\pid_alt.error_i_reg_esr_RNI5BMJZ0Z_16 ));
    InMux I__5923 (
            .O(N__30885),
            .I(bfn_13_23_0_));
    InMux I__5922 (
            .O(N__30882),
            .I(N__30876));
    InMux I__5921 (
            .O(N__30881),
            .I(N__30876));
    LocalMux I__5920 (
            .O(N__30876),
            .I(N__30872));
    InMux I__5919 (
            .O(N__30875),
            .I(N__30869));
    Span4Mux_h I__5918 (
            .O(N__30872),
            .I(N__30866));
    LocalMux I__5917 (
            .O(N__30869),
            .I(N__30863));
    Span4Mux_v I__5916 (
            .O(N__30866),
            .I(N__30860));
    Span4Mux_h I__5915 (
            .O(N__30863),
            .I(N__30857));
    Span4Mux_h I__5914 (
            .O(N__30860),
            .I(N__30854));
    Odrv4 I__5913 (
            .O(N__30857),
            .I(\pid_alt.error_i_reg_esr_RNI7ENJZ0Z_17 ));
    Odrv4 I__5912 (
            .O(N__30854),
            .I(\pid_alt.error_i_reg_esr_RNI7ENJZ0Z_17 ));
    InMux I__5911 (
            .O(N__30849),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_16 ));
    InMux I__5910 (
            .O(N__30846),
            .I(N__30840));
    InMux I__5909 (
            .O(N__30845),
            .I(N__30840));
    LocalMux I__5908 (
            .O(N__30840),
            .I(N__30836));
    InMux I__5907 (
            .O(N__30839),
            .I(N__30833));
    Span4Mux_h I__5906 (
            .O(N__30836),
            .I(N__30830));
    LocalMux I__5905 (
            .O(N__30833),
            .I(N__30827));
    Sp12to4 I__5904 (
            .O(N__30830),
            .I(N__30824));
    Span4Mux_h I__5903 (
            .O(N__30827),
            .I(N__30821));
    Span12Mux_v I__5902 (
            .O(N__30824),
            .I(N__30818));
    Odrv4 I__5901 (
            .O(N__30821),
            .I(\pid_alt.error_i_reg_esr_RNI9HOJZ0Z_18 ));
    Odrv12 I__5900 (
            .O(N__30818),
            .I(\pid_alt.error_i_reg_esr_RNI9HOJZ0Z_18 ));
    InMux I__5899 (
            .O(N__30813),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_17 ));
    InMux I__5898 (
            .O(N__30810),
            .I(N__30804));
    InMux I__5897 (
            .O(N__30809),
            .I(N__30804));
    LocalMux I__5896 (
            .O(N__30804),
            .I(N__30801));
    Span4Mux_h I__5895 (
            .O(N__30801),
            .I(N__30797));
    InMux I__5894 (
            .O(N__30800),
            .I(N__30794));
    Span4Mux_v I__5893 (
            .O(N__30797),
            .I(N__30791));
    LocalMux I__5892 (
            .O(N__30794),
            .I(N__30788));
    Span4Mux_h I__5891 (
            .O(N__30791),
            .I(N__30785));
    Span4Mux_h I__5890 (
            .O(N__30788),
            .I(N__30782));
    Span4Mux_h I__5889 (
            .O(N__30785),
            .I(N__30779));
    Odrv4 I__5888 (
            .O(N__30782),
            .I(\pid_alt.error_i_reg_esr_RNIBKPJZ0Z_19 ));
    Odrv4 I__5887 (
            .O(N__30779),
            .I(\pid_alt.error_i_reg_esr_RNIBKPJZ0Z_19 ));
    InMux I__5886 (
            .O(N__30774),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_18 ));
    InMux I__5885 (
            .O(N__30771),
            .I(N__30767));
    InMux I__5884 (
            .O(N__30770),
            .I(N__30763));
    LocalMux I__5883 (
            .O(N__30767),
            .I(N__30760));
    InMux I__5882 (
            .O(N__30766),
            .I(N__30757));
    LocalMux I__5881 (
            .O(N__30763),
            .I(N__30754));
    Span4Mux_h I__5880 (
            .O(N__30760),
            .I(N__30751));
    LocalMux I__5879 (
            .O(N__30757),
            .I(N__30748));
    Span4Mux_v I__5878 (
            .O(N__30754),
            .I(N__30745));
    Sp12to4 I__5877 (
            .O(N__30751),
            .I(N__30742));
    Span4Mux_h I__5876 (
            .O(N__30748),
            .I(N__30739));
    Span4Mux_h I__5875 (
            .O(N__30745),
            .I(N__30736));
    Span12Mux_v I__5874 (
            .O(N__30742),
            .I(N__30733));
    Odrv4 I__5873 (
            .O(N__30739),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_19_c_RNI4FRJ ));
    Odrv4 I__5872 (
            .O(N__30736),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_19_c_RNI4FRJ ));
    Odrv12 I__5871 (
            .O(N__30733),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_19_c_RNI4FRJ ));
    InMux I__5870 (
            .O(N__30726),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_19 ));
    InMux I__5869 (
            .O(N__30723),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_20 ));
    InMux I__5868 (
            .O(N__30720),
            .I(N__30714));
    InMux I__5867 (
            .O(N__30719),
            .I(N__30707));
    InMux I__5866 (
            .O(N__30718),
            .I(N__30707));
    InMux I__5865 (
            .O(N__30717),
            .I(N__30707));
    LocalMux I__5864 (
            .O(N__30714),
            .I(N__30691));
    LocalMux I__5863 (
            .O(N__30707),
            .I(N__30687));
    InMux I__5862 (
            .O(N__30706),
            .I(N__30684));
    InMux I__5861 (
            .O(N__30705),
            .I(N__30681));
    InMux I__5860 (
            .O(N__30704),
            .I(N__30676));
    InMux I__5859 (
            .O(N__30703),
            .I(N__30676));
    InMux I__5858 (
            .O(N__30702),
            .I(N__30667));
    InMux I__5857 (
            .O(N__30701),
            .I(N__30667));
    InMux I__5856 (
            .O(N__30700),
            .I(N__30667));
    InMux I__5855 (
            .O(N__30699),
            .I(N__30667));
    InMux I__5854 (
            .O(N__30698),
            .I(N__30664));
    InMux I__5853 (
            .O(N__30697),
            .I(N__30655));
    InMux I__5852 (
            .O(N__30696),
            .I(N__30655));
    InMux I__5851 (
            .O(N__30695),
            .I(N__30655));
    InMux I__5850 (
            .O(N__30694),
            .I(N__30655));
    Span4Mux_v I__5849 (
            .O(N__30691),
            .I(N__30652));
    InMux I__5848 (
            .O(N__30690),
            .I(N__30648));
    Span4Mux_h I__5847 (
            .O(N__30687),
            .I(N__30645));
    LocalMux I__5846 (
            .O(N__30684),
            .I(N__30642));
    LocalMux I__5845 (
            .O(N__30681),
            .I(N__30639));
    LocalMux I__5844 (
            .O(N__30676),
            .I(N__30636));
    LocalMux I__5843 (
            .O(N__30667),
            .I(N__30629));
    LocalMux I__5842 (
            .O(N__30664),
            .I(N__30629));
    LocalMux I__5841 (
            .O(N__30655),
            .I(N__30629));
    Span4Mux_v I__5840 (
            .O(N__30652),
            .I(N__30626));
    InMux I__5839 (
            .O(N__30651),
            .I(N__30623));
    LocalMux I__5838 (
            .O(N__30648),
            .I(N__30618));
    Span4Mux_v I__5837 (
            .O(N__30645),
            .I(N__30618));
    Span4Mux_h I__5836 (
            .O(N__30642),
            .I(N__30615));
    Span4Mux_h I__5835 (
            .O(N__30639),
            .I(N__30612));
    Span4Mux_h I__5834 (
            .O(N__30636),
            .I(N__30607));
    Span4Mux_v I__5833 (
            .O(N__30629),
            .I(N__30607));
    Span4Mux_h I__5832 (
            .O(N__30626),
            .I(N__30604));
    LocalMux I__5831 (
            .O(N__30623),
            .I(N__30601));
    Span4Mux_h I__5830 (
            .O(N__30618),
            .I(N__30598));
    Span4Mux_h I__5829 (
            .O(N__30615),
            .I(N__30593));
    Span4Mux_v I__5828 (
            .O(N__30612),
            .I(N__30593));
    Span4Mux_h I__5827 (
            .O(N__30607),
            .I(N__30590));
    Odrv4 I__5826 (
            .O(N__30604),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_20_c_RNISVKK ));
    Odrv12 I__5825 (
            .O(N__30601),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_20_c_RNISVKK ));
    Odrv4 I__5824 (
            .O(N__30598),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_20_c_RNISVKK ));
    Odrv4 I__5823 (
            .O(N__30593),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_20_c_RNISVKK ));
    Odrv4 I__5822 (
            .O(N__30590),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_20_c_RNISVKK ));
    InMux I__5821 (
            .O(N__30579),
            .I(N__30574));
    IoInMux I__5820 (
            .O(N__30578),
            .I(N__30571));
    InMux I__5819 (
            .O(N__30577),
            .I(N__30568));
    LocalMux I__5818 (
            .O(N__30574),
            .I(N__30563));
    LocalMux I__5817 (
            .O(N__30571),
            .I(N__30560));
    LocalMux I__5816 (
            .O(N__30568),
            .I(N__30557));
    InMux I__5815 (
            .O(N__30567),
            .I(N__30552));
    InMux I__5814 (
            .O(N__30566),
            .I(N__30552));
    Span4Mux_v I__5813 (
            .O(N__30563),
            .I(N__30549));
    Span4Mux_s1_v I__5812 (
            .O(N__30560),
            .I(N__30546));
    Span4Mux_v I__5811 (
            .O(N__30557),
            .I(N__30543));
    LocalMux I__5810 (
            .O(N__30552),
            .I(N__30540));
    Span4Mux_h I__5809 (
            .O(N__30549),
            .I(N__30537));
    Span4Mux_v I__5808 (
            .O(N__30546),
            .I(N__30534));
    Span4Mux_v I__5807 (
            .O(N__30543),
            .I(N__30529));
    Span4Mux_h I__5806 (
            .O(N__30540),
            .I(N__30529));
    Sp12to4 I__5805 (
            .O(N__30537),
            .I(N__30525));
    Span4Mux_h I__5804 (
            .O(N__30534),
            .I(N__30520));
    Span4Mux_v I__5803 (
            .O(N__30529),
            .I(N__30520));
    InMux I__5802 (
            .O(N__30528),
            .I(N__30517));
    Span12Mux_v I__5801 (
            .O(N__30525),
            .I(N__30514));
    Odrv4 I__5800 (
            .O(N__30520),
            .I(debug_CH3_20A_c));
    LocalMux I__5799 (
            .O(N__30517),
            .I(debug_CH3_20A_c));
    Odrv12 I__5798 (
            .O(N__30514),
            .I(debug_CH3_20A_c));
    IoInMux I__5797 (
            .O(N__30507),
            .I(N__30504));
    LocalMux I__5796 (
            .O(N__30504),
            .I(N__30501));
    Odrv4 I__5795 (
            .O(N__30501),
            .I(debug_CH3_20A_c_0));
    InMux I__5794 (
            .O(N__30498),
            .I(N__30495));
    LocalMux I__5793 (
            .O(N__30495),
            .I(N__30491));
    InMux I__5792 (
            .O(N__30494),
            .I(N__30488));
    Span4Mux_h I__5791 (
            .O(N__30491),
            .I(N__30485));
    LocalMux I__5790 (
            .O(N__30488),
            .I(\pid_alt.error_i_acummZ0Z_7 ));
    Odrv4 I__5789 (
            .O(N__30485),
            .I(\pid_alt.error_i_acummZ0Z_7 ));
    InMux I__5788 (
            .O(N__30480),
            .I(N__30476));
    InMux I__5787 (
            .O(N__30479),
            .I(N__30472));
    LocalMux I__5786 (
            .O(N__30476),
            .I(N__30469));
    InMux I__5785 (
            .O(N__30475),
            .I(N__30466));
    LocalMux I__5784 (
            .O(N__30472),
            .I(N__30463));
    Span4Mux_v I__5783 (
            .O(N__30469),
            .I(N__30460));
    LocalMux I__5782 (
            .O(N__30466),
            .I(N__30455));
    Span12Mux_v I__5781 (
            .O(N__30463),
            .I(N__30455));
    Span4Mux_h I__5780 (
            .O(N__30460),
            .I(N__30452));
    Odrv12 I__5779 (
            .O(N__30455),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_6_c_RNI3HMQ ));
    Odrv4 I__5778 (
            .O(N__30452),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_6_c_RNI3HMQ ));
    InMux I__5777 (
            .O(N__30447),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_6 ));
    InMux I__5776 (
            .O(N__30444),
            .I(N__30440));
    InMux I__5775 (
            .O(N__30443),
            .I(N__30437));
    LocalMux I__5774 (
            .O(N__30440),
            .I(\pid_alt.error_i_acummZ0Z_8 ));
    LocalMux I__5773 (
            .O(N__30437),
            .I(\pid_alt.error_i_acummZ0Z_8 ));
    InMux I__5772 (
            .O(N__30432),
            .I(N__30426));
    InMux I__5771 (
            .O(N__30431),
            .I(N__30426));
    LocalMux I__5770 (
            .O(N__30426),
            .I(N__30423));
    Span4Mux_h I__5769 (
            .O(N__30423),
            .I(N__30419));
    InMux I__5768 (
            .O(N__30422),
            .I(N__30416));
    Span4Mux_v I__5767 (
            .O(N__30419),
            .I(N__30413));
    LocalMux I__5766 (
            .O(N__30416),
            .I(N__30410));
    Span4Mux_h I__5765 (
            .O(N__30413),
            .I(N__30407));
    Odrv4 I__5764 (
            .O(N__30410),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_7_c_RNI6LNQ ));
    Odrv4 I__5763 (
            .O(N__30407),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_7_c_RNI6LNQ ));
    InMux I__5762 (
            .O(N__30402),
            .I(bfn_13_22_0_));
    CascadeMux I__5761 (
            .O(N__30399),
            .I(N__30396));
    InMux I__5760 (
            .O(N__30396),
            .I(N__30392));
    CascadeMux I__5759 (
            .O(N__30395),
            .I(N__30389));
    LocalMux I__5758 (
            .O(N__30392),
            .I(N__30386));
    InMux I__5757 (
            .O(N__30389),
            .I(N__30383));
    Odrv4 I__5756 (
            .O(N__30386),
            .I(\pid_alt.error_i_acummZ0Z_9 ));
    LocalMux I__5755 (
            .O(N__30383),
            .I(\pid_alt.error_i_acummZ0Z_9 ));
    InMux I__5754 (
            .O(N__30378),
            .I(N__30371));
    InMux I__5753 (
            .O(N__30377),
            .I(N__30371));
    InMux I__5752 (
            .O(N__30376),
            .I(N__30368));
    LocalMux I__5751 (
            .O(N__30371),
            .I(N__30365));
    LocalMux I__5750 (
            .O(N__30368),
            .I(N__30360));
    Span12Mux_v I__5749 (
            .O(N__30365),
            .I(N__30360));
    Odrv12 I__5748 (
            .O(N__30360),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_8_c_RNI9POQ ));
    InMux I__5747 (
            .O(N__30357),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_8 ));
    CascadeMux I__5746 (
            .O(N__30354),
            .I(N__30351));
    InMux I__5745 (
            .O(N__30351),
            .I(N__30347));
    InMux I__5744 (
            .O(N__30350),
            .I(N__30344));
    LocalMux I__5743 (
            .O(N__30347),
            .I(\pid_alt.error_i_acummZ0Z_10 ));
    LocalMux I__5742 (
            .O(N__30344),
            .I(\pid_alt.error_i_acummZ0Z_10 ));
    InMux I__5741 (
            .O(N__30339),
            .I(N__30335));
    InMux I__5740 (
            .O(N__30338),
            .I(N__30331));
    LocalMux I__5739 (
            .O(N__30335),
            .I(N__30328));
    InMux I__5738 (
            .O(N__30334),
            .I(N__30325));
    LocalMux I__5737 (
            .O(N__30331),
            .I(N__30320));
    Span4Mux_h I__5736 (
            .O(N__30328),
            .I(N__30320));
    LocalMux I__5735 (
            .O(N__30325),
            .I(N__30317));
    Span4Mux_v I__5734 (
            .O(N__30320),
            .I(N__30314));
    Span4Mux_h I__5733 (
            .O(N__30317),
            .I(N__30311));
    Span4Mux_h I__5732 (
            .O(N__30314),
            .I(N__30308));
    Odrv4 I__5731 (
            .O(N__30311),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_9_c_RNIQN3F ));
    Odrv4 I__5730 (
            .O(N__30308),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_9_c_RNIQN3F ));
    InMux I__5729 (
            .O(N__30303),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_9 ));
    InMux I__5728 (
            .O(N__30300),
            .I(N__30293));
    InMux I__5727 (
            .O(N__30299),
            .I(N__30293));
    InMux I__5726 (
            .O(N__30298),
            .I(N__30290));
    LocalMux I__5725 (
            .O(N__30293),
            .I(N__30287));
    LocalMux I__5724 (
            .O(N__30290),
            .I(N__30284));
    Sp12to4 I__5723 (
            .O(N__30287),
            .I(N__30281));
    Span4Mux_h I__5722 (
            .O(N__30284),
            .I(N__30278));
    Span12Mux_v I__5721 (
            .O(N__30281),
            .I(N__30275));
    Odrv4 I__5720 (
            .O(N__30278),
            .I(\pid_alt.error_i_reg_esr_RNI4NMPZ0Z_11 ));
    Odrv12 I__5719 (
            .O(N__30275),
            .I(\pid_alt.error_i_reg_esr_RNI4NMPZ0Z_11 ));
    InMux I__5718 (
            .O(N__30270),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_10 ));
    InMux I__5717 (
            .O(N__30267),
            .I(N__30263));
    InMux I__5716 (
            .O(N__30266),
            .I(N__30260));
    LocalMux I__5715 (
            .O(N__30263),
            .I(\pid_alt.error_i_acummZ0Z_12 ));
    LocalMux I__5714 (
            .O(N__30260),
            .I(\pid_alt.error_i_acummZ0Z_12 ));
    InMux I__5713 (
            .O(N__30255),
            .I(N__30251));
    InMux I__5712 (
            .O(N__30254),
            .I(N__30247));
    LocalMux I__5711 (
            .O(N__30251),
            .I(N__30244));
    InMux I__5710 (
            .O(N__30250),
            .I(N__30241));
    LocalMux I__5709 (
            .O(N__30247),
            .I(N__30238));
    Sp12to4 I__5708 (
            .O(N__30244),
            .I(N__30233));
    LocalMux I__5707 (
            .O(N__30241),
            .I(N__30233));
    Span4Mux_h I__5706 (
            .O(N__30238),
            .I(N__30230));
    Span12Mux_v I__5705 (
            .O(N__30233),
            .I(N__30227));
    Odrv4 I__5704 (
            .O(N__30230),
            .I(\pid_alt.error_i_reg_esr_RNI7RNPZ0Z_12 ));
    Odrv12 I__5703 (
            .O(N__30227),
            .I(\pid_alt.error_i_reg_esr_RNI7RNPZ0Z_12 ));
    InMux I__5702 (
            .O(N__30222),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_11 ));
    InMux I__5701 (
            .O(N__30219),
            .I(N__30216));
    LocalMux I__5700 (
            .O(N__30216),
            .I(N__30211));
    InMux I__5699 (
            .O(N__30215),
            .I(N__30206));
    InMux I__5698 (
            .O(N__30214),
            .I(N__30206));
    Span4Mux_h I__5697 (
            .O(N__30211),
            .I(N__30203));
    LocalMux I__5696 (
            .O(N__30206),
            .I(N__30200));
    Span4Mux_h I__5695 (
            .O(N__30203),
            .I(N__30197));
    Span12Mux_v I__5694 (
            .O(N__30200),
            .I(N__30194));
    Odrv4 I__5693 (
            .O(N__30197),
            .I(\pid_alt.error_i_acumm_esr_RNIJ6LMZ0Z_13 ));
    Odrv12 I__5692 (
            .O(N__30194),
            .I(\pid_alt.error_i_acumm_esr_RNIJ6LMZ0Z_13 ));
    InMux I__5691 (
            .O(N__30189),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_12 ));
    InMux I__5690 (
            .O(N__30186),
            .I(N__30180));
    InMux I__5689 (
            .O(N__30185),
            .I(N__30180));
    LocalMux I__5688 (
            .O(N__30180),
            .I(N__30176));
    InMux I__5687 (
            .O(N__30179),
            .I(N__30173));
    Span4Mux_h I__5686 (
            .O(N__30176),
            .I(N__30170));
    LocalMux I__5685 (
            .O(N__30173),
            .I(N__30167));
    Span4Mux_v I__5684 (
            .O(N__30170),
            .I(N__30164));
    Span4Mux_v I__5683 (
            .O(N__30167),
            .I(N__30159));
    Span4Mux_h I__5682 (
            .O(N__30164),
            .I(N__30159));
    Odrv4 I__5681 (
            .O(N__30159),
            .I(\pid_alt.error_i_reg_esr_RNI15KJZ0Z_14 ));
    InMux I__5680 (
            .O(N__30156),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_13 ));
    InMux I__5679 (
            .O(N__30153),
            .I(N__30150));
    LocalMux I__5678 (
            .O(N__30150),
            .I(N__30147));
    Span4Mux_v I__5677 (
            .O(N__30147),
            .I(N__30144));
    Odrv4 I__5676 (
            .O(N__30144),
            .I(scaler_3_data_14));
    InMux I__5675 (
            .O(N__30141),
            .I(bfn_13_20_0_));
    InMux I__5674 (
            .O(N__30138),
            .I(N__30134));
    CascadeMux I__5673 (
            .O(N__30137),
            .I(N__30131));
    LocalMux I__5672 (
            .O(N__30134),
            .I(N__30128));
    InMux I__5671 (
            .O(N__30131),
            .I(N__30125));
    Span4Mux_v I__5670 (
            .O(N__30128),
            .I(N__30120));
    LocalMux I__5669 (
            .O(N__30125),
            .I(N__30120));
    Span4Mux_h I__5668 (
            .O(N__30120),
            .I(N__30117));
    Span4Mux_v I__5667 (
            .O(N__30117),
            .I(N__30114));
    Span4Mux_h I__5666 (
            .O(N__30114),
            .I(N__30111));
    Odrv4 I__5665 (
            .O(N__30111),
            .I(\pid_alt.un1_pid_prereg_0 ));
    InMux I__5664 (
            .O(N__30108),
            .I(N__30105));
    LocalMux I__5663 (
            .O(N__30105),
            .I(\pid_alt.error_i_acummZ0Z_1 ));
    CascadeMux I__5662 (
            .O(N__30102),
            .I(N__30098));
    CascadeMux I__5661 (
            .O(N__30101),
            .I(N__30095));
    InMux I__5660 (
            .O(N__30098),
            .I(N__30092));
    InMux I__5659 (
            .O(N__30095),
            .I(N__30089));
    LocalMux I__5658 (
            .O(N__30092),
            .I(N__30086));
    LocalMux I__5657 (
            .O(N__30089),
            .I(N__30082));
    Span4Mux_v I__5656 (
            .O(N__30086),
            .I(N__30079));
    InMux I__5655 (
            .O(N__30085),
            .I(N__30076));
    Span4Mux_h I__5654 (
            .O(N__30082),
            .I(N__30073));
    Sp12to4 I__5653 (
            .O(N__30079),
            .I(N__30070));
    LocalMux I__5652 (
            .O(N__30076),
            .I(N__30067));
    Span4Mux_v I__5651 (
            .O(N__30073),
            .I(N__30064));
    Span12Mux_v I__5650 (
            .O(N__30070),
            .I(N__30061));
    Span4Mux_h I__5649 (
            .O(N__30067),
            .I(N__30058));
    Span4Mux_h I__5648 (
            .O(N__30064),
            .I(N__30055));
    Odrv12 I__5647 (
            .O(N__30061),
            .I(\pid_alt.error_i_acumm_esr_RNIQMD91Z0Z_1 ));
    Odrv4 I__5646 (
            .O(N__30058),
            .I(\pid_alt.error_i_acumm_esr_RNIQMD91Z0Z_1 ));
    Odrv4 I__5645 (
            .O(N__30055),
            .I(\pid_alt.error_i_acumm_esr_RNIQMD91Z0Z_1 ));
    InMux I__5644 (
            .O(N__30048),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_0 ));
    InMux I__5643 (
            .O(N__30045),
            .I(N__30042));
    LocalMux I__5642 (
            .O(N__30042),
            .I(\pid_alt.error_i_acummZ0Z_2 ));
    InMux I__5641 (
            .O(N__30039),
            .I(N__30036));
    LocalMux I__5640 (
            .O(N__30036),
            .I(N__30032));
    CascadeMux I__5639 (
            .O(N__30035),
            .I(N__30029));
    Span4Mux_h I__5638 (
            .O(N__30032),
            .I(N__30025));
    InMux I__5637 (
            .O(N__30029),
            .I(N__30022));
    InMux I__5636 (
            .O(N__30028),
            .I(N__30019));
    Sp12to4 I__5635 (
            .O(N__30025),
            .I(N__30014));
    LocalMux I__5634 (
            .O(N__30022),
            .I(N__30014));
    LocalMux I__5633 (
            .O(N__30019),
            .I(N__30009));
    Span12Mux_v I__5632 (
            .O(N__30014),
            .I(N__30009));
    Odrv12 I__5631 (
            .O(N__30009),
            .I(\pid_alt.error_i_acumm_esr_RNITQE91Z0Z_2 ));
    InMux I__5630 (
            .O(N__30006),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_1 ));
    InMux I__5629 (
            .O(N__30003),
            .I(N__30000));
    LocalMux I__5628 (
            .O(N__30000),
            .I(\pid_alt.error_i_acummZ0Z_3 ));
    InMux I__5627 (
            .O(N__29997),
            .I(N__29993));
    CascadeMux I__5626 (
            .O(N__29996),
            .I(N__29990));
    LocalMux I__5625 (
            .O(N__29993),
            .I(N__29986));
    InMux I__5624 (
            .O(N__29990),
            .I(N__29983));
    InMux I__5623 (
            .O(N__29989),
            .I(N__29980));
    Span4Mux_h I__5622 (
            .O(N__29986),
            .I(N__29975));
    LocalMux I__5621 (
            .O(N__29983),
            .I(N__29975));
    LocalMux I__5620 (
            .O(N__29980),
            .I(N__29972));
    Span4Mux_h I__5619 (
            .O(N__29975),
            .I(N__29969));
    Span4Mux_v I__5618 (
            .O(N__29972),
            .I(N__29964));
    Span4Mux_v I__5617 (
            .O(N__29969),
            .I(N__29964));
    Span4Mux_h I__5616 (
            .O(N__29964),
            .I(N__29961));
    Odrv4 I__5615 (
            .O(N__29961),
            .I(\pid_alt.error_i_acumm_esr_RNI0VF91Z0Z_3 ));
    InMux I__5614 (
            .O(N__29958),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_2 ));
    InMux I__5613 (
            .O(N__29955),
            .I(N__29952));
    LocalMux I__5612 (
            .O(N__29952),
            .I(\pid_alt.error_i_acummZ0Z_4 ));
    InMux I__5611 (
            .O(N__29949),
            .I(N__29940));
    InMux I__5610 (
            .O(N__29948),
            .I(N__29940));
    InMux I__5609 (
            .O(N__29947),
            .I(N__29940));
    LocalMux I__5608 (
            .O(N__29940),
            .I(N__29937));
    Span4Mux_h I__5607 (
            .O(N__29937),
            .I(N__29934));
    Span4Mux_v I__5606 (
            .O(N__29934),
            .I(N__29931));
    Odrv4 I__5605 (
            .O(N__29931),
            .I(\pid_alt.error_i_acumm_esr_RNI33H91Z0Z_4 ));
    InMux I__5604 (
            .O(N__29928),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_3 ));
    CascadeMux I__5603 (
            .O(N__29925),
            .I(N__29921));
    InMux I__5602 (
            .O(N__29924),
            .I(N__29918));
    InMux I__5601 (
            .O(N__29921),
            .I(N__29915));
    LocalMux I__5600 (
            .O(N__29918),
            .I(\pid_alt.error_i_acummZ0Z_5 ));
    LocalMux I__5599 (
            .O(N__29915),
            .I(\pid_alt.error_i_acummZ0Z_5 ));
    InMux I__5598 (
            .O(N__29910),
            .I(N__29907));
    LocalMux I__5597 (
            .O(N__29907),
            .I(N__29902));
    InMux I__5596 (
            .O(N__29906),
            .I(N__29897));
    InMux I__5595 (
            .O(N__29905),
            .I(N__29897));
    Span4Mux_h I__5594 (
            .O(N__29902),
            .I(N__29894));
    LocalMux I__5593 (
            .O(N__29897),
            .I(N__29891));
    Sp12to4 I__5592 (
            .O(N__29894),
            .I(N__29886));
    Span12Mux_h I__5591 (
            .O(N__29891),
            .I(N__29886));
    Odrv12 I__5590 (
            .O(N__29886),
            .I(\pid_alt.error_i_reg_esr_RNIT8KA1Z0Z_5 ));
    InMux I__5589 (
            .O(N__29883),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_4 ));
    InMux I__5588 (
            .O(N__29880),
            .I(N__29874));
    InMux I__5587 (
            .O(N__29879),
            .I(N__29874));
    LocalMux I__5586 (
            .O(N__29874),
            .I(N__29871));
    Span4Mux_h I__5585 (
            .O(N__29871),
            .I(N__29867));
    InMux I__5584 (
            .O(N__29870),
            .I(N__29864));
    Span4Mux_v I__5583 (
            .O(N__29867),
            .I(N__29861));
    LocalMux I__5582 (
            .O(N__29864),
            .I(N__29858));
    Span4Mux_h I__5581 (
            .O(N__29861),
            .I(N__29855));
    Odrv4 I__5580 (
            .O(N__29858),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_5_c_RNI0DLQ ));
    Odrv4 I__5579 (
            .O(N__29855),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_5_c_RNI0DLQ ));
    InMux I__5578 (
            .O(N__29850),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_5 ));
    InMux I__5577 (
            .O(N__29847),
            .I(N__29844));
    LocalMux I__5576 (
            .O(N__29844),
            .I(scaler_4_data_14));
    InMux I__5575 (
            .O(N__29841),
            .I(bfn_13_18_0_));
    InMux I__5574 (
            .O(N__29838),
            .I(\ppm_encoder_1.un1_elevator_cry_6 ));
    InMux I__5573 (
            .O(N__29835),
            .I(N__29831));
    InMux I__5572 (
            .O(N__29834),
            .I(N__29828));
    LocalMux I__5571 (
            .O(N__29831),
            .I(N__29825));
    LocalMux I__5570 (
            .O(N__29828),
            .I(N__29820));
    Span4Mux_v I__5569 (
            .O(N__29825),
            .I(N__29820));
    Odrv4 I__5568 (
            .O(N__29820),
            .I(scaler_3_data_8));
    InMux I__5567 (
            .O(N__29817),
            .I(N__29814));
    LocalMux I__5566 (
            .O(N__29814),
            .I(N__29811));
    Odrv12 I__5565 (
            .O(N__29811),
            .I(\ppm_encoder_1.un1_elevator_cry_7_THRU_CO ));
    InMux I__5564 (
            .O(N__29808),
            .I(\ppm_encoder_1.un1_elevator_cry_7 ));
    InMux I__5563 (
            .O(N__29805),
            .I(\ppm_encoder_1.un1_elevator_cry_8 ));
    InMux I__5562 (
            .O(N__29802),
            .I(\ppm_encoder_1.un1_elevator_cry_9 ));
    InMux I__5561 (
            .O(N__29799),
            .I(\ppm_encoder_1.un1_elevator_cry_10 ));
    InMux I__5560 (
            .O(N__29796),
            .I(\ppm_encoder_1.un1_elevator_cry_11 ));
    InMux I__5559 (
            .O(N__29793),
            .I(\ppm_encoder_1.un1_elevator_cry_12 ));
    InMux I__5558 (
            .O(N__29790),
            .I(N__29786));
    InMux I__5557 (
            .O(N__29789),
            .I(N__29783));
    LocalMux I__5556 (
            .O(N__29786),
            .I(scaler_4_data_6));
    LocalMux I__5555 (
            .O(N__29783),
            .I(scaler_4_data_6));
    InMux I__5554 (
            .O(N__29778),
            .I(N__29774));
    InMux I__5553 (
            .O(N__29777),
            .I(N__29771));
    LocalMux I__5552 (
            .O(N__29774),
            .I(scaler_4_data_7));
    LocalMux I__5551 (
            .O(N__29771),
            .I(scaler_4_data_7));
    InMux I__5550 (
            .O(N__29766),
            .I(N__29763));
    LocalMux I__5549 (
            .O(N__29763),
            .I(\ppm_encoder_1.un1_rudder_cry_6_THRU_CO ));
    InMux I__5548 (
            .O(N__29760),
            .I(\ppm_encoder_1.un1_rudder_cry_6 ));
    InMux I__5547 (
            .O(N__29757),
            .I(\ppm_encoder_1.un1_rudder_cry_7 ));
    InMux I__5546 (
            .O(N__29754),
            .I(N__29750));
    InMux I__5545 (
            .O(N__29753),
            .I(N__29747));
    LocalMux I__5544 (
            .O(N__29750),
            .I(scaler_4_data_9));
    LocalMux I__5543 (
            .O(N__29747),
            .I(scaler_4_data_9));
    InMux I__5542 (
            .O(N__29742),
            .I(N__29739));
    LocalMux I__5541 (
            .O(N__29739),
            .I(\ppm_encoder_1.un1_rudder_cry_8_THRU_CO ));
    InMux I__5540 (
            .O(N__29736),
            .I(\ppm_encoder_1.un1_rudder_cry_8 ));
    InMux I__5539 (
            .O(N__29733),
            .I(\ppm_encoder_1.un1_rudder_cry_9 ));
    InMux I__5538 (
            .O(N__29730),
            .I(\ppm_encoder_1.un1_rudder_cry_10 ));
    InMux I__5537 (
            .O(N__29727),
            .I(\ppm_encoder_1.un1_rudder_cry_11 ));
    InMux I__5536 (
            .O(N__29724),
            .I(\ppm_encoder_1.un1_rudder_cry_12 ));
    InMux I__5535 (
            .O(N__29721),
            .I(N__29718));
    LocalMux I__5534 (
            .O(N__29718),
            .I(N__29715));
    Span4Mux_v I__5533 (
            .O(N__29715),
            .I(N__29709));
    CascadeMux I__5532 (
            .O(N__29714),
            .I(N__29706));
    InMux I__5531 (
            .O(N__29713),
            .I(N__29701));
    InMux I__5530 (
            .O(N__29712),
            .I(N__29698));
    Span4Mux_h I__5529 (
            .O(N__29709),
            .I(N__29695));
    InMux I__5528 (
            .O(N__29706),
            .I(N__29688));
    InMux I__5527 (
            .O(N__29705),
            .I(N__29688));
    InMux I__5526 (
            .O(N__29704),
            .I(N__29688));
    LocalMux I__5525 (
            .O(N__29701),
            .I(N__29683));
    LocalMux I__5524 (
            .O(N__29698),
            .I(N__29683));
    Odrv4 I__5523 (
            .O(N__29695),
            .I(\dron_frame_decoder_1.stateZ0Z_6 ));
    LocalMux I__5522 (
            .O(N__29688),
            .I(\dron_frame_decoder_1.stateZ0Z_6 ));
    Odrv4 I__5521 (
            .O(N__29683),
            .I(\dron_frame_decoder_1.stateZ0Z_6 ));
    InMux I__5520 (
            .O(N__29676),
            .I(N__29673));
    LocalMux I__5519 (
            .O(N__29673),
            .I(N__29669));
    InMux I__5518 (
            .O(N__29672),
            .I(N__29664));
    Span4Mux_v I__5517 (
            .O(N__29669),
            .I(N__29658));
    InMux I__5516 (
            .O(N__29668),
            .I(N__29654));
    InMux I__5515 (
            .O(N__29667),
            .I(N__29651));
    LocalMux I__5514 (
            .O(N__29664),
            .I(N__29648));
    CascadeMux I__5513 (
            .O(N__29663),
            .I(N__29644));
    InMux I__5512 (
            .O(N__29662),
            .I(N__29637));
    InMux I__5511 (
            .O(N__29661),
            .I(N__29637));
    Span4Mux_h I__5510 (
            .O(N__29658),
            .I(N__29634));
    InMux I__5509 (
            .O(N__29657),
            .I(N__29631));
    LocalMux I__5508 (
            .O(N__29654),
            .I(N__29628));
    LocalMux I__5507 (
            .O(N__29651),
            .I(N__29623));
    Span4Mux_h I__5506 (
            .O(N__29648),
            .I(N__29623));
    InMux I__5505 (
            .O(N__29647),
            .I(N__29614));
    InMux I__5504 (
            .O(N__29644),
            .I(N__29614));
    InMux I__5503 (
            .O(N__29643),
            .I(N__29614));
    InMux I__5502 (
            .O(N__29642),
            .I(N__29614));
    LocalMux I__5501 (
            .O(N__29637),
            .I(uart_drone_data_rdy));
    Odrv4 I__5500 (
            .O(N__29634),
            .I(uart_drone_data_rdy));
    LocalMux I__5499 (
            .O(N__29631),
            .I(uart_drone_data_rdy));
    Odrv4 I__5498 (
            .O(N__29628),
            .I(uart_drone_data_rdy));
    Odrv4 I__5497 (
            .O(N__29623),
            .I(uart_drone_data_rdy));
    LocalMux I__5496 (
            .O(N__29614),
            .I(uart_drone_data_rdy));
    InMux I__5495 (
            .O(N__29601),
            .I(N__29597));
    IoInMux I__5494 (
            .O(N__29600),
            .I(N__29594));
    LocalMux I__5493 (
            .O(N__29597),
            .I(N__29591));
    LocalMux I__5492 (
            .O(N__29594),
            .I(N__29587));
    Span4Mux_v I__5491 (
            .O(N__29591),
            .I(N__29584));
    InMux I__5490 (
            .O(N__29590),
            .I(N__29581));
    Span12Mux_s2_v I__5489 (
            .O(N__29587),
            .I(N__29578));
    Span4Mux_h I__5488 (
            .O(N__29584),
            .I(N__29572));
    LocalMux I__5487 (
            .O(N__29581),
            .I(N__29572));
    Span12Mux_v I__5486 (
            .O(N__29578),
            .I(N__29569));
    InMux I__5485 (
            .O(N__29577),
            .I(N__29566));
    Span4Mux_h I__5484 (
            .O(N__29572),
            .I(N__29563));
    Odrv12 I__5483 (
            .O(N__29569),
            .I(debug_CH1_0A_c));
    LocalMux I__5482 (
            .O(N__29566),
            .I(debug_CH1_0A_c));
    Odrv4 I__5481 (
            .O(N__29563),
            .I(debug_CH1_0A_c));
    InMux I__5480 (
            .O(N__29556),
            .I(N__29553));
    LocalMux I__5479 (
            .O(N__29553),
            .I(N__29547));
    InMux I__5478 (
            .O(N__29552),
            .I(N__29544));
    InMux I__5477 (
            .O(N__29551),
            .I(N__29541));
    CascadeMux I__5476 (
            .O(N__29550),
            .I(N__29538));
    Span4Mux_h I__5475 (
            .O(N__29547),
            .I(N__29535));
    LocalMux I__5474 (
            .O(N__29544),
            .I(N__29532));
    LocalMux I__5473 (
            .O(N__29541),
            .I(N__29529));
    InMux I__5472 (
            .O(N__29538),
            .I(N__29526));
    Odrv4 I__5471 (
            .O(N__29535),
            .I(frame_decoder_OFF4data_0));
    Odrv4 I__5470 (
            .O(N__29532),
            .I(frame_decoder_OFF4data_0));
    Odrv4 I__5469 (
            .O(N__29529),
            .I(frame_decoder_OFF4data_0));
    LocalMux I__5468 (
            .O(N__29526),
            .I(frame_decoder_OFF4data_0));
    InMux I__5467 (
            .O(N__29517),
            .I(N__29514));
    LocalMux I__5466 (
            .O(N__29514),
            .I(N__29509));
    InMux I__5465 (
            .O(N__29513),
            .I(N__29506));
    InMux I__5464 (
            .O(N__29512),
            .I(N__29503));
    Span4Mux_h I__5463 (
            .O(N__29509),
            .I(N__29500));
    LocalMux I__5462 (
            .O(N__29506),
            .I(N__29497));
    LocalMux I__5461 (
            .O(N__29503),
            .I(N__29494));
    Span4Mux_v I__5460 (
            .O(N__29500),
            .I(N__29488));
    Span4Mux_h I__5459 (
            .O(N__29497),
            .I(N__29488));
    Span4Mux_v I__5458 (
            .O(N__29494),
            .I(N__29485));
    InMux I__5457 (
            .O(N__29493),
            .I(N__29482));
    Odrv4 I__5456 (
            .O(N__29488),
            .I(frame_decoder_CH4data_0));
    Odrv4 I__5455 (
            .O(N__29485),
            .I(frame_decoder_CH4data_0));
    LocalMux I__5454 (
            .O(N__29482),
            .I(frame_decoder_CH4data_0));
    InMux I__5453 (
            .O(N__29475),
            .I(N__29471));
    CascadeMux I__5452 (
            .O(N__29474),
            .I(N__29468));
    LocalMux I__5451 (
            .O(N__29471),
            .I(N__29465));
    InMux I__5450 (
            .O(N__29468),
            .I(N__29462));
    Odrv12 I__5449 (
            .O(N__29465),
            .I(scaler_4_data_4));
    LocalMux I__5448 (
            .O(N__29462),
            .I(scaler_4_data_4));
    IoInMux I__5447 (
            .O(N__29457),
            .I(N__29454));
    LocalMux I__5446 (
            .O(N__29454),
            .I(N__29450));
    CascadeMux I__5445 (
            .O(N__29453),
            .I(N__29447));
    Span12Mux_s3_v I__5444 (
            .O(N__29450),
            .I(N__29444));
    InMux I__5443 (
            .O(N__29447),
            .I(N__29441));
    Odrv12 I__5442 (
            .O(N__29444),
            .I(ppm_output_c));
    LocalMux I__5441 (
            .O(N__29441),
            .I(ppm_output_c));
    InMux I__5440 (
            .O(N__29436),
            .I(N__29432));
    InMux I__5439 (
            .O(N__29435),
            .I(N__29429));
    LocalMux I__5438 (
            .O(N__29432),
            .I(N__29424));
    LocalMux I__5437 (
            .O(N__29429),
            .I(N__29424));
    Span4Mux_v I__5436 (
            .O(N__29424),
            .I(N__29421));
    Odrv4 I__5435 (
            .O(N__29421),
            .I(throttle_command_10));
    InMux I__5434 (
            .O(N__29418),
            .I(N__29415));
    LocalMux I__5433 (
            .O(N__29415),
            .I(N__29412));
    Odrv4 I__5432 (
            .O(N__29412),
            .I(\ppm_encoder_1.un1_throttle_cry_9_THRU_CO ));
    InMux I__5431 (
            .O(N__29409),
            .I(N__29406));
    LocalMux I__5430 (
            .O(N__29406),
            .I(N__29403));
    Odrv12 I__5429 (
            .O(N__29403),
            .I(\ppm_encoder_1.un1_throttle_cry_3_THRU_CO ));
    InMux I__5428 (
            .O(N__29400),
            .I(N__29397));
    LocalMux I__5427 (
            .O(N__29397),
            .I(N__29393));
    CascadeMux I__5426 (
            .O(N__29396),
            .I(N__29389));
    Span4Mux_h I__5425 (
            .O(N__29393),
            .I(N__29386));
    InMux I__5424 (
            .O(N__29392),
            .I(N__29383));
    InMux I__5423 (
            .O(N__29389),
            .I(N__29380));
    Span4Mux_h I__5422 (
            .O(N__29386),
            .I(N__29377));
    LocalMux I__5421 (
            .O(N__29383),
            .I(N__29374));
    LocalMux I__5420 (
            .O(N__29380),
            .I(throttle_command_4));
    Odrv4 I__5419 (
            .O(N__29377),
            .I(throttle_command_4));
    Odrv12 I__5418 (
            .O(N__29374),
            .I(throttle_command_4));
    InMux I__5417 (
            .O(N__29367),
            .I(\ppm_encoder_1.un1_throttle_cry_8 ));
    InMux I__5416 (
            .O(N__29364),
            .I(\ppm_encoder_1.un1_throttle_cry_9 ));
    InMux I__5415 (
            .O(N__29361),
            .I(\ppm_encoder_1.un1_throttle_cry_10 ));
    InMux I__5414 (
            .O(N__29358),
            .I(\ppm_encoder_1.un1_throttle_cry_11 ));
    InMux I__5413 (
            .O(N__29355),
            .I(\ppm_encoder_1.un1_throttle_cry_12 ));
    InMux I__5412 (
            .O(N__29352),
            .I(\ppm_encoder_1.un1_throttle_cry_13 ));
    InMux I__5411 (
            .O(N__29349),
            .I(N__29346));
    LocalMux I__5410 (
            .O(N__29346),
            .I(N__29342));
    CascadeMux I__5409 (
            .O(N__29345),
            .I(N__29338));
    Span4Mux_v I__5408 (
            .O(N__29342),
            .I(N__29335));
    InMux I__5407 (
            .O(N__29341),
            .I(N__29332));
    InMux I__5406 (
            .O(N__29338),
            .I(N__29329));
    Span4Mux_h I__5405 (
            .O(N__29335),
            .I(N__29324));
    LocalMux I__5404 (
            .O(N__29332),
            .I(N__29324));
    LocalMux I__5403 (
            .O(N__29329),
            .I(throttle_command_2));
    Odrv4 I__5402 (
            .O(N__29324),
            .I(throttle_command_2));
    InMux I__5401 (
            .O(N__29319),
            .I(N__29316));
    LocalMux I__5400 (
            .O(N__29316),
            .I(N__29313));
    Odrv4 I__5399 (
            .O(N__29313),
            .I(\ppm_encoder_1.un1_throttle_cry_1_THRU_CO ));
    InMux I__5398 (
            .O(N__29310),
            .I(N__29307));
    LocalMux I__5397 (
            .O(N__29307),
            .I(N__29304));
    Odrv4 I__5396 (
            .O(N__29304),
            .I(\ppm_encoder_1.un1_throttle_cry_0_THRU_CO ));
    InMux I__5395 (
            .O(N__29301),
            .I(N__29297));
    CascadeMux I__5394 (
            .O(N__29300),
            .I(N__29293));
    LocalMux I__5393 (
            .O(N__29297),
            .I(N__29290));
    InMux I__5392 (
            .O(N__29296),
            .I(N__29287));
    InMux I__5391 (
            .O(N__29293),
            .I(N__29284));
    Span4Mux_h I__5390 (
            .O(N__29290),
            .I(N__29281));
    LocalMux I__5389 (
            .O(N__29287),
            .I(N__29278));
    LocalMux I__5388 (
            .O(N__29284),
            .I(throttle_command_1));
    Odrv4 I__5387 (
            .O(N__29281),
            .I(throttle_command_1));
    Odrv4 I__5386 (
            .O(N__29278),
            .I(throttle_command_1));
    InMux I__5385 (
            .O(N__29271),
            .I(\ppm_encoder_1.un1_throttle_cry_0 ));
    InMux I__5384 (
            .O(N__29268),
            .I(\ppm_encoder_1.un1_throttle_cry_1 ));
    InMux I__5383 (
            .O(N__29265),
            .I(\ppm_encoder_1.un1_throttle_cry_2 ));
    InMux I__5382 (
            .O(N__29262),
            .I(\ppm_encoder_1.un1_throttle_cry_3 ));
    InMux I__5381 (
            .O(N__29259),
            .I(N__29255));
    InMux I__5380 (
            .O(N__29258),
            .I(N__29252));
    LocalMux I__5379 (
            .O(N__29255),
            .I(N__29249));
    LocalMux I__5378 (
            .O(N__29252),
            .I(N__29246));
    Span4Mux_h I__5377 (
            .O(N__29249),
            .I(N__29243));
    Span4Mux_h I__5376 (
            .O(N__29246),
            .I(N__29240));
    Odrv4 I__5375 (
            .O(N__29243),
            .I(throttle_command_5));
    Odrv4 I__5374 (
            .O(N__29240),
            .I(throttle_command_5));
    InMux I__5373 (
            .O(N__29235),
            .I(N__29232));
    LocalMux I__5372 (
            .O(N__29232),
            .I(N__29229));
    Odrv4 I__5371 (
            .O(N__29229),
            .I(\ppm_encoder_1.un1_throttle_cry_4_THRU_CO ));
    InMux I__5370 (
            .O(N__29226),
            .I(\ppm_encoder_1.un1_throttle_cry_4 ));
    InMux I__5369 (
            .O(N__29223),
            .I(\ppm_encoder_1.un1_throttle_cry_5 ));
    InMux I__5368 (
            .O(N__29220),
            .I(\ppm_encoder_1.un1_throttle_cry_6 ));
    InMux I__5367 (
            .O(N__29217),
            .I(bfn_13_14_0_));
    InMux I__5366 (
            .O(N__29214),
            .I(N__29211));
    LocalMux I__5365 (
            .O(N__29211),
            .I(N__29208));
    Odrv12 I__5364 (
            .O(N__29208),
            .I(\uart_pc.data_Auxce_0_0_0 ));
    CascadeMux I__5363 (
            .O(N__29205),
            .I(N__29202));
    InMux I__5362 (
            .O(N__29202),
            .I(N__29199));
    LocalMux I__5361 (
            .O(N__29199),
            .I(N__29196));
    Odrv4 I__5360 (
            .O(N__29196),
            .I(\uart_pc.data_Auxce_0_1 ));
    InMux I__5359 (
            .O(N__29193),
            .I(N__29190));
    LocalMux I__5358 (
            .O(N__29190),
            .I(N__29187));
    Span4Mux_h I__5357 (
            .O(N__29187),
            .I(N__29184));
    Odrv4 I__5356 (
            .O(N__29184),
            .I(\uart_pc.data_Auxce_0_0_4 ));
    InMux I__5355 (
            .O(N__29181),
            .I(N__29177));
    CascadeMux I__5354 (
            .O(N__29180),
            .I(N__29174));
    LocalMux I__5353 (
            .O(N__29177),
            .I(N__29171));
    InMux I__5352 (
            .O(N__29174),
            .I(N__29168));
    Odrv4 I__5351 (
            .O(N__29171),
            .I(scaler_2_data_4));
    LocalMux I__5350 (
            .O(N__29168),
            .I(scaler_2_data_4));
    InMux I__5349 (
            .O(N__29163),
            .I(N__29160));
    LocalMux I__5348 (
            .O(N__29160),
            .I(scaler_2_data_5));
    InMux I__5347 (
            .O(N__29157),
            .I(N__29153));
    CascadeMux I__5346 (
            .O(N__29156),
            .I(N__29150));
    LocalMux I__5345 (
            .O(N__29153),
            .I(N__29147));
    InMux I__5344 (
            .O(N__29150),
            .I(N__29144));
    Odrv4 I__5343 (
            .O(N__29147),
            .I(scaler_3_data_4));
    LocalMux I__5342 (
            .O(N__29144),
            .I(scaler_3_data_4));
    InMux I__5341 (
            .O(N__29139),
            .I(N__29136));
    LocalMux I__5340 (
            .O(N__29136),
            .I(scaler_3_data_5));
    InMux I__5339 (
            .O(N__29133),
            .I(N__29130));
    LocalMux I__5338 (
            .O(N__29130),
            .I(scaler_4_data_5));
    CascadeMux I__5337 (
            .O(N__29127),
            .I(N__29124));
    InMux I__5336 (
            .O(N__29124),
            .I(N__29120));
    InMux I__5335 (
            .O(N__29123),
            .I(N__29117));
    LocalMux I__5334 (
            .O(N__29120),
            .I(N__29114));
    LocalMux I__5333 (
            .O(N__29117),
            .I(\uart_pc.data_AuxZ0Z_7 ));
    Odrv4 I__5332 (
            .O(N__29114),
            .I(\uart_pc.data_AuxZ0Z_7 ));
    SRMux I__5331 (
            .O(N__29109),
            .I(N__29106));
    LocalMux I__5330 (
            .O(N__29106),
            .I(N__29103));
    Odrv12 I__5329 (
            .O(N__29103),
            .I(\uart_pc.state_RNIEAGSZ0Z_4 ));
    InMux I__5328 (
            .O(N__29100),
            .I(N__29097));
    LocalMux I__5327 (
            .O(N__29097),
            .I(\uart_pc.data_Auxce_0_3 ));
    InMux I__5326 (
            .O(N__29094),
            .I(N__29091));
    LocalMux I__5325 (
            .O(N__29091),
            .I(\uart_pc.data_Auxce_0_0_2 ));
    InMux I__5324 (
            .O(N__29088),
            .I(N__29085));
    LocalMux I__5323 (
            .O(N__29085),
            .I(\uart_pc.data_Auxce_0_5 ));
    InMux I__5322 (
            .O(N__29082),
            .I(N__29076));
    CascadeMux I__5321 (
            .O(N__29081),
            .I(N__29073));
    InMux I__5320 (
            .O(N__29080),
            .I(N__29070));
    InMux I__5319 (
            .O(N__29079),
            .I(N__29067));
    LocalMux I__5318 (
            .O(N__29076),
            .I(N__29064));
    InMux I__5317 (
            .O(N__29073),
            .I(N__29061));
    LocalMux I__5316 (
            .O(N__29070),
            .I(frame_decoder_OFF2data_0));
    LocalMux I__5315 (
            .O(N__29067),
            .I(frame_decoder_OFF2data_0));
    Odrv12 I__5314 (
            .O(N__29064),
            .I(frame_decoder_OFF2data_0));
    LocalMux I__5313 (
            .O(N__29061),
            .I(frame_decoder_OFF2data_0));
    InMux I__5312 (
            .O(N__29052),
            .I(N__29048));
    InMux I__5311 (
            .O(N__29051),
            .I(N__29045));
    LocalMux I__5310 (
            .O(N__29048),
            .I(N__29039));
    LocalMux I__5309 (
            .O(N__29045),
            .I(N__29039));
    InMux I__5308 (
            .O(N__29044),
            .I(N__29036));
    Span4Mux_v I__5307 (
            .O(N__29039),
            .I(N__29032));
    LocalMux I__5306 (
            .O(N__29036),
            .I(N__29029));
    InMux I__5305 (
            .O(N__29035),
            .I(N__29026));
    Odrv4 I__5304 (
            .O(N__29032),
            .I(frame_decoder_CH2data_0));
    Odrv4 I__5303 (
            .O(N__29029),
            .I(frame_decoder_CH2data_0));
    LocalMux I__5302 (
            .O(N__29026),
            .I(frame_decoder_CH2data_0));
    InMux I__5301 (
            .O(N__29019),
            .I(N__29016));
    LocalMux I__5300 (
            .O(N__29016),
            .I(N__29011));
    CascadeMux I__5299 (
            .O(N__29015),
            .I(N__29008));
    InMux I__5298 (
            .O(N__29014),
            .I(N__29004));
    Span4Mux_h I__5297 (
            .O(N__29011),
            .I(N__29001));
    InMux I__5296 (
            .O(N__29008),
            .I(N__28996));
    InMux I__5295 (
            .O(N__29007),
            .I(N__28996));
    LocalMux I__5294 (
            .O(N__29004),
            .I(\scaler_3.un2_source_data_0 ));
    Odrv4 I__5293 (
            .O(N__29001),
            .I(\scaler_3.un2_source_data_0 ));
    LocalMux I__5292 (
            .O(N__28996),
            .I(\scaler_3.un2_source_data_0 ));
    InMux I__5291 (
            .O(N__28989),
            .I(N__28985));
    InMux I__5290 (
            .O(N__28988),
            .I(N__28982));
    LocalMux I__5289 (
            .O(N__28985),
            .I(N__28975));
    LocalMux I__5288 (
            .O(N__28982),
            .I(N__28975));
    InMux I__5287 (
            .O(N__28981),
            .I(N__28972));
    CascadeMux I__5286 (
            .O(N__28980),
            .I(N__28969));
    Span4Mux_v I__5285 (
            .O(N__28975),
            .I(N__28966));
    LocalMux I__5284 (
            .O(N__28972),
            .I(N__28963));
    InMux I__5283 (
            .O(N__28969),
            .I(N__28960));
    Odrv4 I__5282 (
            .O(N__28966),
            .I(frame_decoder_OFF3data_0));
    Odrv4 I__5281 (
            .O(N__28963),
            .I(frame_decoder_OFF3data_0));
    LocalMux I__5280 (
            .O(N__28960),
            .I(frame_decoder_OFF3data_0));
    InMux I__5279 (
            .O(N__28953),
            .I(N__28949));
    InMux I__5278 (
            .O(N__28952),
            .I(N__28946));
    LocalMux I__5277 (
            .O(N__28949),
            .I(N__28939));
    LocalMux I__5276 (
            .O(N__28946),
            .I(N__28939));
    InMux I__5275 (
            .O(N__28945),
            .I(N__28936));
    InMux I__5274 (
            .O(N__28944),
            .I(N__28933));
    Span4Mux_v I__5273 (
            .O(N__28939),
            .I(N__28930));
    LocalMux I__5272 (
            .O(N__28936),
            .I(N__28927));
    LocalMux I__5271 (
            .O(N__28933),
            .I(N__28924));
    Odrv4 I__5270 (
            .O(N__28930),
            .I(frame_decoder_CH3data_0));
    Odrv12 I__5269 (
            .O(N__28927),
            .I(frame_decoder_CH3data_0));
    Odrv4 I__5268 (
            .O(N__28924),
            .I(frame_decoder_CH3data_0));
    InMux I__5267 (
            .O(N__28917),
            .I(N__28914));
    LocalMux I__5266 (
            .O(N__28914),
            .I(N__28910));
    InMux I__5265 (
            .O(N__28913),
            .I(N__28906));
    Span4Mux_v I__5264 (
            .O(N__28910),
            .I(N__28903));
    CascadeMux I__5263 (
            .O(N__28909),
            .I(N__28900));
    LocalMux I__5262 (
            .O(N__28906),
            .I(N__28896));
    Span4Mux_v I__5261 (
            .O(N__28903),
            .I(N__28893));
    InMux I__5260 (
            .O(N__28900),
            .I(N__28888));
    InMux I__5259 (
            .O(N__28899),
            .I(N__28888));
    Odrv4 I__5258 (
            .O(N__28896),
            .I(\scaler_4.un2_source_data_0 ));
    Odrv4 I__5257 (
            .O(N__28893),
            .I(\scaler_4.un2_source_data_0 ));
    LocalMux I__5256 (
            .O(N__28888),
            .I(\scaler_4.un2_source_data_0 ));
    CascadeMux I__5255 (
            .O(N__28881),
            .I(\reset_module_System.count_1_1_cascade_ ));
    CascadeMux I__5254 (
            .O(N__28878),
            .I(N__28875));
    InMux I__5253 (
            .O(N__28875),
            .I(N__28871));
    CascadeMux I__5252 (
            .O(N__28874),
            .I(N__28868));
    LocalMux I__5251 (
            .O(N__28871),
            .I(N__28865));
    InMux I__5250 (
            .O(N__28868),
            .I(N__28862));
    Odrv4 I__5249 (
            .O(N__28865),
            .I(\uart_pc.data_AuxZ1Z_0 ));
    LocalMux I__5248 (
            .O(N__28862),
            .I(\uart_pc.data_AuxZ1Z_0 ));
    CascadeMux I__5247 (
            .O(N__28857),
            .I(N__28854));
    InMux I__5246 (
            .O(N__28854),
            .I(N__28850));
    InMux I__5245 (
            .O(N__28853),
            .I(N__28847));
    LocalMux I__5244 (
            .O(N__28850),
            .I(\uart_pc.data_AuxZ1Z_1 ));
    LocalMux I__5243 (
            .O(N__28847),
            .I(\uart_pc.data_AuxZ1Z_1 ));
    CascadeMux I__5242 (
            .O(N__28842),
            .I(N__28838));
    CascadeMux I__5241 (
            .O(N__28841),
            .I(N__28835));
    InMux I__5240 (
            .O(N__28838),
            .I(N__28832));
    InMux I__5239 (
            .O(N__28835),
            .I(N__28829));
    LocalMux I__5238 (
            .O(N__28832),
            .I(\uart_pc.data_AuxZ1Z_2 ));
    LocalMux I__5237 (
            .O(N__28829),
            .I(\uart_pc.data_AuxZ1Z_2 ));
    CascadeMux I__5236 (
            .O(N__28824),
            .I(N__28821));
    InMux I__5235 (
            .O(N__28821),
            .I(N__28818));
    LocalMux I__5234 (
            .O(N__28818),
            .I(N__28814));
    CascadeMux I__5233 (
            .O(N__28817),
            .I(N__28811));
    Span4Mux_v I__5232 (
            .O(N__28814),
            .I(N__28808));
    InMux I__5231 (
            .O(N__28811),
            .I(N__28805));
    Odrv4 I__5230 (
            .O(N__28808),
            .I(\uart_pc.data_AuxZ0Z_4 ));
    LocalMux I__5229 (
            .O(N__28805),
            .I(\uart_pc.data_AuxZ0Z_4 ));
    CascadeMux I__5228 (
            .O(N__28800),
            .I(N__28796));
    CascadeMux I__5227 (
            .O(N__28799),
            .I(N__28793));
    InMux I__5226 (
            .O(N__28796),
            .I(N__28790));
    InMux I__5225 (
            .O(N__28793),
            .I(N__28787));
    LocalMux I__5224 (
            .O(N__28790),
            .I(\uart_pc.data_AuxZ0Z_5 ));
    LocalMux I__5223 (
            .O(N__28787),
            .I(\uart_pc.data_AuxZ0Z_5 ));
    CascadeMux I__5222 (
            .O(N__28782),
            .I(N__28778));
    InMux I__5221 (
            .O(N__28781),
            .I(N__28775));
    InMux I__5220 (
            .O(N__28778),
            .I(N__28772));
    LocalMux I__5219 (
            .O(N__28775),
            .I(\uart_pc.data_AuxZ0Z_6 ));
    LocalMux I__5218 (
            .O(N__28772),
            .I(\uart_pc.data_AuxZ0Z_6 ));
    InMux I__5217 (
            .O(N__28767),
            .I(N__28743));
    InMux I__5216 (
            .O(N__28766),
            .I(N__28743));
    InMux I__5215 (
            .O(N__28765),
            .I(N__28743));
    InMux I__5214 (
            .O(N__28764),
            .I(N__28743));
    InMux I__5213 (
            .O(N__28763),
            .I(N__28743));
    InMux I__5212 (
            .O(N__28762),
            .I(N__28743));
    InMux I__5211 (
            .O(N__28761),
            .I(N__28743));
    InMux I__5210 (
            .O(N__28760),
            .I(N__28743));
    LocalMux I__5209 (
            .O(N__28743),
            .I(N__28740));
    Span4Mux_h I__5208 (
            .O(N__28740),
            .I(N__28737));
    Odrv4 I__5207 (
            .O(N__28737),
            .I(\uart_pc.un1_state_2_0 ));
    InMux I__5206 (
            .O(N__28734),
            .I(N__28729));
    InMux I__5205 (
            .O(N__28733),
            .I(N__28724));
    InMux I__5204 (
            .O(N__28732),
            .I(N__28724));
    LocalMux I__5203 (
            .O(N__28729),
            .I(\pid_alt.error_i_acumm_preregZ0Z_8 ));
    LocalMux I__5202 (
            .O(N__28724),
            .I(\pid_alt.error_i_acumm_preregZ0Z_8 ));
    CascadeMux I__5201 (
            .O(N__28719),
            .I(N__28714));
    CascadeMux I__5200 (
            .O(N__28718),
            .I(N__28711));
    InMux I__5199 (
            .O(N__28717),
            .I(N__28708));
    InMux I__5198 (
            .O(N__28714),
            .I(N__28703));
    InMux I__5197 (
            .O(N__28711),
            .I(N__28703));
    LocalMux I__5196 (
            .O(N__28708),
            .I(\pid_alt.error_i_acumm_preregZ0Z_9 ));
    LocalMux I__5195 (
            .O(N__28703),
            .I(\pid_alt.error_i_acumm_preregZ0Z_9 ));
    InMux I__5194 (
            .O(N__28698),
            .I(N__28691));
    InMux I__5193 (
            .O(N__28697),
            .I(N__28691));
    InMux I__5192 (
            .O(N__28696),
            .I(N__28688));
    LocalMux I__5191 (
            .O(N__28691),
            .I(\pid_alt.error_i_acumm_preregZ0Z_10 ));
    LocalMux I__5190 (
            .O(N__28688),
            .I(\pid_alt.error_i_acumm_preregZ0Z_10 ));
    CascadeMux I__5189 (
            .O(N__28683),
            .I(N__28680));
    InMux I__5188 (
            .O(N__28680),
            .I(N__28677));
    LocalMux I__5187 (
            .O(N__28677),
            .I(\pid_alt.m35_e_2 ));
    CascadeMux I__5186 (
            .O(N__28674),
            .I(N__28669));
    CascadeMux I__5185 (
            .O(N__28673),
            .I(N__28664));
    CascadeMux I__5184 (
            .O(N__28672),
            .I(N__28661));
    InMux I__5183 (
            .O(N__28669),
            .I(N__28649));
    InMux I__5182 (
            .O(N__28668),
            .I(N__28649));
    InMux I__5181 (
            .O(N__28667),
            .I(N__28649));
    InMux I__5180 (
            .O(N__28664),
            .I(N__28649));
    InMux I__5179 (
            .O(N__28661),
            .I(N__28649));
    InMux I__5178 (
            .O(N__28660),
            .I(N__28646));
    LocalMux I__5177 (
            .O(N__28649),
            .I(\pid_alt.N_62_mux ));
    LocalMux I__5176 (
            .O(N__28646),
            .I(\pid_alt.N_62_mux ));
    CascadeMux I__5175 (
            .O(N__28641),
            .I(N__28638));
    InMux I__5174 (
            .O(N__28638),
            .I(N__28633));
    InMux I__5173 (
            .O(N__28637),
            .I(N__28630));
    InMux I__5172 (
            .O(N__28636),
            .I(N__28627));
    LocalMux I__5171 (
            .O(N__28633),
            .I(N__28621));
    LocalMux I__5170 (
            .O(N__28630),
            .I(N__28621));
    LocalMux I__5169 (
            .O(N__28627),
            .I(N__28618));
    InMux I__5168 (
            .O(N__28626),
            .I(N__28615));
    Span4Mux_v I__5167 (
            .O(N__28621),
            .I(N__28608));
    Span4Mux_v I__5166 (
            .O(N__28618),
            .I(N__28608));
    LocalMux I__5165 (
            .O(N__28615),
            .I(N__28608));
    Span4Mux_v I__5164 (
            .O(N__28608),
            .I(N__28605));
    Odrv4 I__5163 (
            .O(N__28605),
            .I(\pid_alt.error_i_acumm7lto5 ));
    CascadeMux I__5162 (
            .O(N__28602),
            .I(N__28599));
    InMux I__5161 (
            .O(N__28599),
            .I(N__28596));
    LocalMux I__5160 (
            .O(N__28596),
            .I(N__28591));
    InMux I__5159 (
            .O(N__28595),
            .I(N__28588));
    InMux I__5158 (
            .O(N__28594),
            .I(N__28585));
    Odrv4 I__5157 (
            .O(N__28591),
            .I(\pid_alt.error_i_acumm7lto12 ));
    LocalMux I__5156 (
            .O(N__28588),
            .I(\pid_alt.error_i_acumm7lto12 ));
    LocalMux I__5155 (
            .O(N__28585),
            .I(\pid_alt.error_i_acumm7lto12 ));
    InMux I__5154 (
            .O(N__28578),
            .I(N__28575));
    LocalMux I__5153 (
            .O(N__28575),
            .I(N__28570));
    InMux I__5152 (
            .O(N__28574),
            .I(N__28565));
    InMux I__5151 (
            .O(N__28573),
            .I(N__28565));
    Odrv4 I__5150 (
            .O(N__28570),
            .I(\pid_alt.N_9_0 ));
    LocalMux I__5149 (
            .O(N__28565),
            .I(\pid_alt.N_9_0 ));
    InMux I__5148 (
            .O(N__28560),
            .I(N__28557));
    LocalMux I__5147 (
            .O(N__28557),
            .I(N__28554));
    Span4Mux_h I__5146 (
            .O(N__28554),
            .I(N__28549));
    InMux I__5145 (
            .O(N__28553),
            .I(N__28544));
    InMux I__5144 (
            .O(N__28552),
            .I(N__28544));
    Odrv4 I__5143 (
            .O(N__28549),
            .I(\pid_alt.error_i_acumm_preregZ0Z_7 ));
    LocalMux I__5142 (
            .O(N__28544),
            .I(\pid_alt.error_i_acumm_preregZ0Z_7 ));
    CascadeMux I__5141 (
            .O(N__28539),
            .I(N__28536));
    InMux I__5140 (
            .O(N__28536),
            .I(N__28530));
    InMux I__5139 (
            .O(N__28535),
            .I(N__28530));
    LocalMux I__5138 (
            .O(N__28530),
            .I(\uart_pc.N_144_1 ));
    CascadeMux I__5137 (
            .O(N__28527),
            .I(N__28524));
    InMux I__5136 (
            .O(N__28524),
            .I(N__28517));
    InMux I__5135 (
            .O(N__28523),
            .I(N__28508));
    InMux I__5134 (
            .O(N__28522),
            .I(N__28508));
    InMux I__5133 (
            .O(N__28521),
            .I(N__28508));
    InMux I__5132 (
            .O(N__28520),
            .I(N__28508));
    LocalMux I__5131 (
            .O(N__28517),
            .I(N__28502));
    LocalMux I__5130 (
            .O(N__28508),
            .I(N__28502));
    InMux I__5129 (
            .O(N__28507),
            .I(N__28499));
    Span4Mux_v I__5128 (
            .O(N__28502),
            .I(N__28494));
    LocalMux I__5127 (
            .O(N__28499),
            .I(N__28494));
    Span4Mux_v I__5126 (
            .O(N__28494),
            .I(N__28491));
    Odrv4 I__5125 (
            .O(N__28491),
            .I(\pid_alt.error_i_acumm7lto4 ));
    InMux I__5124 (
            .O(N__28488),
            .I(N__28484));
    InMux I__5123 (
            .O(N__28487),
            .I(N__28481));
    LocalMux I__5122 (
            .O(N__28484),
            .I(N__28478));
    LocalMux I__5121 (
            .O(N__28481),
            .I(\pid_alt.error_i_acumm_preregZ0Z_2 ));
    Odrv4 I__5120 (
            .O(N__28478),
            .I(\pid_alt.error_i_acumm_preregZ0Z_2 ));
    InMux I__5119 (
            .O(N__28473),
            .I(N__28470));
    LocalMux I__5118 (
            .O(N__28470),
            .I(\pid_alt.m21_e_8 ));
    CascadeMux I__5117 (
            .O(N__28467),
            .I(N__28463));
    CascadeMux I__5116 (
            .O(N__28466),
            .I(N__28460));
    InMux I__5115 (
            .O(N__28463),
            .I(N__28457));
    InMux I__5114 (
            .O(N__28460),
            .I(N__28454));
    LocalMux I__5113 (
            .O(N__28457),
            .I(N__28451));
    LocalMux I__5112 (
            .O(N__28454),
            .I(N__28448));
    Span4Mux_v I__5111 (
            .O(N__28451),
            .I(N__28443));
    Span4Mux_h I__5110 (
            .O(N__28448),
            .I(N__28443));
    Span4Mux_h I__5109 (
            .O(N__28443),
            .I(N__28440));
    Odrv4 I__5108 (
            .O(N__28440),
            .I(\pid_alt.error_i_acumm_preregZ0Z_3 ));
    InMux I__5107 (
            .O(N__28437),
            .I(N__28434));
    LocalMux I__5106 (
            .O(N__28434),
            .I(N__28431));
    Odrv4 I__5105 (
            .O(N__28431),
            .I(\pid_alt.m21_e_2 ));
    CascadeMux I__5104 (
            .O(N__28428),
            .I(\pid_alt.m21_e_10_cascade_ ));
    InMux I__5103 (
            .O(N__28425),
            .I(N__28422));
    LocalMux I__5102 (
            .O(N__28422),
            .I(N__28419));
    Odrv4 I__5101 (
            .O(N__28419),
            .I(\pid_alt.N_138 ));
    InMux I__5100 (
            .O(N__28416),
            .I(N__28413));
    LocalMux I__5099 (
            .O(N__28413),
            .I(N__28410));
    Odrv4 I__5098 (
            .O(N__28410),
            .I(\pid_alt.m35_e_3 ));
    CascadeMux I__5097 (
            .O(N__28407),
            .I(\pid_alt.N_62_mux_cascade_ ));
    InMux I__5096 (
            .O(N__28404),
            .I(N__28392));
    InMux I__5095 (
            .O(N__28403),
            .I(N__28392));
    InMux I__5094 (
            .O(N__28402),
            .I(N__28392));
    InMux I__5093 (
            .O(N__28401),
            .I(N__28392));
    LocalMux I__5092 (
            .O(N__28392),
            .I(\pid_alt.N_129 ));
    InMux I__5091 (
            .O(N__28389),
            .I(N__28385));
    InMux I__5090 (
            .O(N__28388),
            .I(N__28382));
    LocalMux I__5089 (
            .O(N__28385),
            .I(N__28379));
    LocalMux I__5088 (
            .O(N__28382),
            .I(\pid_alt.error_i_acumm_preregZ0Z_1 ));
    Odrv4 I__5087 (
            .O(N__28379),
            .I(\pid_alt.error_i_acumm_preregZ0Z_1 ));
    CascadeMux I__5086 (
            .O(N__28374),
            .I(\pid_alt.m21_e_0_cascade_ ));
    InMux I__5085 (
            .O(N__28371),
            .I(N__28368));
    LocalMux I__5084 (
            .O(N__28368),
            .I(\pid_alt.m21_e_9 ));
    InMux I__5083 (
            .O(N__28365),
            .I(\scaler_4.un2_source_data_0_cry_9 ));
    CascadeMux I__5082 (
            .O(N__28362),
            .I(\pid_alt.un1_reset_1_0_i_cascade_ ));
    CascadeMux I__5081 (
            .O(N__28359),
            .I(N__28356));
    InMux I__5080 (
            .O(N__28356),
            .I(N__28353));
    LocalMux I__5079 (
            .O(N__28353),
            .I(N__28350));
    Odrv4 I__5078 (
            .O(N__28350),
            .I(\scaler_4.un2_source_data_0_cry_1_c_RNO_1 ));
    InMux I__5077 (
            .O(N__28347),
            .I(\scaler_4.un2_source_data_0_cry_1 ));
    CascadeMux I__5076 (
            .O(N__28344),
            .I(N__28341));
    InMux I__5075 (
            .O(N__28341),
            .I(N__28335));
    InMux I__5074 (
            .O(N__28340),
            .I(N__28335));
    LocalMux I__5073 (
            .O(N__28335),
            .I(\scaler_4.un3_source_data_0_cry_1_c_RNI74CL ));
    InMux I__5072 (
            .O(N__28332),
            .I(\scaler_4.un2_source_data_0_cry_2 ));
    CascadeMux I__5071 (
            .O(N__28329),
            .I(N__28326));
    InMux I__5070 (
            .O(N__28326),
            .I(N__28320));
    InMux I__5069 (
            .O(N__28325),
            .I(N__28320));
    LocalMux I__5068 (
            .O(N__28320),
            .I(\scaler_4.un3_source_data_0_cry_2_c_RNIA8DL ));
    InMux I__5067 (
            .O(N__28317),
            .I(\scaler_4.un2_source_data_0_cry_3 ));
    CascadeMux I__5066 (
            .O(N__28314),
            .I(N__28311));
    InMux I__5065 (
            .O(N__28311),
            .I(N__28305));
    InMux I__5064 (
            .O(N__28310),
            .I(N__28305));
    LocalMux I__5063 (
            .O(N__28305),
            .I(\scaler_4.un3_source_data_0_cry_3_c_RNIDCEL ));
    InMux I__5062 (
            .O(N__28302),
            .I(\scaler_4.un2_source_data_0_cry_4 ));
    CascadeMux I__5061 (
            .O(N__28299),
            .I(N__28296));
    InMux I__5060 (
            .O(N__28296),
            .I(N__28290));
    InMux I__5059 (
            .O(N__28295),
            .I(N__28290));
    LocalMux I__5058 (
            .O(N__28290),
            .I(\scaler_4.un3_source_data_0_cry_4_c_RNIGGFL ));
    InMux I__5057 (
            .O(N__28287),
            .I(\scaler_4.un2_source_data_0_cry_5 ));
    CascadeMux I__5056 (
            .O(N__28284),
            .I(N__28281));
    InMux I__5055 (
            .O(N__28281),
            .I(N__28275));
    InMux I__5054 (
            .O(N__28280),
            .I(N__28275));
    LocalMux I__5053 (
            .O(N__28275),
            .I(\scaler_4.un3_source_data_0_cry_5_c_RNIJKGL ));
    InMux I__5052 (
            .O(N__28272),
            .I(\scaler_4.un2_source_data_0_cry_6 ));
    CascadeMux I__5051 (
            .O(N__28269),
            .I(N__28266));
    InMux I__5050 (
            .O(N__28266),
            .I(N__28260));
    InMux I__5049 (
            .O(N__28265),
            .I(N__28260));
    LocalMux I__5048 (
            .O(N__28260),
            .I(\scaler_4.un3_source_data_0_cry_6_c_RNIOUNN ));
    InMux I__5047 (
            .O(N__28257),
            .I(\scaler_4.un2_source_data_0_cry_7 ));
    InMux I__5046 (
            .O(N__28254),
            .I(N__28250));
    InMux I__5045 (
            .O(N__28253),
            .I(N__28247));
    LocalMux I__5044 (
            .O(N__28250),
            .I(\scaler_4.un3_source_data_0_cry_7_c_RNIP0PN ));
    LocalMux I__5043 (
            .O(N__28247),
            .I(\scaler_4.un3_source_data_0_cry_7_c_RNIP0PN ));
    CascadeMux I__5042 (
            .O(N__28242),
            .I(N__28239));
    InMux I__5041 (
            .O(N__28239),
            .I(N__28236));
    LocalMux I__5040 (
            .O(N__28236),
            .I(\scaler_4.un3_source_data_0_cry_8_c_RNIS918 ));
    InMux I__5039 (
            .O(N__28233),
            .I(bfn_12_17_0_));
    CascadeMux I__5038 (
            .O(N__28230),
            .I(N__28227));
    InMux I__5037 (
            .O(N__28227),
            .I(N__28221));
    InMux I__5036 (
            .O(N__28226),
            .I(N__28221));
    LocalMux I__5035 (
            .O(N__28221),
            .I(\scaler_3.un3_source_data_0_cry_1_c_RNI44VK ));
    InMux I__5034 (
            .O(N__28218),
            .I(\scaler_3.un2_source_data_0_cry_2 ));
    CascadeMux I__5033 (
            .O(N__28215),
            .I(N__28212));
    InMux I__5032 (
            .O(N__28212),
            .I(N__28206));
    InMux I__5031 (
            .O(N__28211),
            .I(N__28206));
    LocalMux I__5030 (
            .O(N__28206),
            .I(\scaler_3.un3_source_data_0_cry_2_c_RNI780L ));
    InMux I__5029 (
            .O(N__28203),
            .I(\scaler_3.un2_source_data_0_cry_3 ));
    CascadeMux I__5028 (
            .O(N__28200),
            .I(N__28197));
    InMux I__5027 (
            .O(N__28197),
            .I(N__28191));
    InMux I__5026 (
            .O(N__28196),
            .I(N__28191));
    LocalMux I__5025 (
            .O(N__28191),
            .I(\scaler_3.un3_source_data_0_cry_3_c_RNIAC1L ));
    InMux I__5024 (
            .O(N__28188),
            .I(\scaler_3.un2_source_data_0_cry_4 ));
    CascadeMux I__5023 (
            .O(N__28185),
            .I(N__28182));
    InMux I__5022 (
            .O(N__28182),
            .I(N__28176));
    InMux I__5021 (
            .O(N__28181),
            .I(N__28176));
    LocalMux I__5020 (
            .O(N__28176),
            .I(\scaler_3.un3_source_data_0_cry_4_c_RNIDG2L ));
    InMux I__5019 (
            .O(N__28173),
            .I(\scaler_3.un2_source_data_0_cry_5 ));
    CascadeMux I__5018 (
            .O(N__28170),
            .I(N__28167));
    InMux I__5017 (
            .O(N__28167),
            .I(N__28161));
    InMux I__5016 (
            .O(N__28166),
            .I(N__28161));
    LocalMux I__5015 (
            .O(N__28161),
            .I(\scaler_3.un3_source_data_0_cry_5_c_RNIGK3L ));
    InMux I__5014 (
            .O(N__28158),
            .I(\scaler_3.un2_source_data_0_cry_6 ));
    CascadeMux I__5013 (
            .O(N__28155),
            .I(N__28152));
    InMux I__5012 (
            .O(N__28152),
            .I(N__28146));
    InMux I__5011 (
            .O(N__28151),
            .I(N__28146));
    LocalMux I__5010 (
            .O(N__28146),
            .I(\scaler_3.un3_source_data_0_cry_6_c_RNILUAN ));
    InMux I__5009 (
            .O(N__28143),
            .I(\scaler_3.un2_source_data_0_cry_7 ));
    InMux I__5008 (
            .O(N__28140),
            .I(N__28136));
    InMux I__5007 (
            .O(N__28139),
            .I(N__28133));
    LocalMux I__5006 (
            .O(N__28136),
            .I(\scaler_3.un3_source_data_0_cry_7_c_RNIM0CN ));
    LocalMux I__5005 (
            .O(N__28133),
            .I(\scaler_3.un3_source_data_0_cry_7_c_RNIM0CN ));
    CascadeMux I__5004 (
            .O(N__28128),
            .I(N__28125));
    InMux I__5003 (
            .O(N__28125),
            .I(N__28122));
    LocalMux I__5002 (
            .O(N__28122),
            .I(\scaler_3.un3_source_data_0_cry_8_c_RNIRV25 ));
    InMux I__5001 (
            .O(N__28119),
            .I(bfn_12_15_0_));
    InMux I__5000 (
            .O(N__28116),
            .I(\scaler_3.un2_source_data_0_cry_9 ));
    InMux I__4999 (
            .O(N__28113),
            .I(bfn_12_12_0_));
    InMux I__4998 (
            .O(N__28110),
            .I(\scaler_2.un3_source_data_0_cry_8 ));
    InMux I__4997 (
            .O(N__28107),
            .I(N__28104));
    LocalMux I__4996 (
            .O(N__28104),
            .I(N__28100));
    InMux I__4995 (
            .O(N__28103),
            .I(N__28097));
    Odrv4 I__4994 (
            .O(N__28100),
            .I(frame_decoder_OFF2data_7));
    LocalMux I__4993 (
            .O(N__28097),
            .I(frame_decoder_OFF2data_7));
    InMux I__4992 (
            .O(N__28092),
            .I(N__28088));
    InMux I__4991 (
            .O(N__28091),
            .I(N__28085));
    LocalMux I__4990 (
            .O(N__28088),
            .I(frame_decoder_CH2data_7));
    LocalMux I__4989 (
            .O(N__28085),
            .I(frame_decoder_CH2data_7));
    InMux I__4988 (
            .O(N__28080),
            .I(N__28077));
    LocalMux I__4987 (
            .O(N__28077),
            .I(\scaler_2.N_1227_i_l_ofxZ0 ));
    InMux I__4986 (
            .O(N__28074),
            .I(N__28069));
    CascadeMux I__4985 (
            .O(N__28073),
            .I(N__28062));
    CascadeMux I__4984 (
            .O(N__28072),
            .I(N__28059));
    LocalMux I__4983 (
            .O(N__28069),
            .I(N__28054));
    InMux I__4982 (
            .O(N__28068),
            .I(N__28051));
    CascadeMux I__4981 (
            .O(N__28067),
            .I(N__28048));
    InMux I__4980 (
            .O(N__28066),
            .I(N__28044));
    InMux I__4979 (
            .O(N__28065),
            .I(N__28032));
    InMux I__4978 (
            .O(N__28062),
            .I(N__28032));
    InMux I__4977 (
            .O(N__28059),
            .I(N__28032));
    InMux I__4976 (
            .O(N__28058),
            .I(N__28032));
    InMux I__4975 (
            .O(N__28057),
            .I(N__28032));
    Span4Mux_h I__4974 (
            .O(N__28054),
            .I(N__28027));
    LocalMux I__4973 (
            .O(N__28051),
            .I(N__28027));
    InMux I__4972 (
            .O(N__28048),
            .I(N__28022));
    InMux I__4971 (
            .O(N__28047),
            .I(N__28022));
    LocalMux I__4970 (
            .O(N__28044),
            .I(N__28019));
    InMux I__4969 (
            .O(N__28043),
            .I(N__28016));
    LocalMux I__4968 (
            .O(N__28032),
            .I(N__28011));
    Span4Mux_h I__4967 (
            .O(N__28027),
            .I(N__28011));
    LocalMux I__4966 (
            .O(N__28022),
            .I(N__28008));
    Span4Mux_v I__4965 (
            .O(N__28019),
            .I(N__28005));
    LocalMux I__4964 (
            .O(N__28016),
            .I(N__28002));
    Span4Mux_v I__4963 (
            .O(N__28011),
            .I(N__27999));
    Span4Mux_v I__4962 (
            .O(N__28008),
            .I(N__27992));
    Span4Mux_h I__4961 (
            .O(N__28005),
            .I(N__27992));
    Span4Mux_v I__4960 (
            .O(N__28002),
            .I(N__27992));
    Odrv4 I__4959 (
            .O(N__27999),
            .I(\pid_alt.pid_preregZ0Z_30 ));
    Odrv4 I__4958 (
            .O(N__27992),
            .I(\pid_alt.pid_preregZ0Z_30 ));
    InMux I__4957 (
            .O(N__27987),
            .I(N__27984));
    LocalMux I__4956 (
            .O(N__27984),
            .I(N__27981));
    Span4Mux_h I__4955 (
            .O(N__27981),
            .I(N__27972));
    InMux I__4954 (
            .O(N__27980),
            .I(N__27969));
    InMux I__4953 (
            .O(N__27979),
            .I(N__27958));
    InMux I__4952 (
            .O(N__27978),
            .I(N__27958));
    InMux I__4951 (
            .O(N__27977),
            .I(N__27958));
    InMux I__4950 (
            .O(N__27976),
            .I(N__27958));
    InMux I__4949 (
            .O(N__27975),
            .I(N__27958));
    Odrv4 I__4948 (
            .O(N__27972),
            .I(\pid_alt.N_106 ));
    LocalMux I__4947 (
            .O(N__27969),
            .I(\pid_alt.N_106 ));
    LocalMux I__4946 (
            .O(N__27958),
            .I(\pid_alt.N_106 ));
    InMux I__4945 (
            .O(N__27951),
            .I(N__27948));
    LocalMux I__4944 (
            .O(N__27948),
            .I(N__27944));
    InMux I__4943 (
            .O(N__27947),
            .I(N__27941));
    Span4Mux_h I__4942 (
            .O(N__27944),
            .I(N__27937));
    LocalMux I__4941 (
            .O(N__27941),
            .I(N__27934));
    InMux I__4940 (
            .O(N__27940),
            .I(N__27931));
    Span4Mux_h I__4939 (
            .O(N__27937),
            .I(N__27928));
    Span4Mux_h I__4938 (
            .O(N__27934),
            .I(N__27923));
    LocalMux I__4937 (
            .O(N__27931),
            .I(N__27923));
    Odrv4 I__4936 (
            .O(N__27928),
            .I(\pid_alt.pid_preregZ0Z_9 ));
    Odrv4 I__4935 (
            .O(N__27923),
            .I(\pid_alt.pid_preregZ0Z_9 ));
    CEMux I__4934 (
            .O(N__27918),
            .I(N__27914));
    CEMux I__4933 (
            .O(N__27917),
            .I(N__27909));
    LocalMux I__4932 (
            .O(N__27914),
            .I(N__27906));
    CEMux I__4931 (
            .O(N__27913),
            .I(N__27903));
    CEMux I__4930 (
            .O(N__27912),
            .I(N__27900));
    LocalMux I__4929 (
            .O(N__27909),
            .I(N__27897));
    Span4Mux_h I__4928 (
            .O(N__27906),
            .I(N__27894));
    LocalMux I__4927 (
            .O(N__27903),
            .I(N__27891));
    LocalMux I__4926 (
            .O(N__27900),
            .I(N__27888));
    Span4Mux_v I__4925 (
            .O(N__27897),
            .I(N__27885));
    Odrv4 I__4924 (
            .O(N__27894),
            .I(\pid_alt.N_96_i_1 ));
    Odrv4 I__4923 (
            .O(N__27891),
            .I(\pid_alt.N_96_i_1 ));
    Odrv12 I__4922 (
            .O(N__27888),
            .I(\pid_alt.N_96_i_1 ));
    Odrv4 I__4921 (
            .O(N__27885),
            .I(\pid_alt.N_96_i_1 ));
    SRMux I__4920 (
            .O(N__27876),
            .I(N__27872));
    SRMux I__4919 (
            .O(N__27875),
            .I(N__27869));
    LocalMux I__4918 (
            .O(N__27872),
            .I(N__27866));
    LocalMux I__4917 (
            .O(N__27869),
            .I(N__27859));
    Span4Mux_v I__4916 (
            .O(N__27866),
            .I(N__27856));
    SRMux I__4915 (
            .O(N__27865),
            .I(N__27853));
    SRMux I__4914 (
            .O(N__27864),
            .I(N__27850));
    SRMux I__4913 (
            .O(N__27863),
            .I(N__27847));
    SRMux I__4912 (
            .O(N__27862),
            .I(N__27844));
    Span4Mux_v I__4911 (
            .O(N__27859),
            .I(N__27841));
    Span4Mux_h I__4910 (
            .O(N__27856),
            .I(N__27838));
    LocalMux I__4909 (
            .O(N__27853),
            .I(\pid_alt.un1_reset_0_i ));
    LocalMux I__4908 (
            .O(N__27850),
            .I(\pid_alt.un1_reset_0_i ));
    LocalMux I__4907 (
            .O(N__27847),
            .I(\pid_alt.un1_reset_0_i ));
    LocalMux I__4906 (
            .O(N__27844),
            .I(\pid_alt.un1_reset_0_i ));
    Odrv4 I__4905 (
            .O(N__27841),
            .I(\pid_alt.un1_reset_0_i ));
    Odrv4 I__4904 (
            .O(N__27838),
            .I(\pid_alt.un1_reset_0_i ));
    CascadeMux I__4903 (
            .O(N__27825),
            .I(N__27822));
    InMux I__4902 (
            .O(N__27822),
            .I(N__27819));
    LocalMux I__4901 (
            .O(N__27819),
            .I(N__27816));
    Odrv12 I__4900 (
            .O(N__27816),
            .I(\scaler_3.un2_source_data_0_cry_1_c_RNO_0 ));
    InMux I__4899 (
            .O(N__27813),
            .I(\scaler_3.un2_source_data_0_cry_1 ));
    InMux I__4898 (
            .O(N__27810),
            .I(N__27807));
    LocalMux I__4897 (
            .O(N__27807),
            .I(frame_decoder_CH2data_1));
    CascadeMux I__4896 (
            .O(N__27804),
            .I(N__27801));
    InMux I__4895 (
            .O(N__27801),
            .I(N__27798));
    LocalMux I__4894 (
            .O(N__27798),
            .I(frame_decoder_OFF2data_1));
    InMux I__4893 (
            .O(N__27795),
            .I(\scaler_2.un3_source_data_0_cry_0 ));
    InMux I__4892 (
            .O(N__27792),
            .I(N__27789));
    LocalMux I__4891 (
            .O(N__27789),
            .I(frame_decoder_CH2data_2));
    CascadeMux I__4890 (
            .O(N__27786),
            .I(N__27783));
    InMux I__4889 (
            .O(N__27783),
            .I(N__27780));
    LocalMux I__4888 (
            .O(N__27780),
            .I(frame_decoder_OFF2data_2));
    InMux I__4887 (
            .O(N__27777),
            .I(\scaler_2.un3_source_data_0_cry_1 ));
    InMux I__4886 (
            .O(N__27774),
            .I(N__27771));
    LocalMux I__4885 (
            .O(N__27771),
            .I(frame_decoder_CH2data_3));
    CascadeMux I__4884 (
            .O(N__27768),
            .I(N__27765));
    InMux I__4883 (
            .O(N__27765),
            .I(N__27762));
    LocalMux I__4882 (
            .O(N__27762),
            .I(frame_decoder_OFF2data_3));
    InMux I__4881 (
            .O(N__27759),
            .I(\scaler_2.un3_source_data_0_cry_2 ));
    InMux I__4880 (
            .O(N__27756),
            .I(N__27753));
    LocalMux I__4879 (
            .O(N__27753),
            .I(frame_decoder_CH2data_4));
    CascadeMux I__4878 (
            .O(N__27750),
            .I(N__27747));
    InMux I__4877 (
            .O(N__27747),
            .I(N__27744));
    LocalMux I__4876 (
            .O(N__27744),
            .I(frame_decoder_OFF2data_4));
    InMux I__4875 (
            .O(N__27741),
            .I(\scaler_2.un3_source_data_0_cry_3 ));
    InMux I__4874 (
            .O(N__27738),
            .I(N__27735));
    LocalMux I__4873 (
            .O(N__27735),
            .I(frame_decoder_CH2data_5));
    CascadeMux I__4872 (
            .O(N__27732),
            .I(N__27729));
    InMux I__4871 (
            .O(N__27729),
            .I(N__27726));
    LocalMux I__4870 (
            .O(N__27726),
            .I(frame_decoder_OFF2data_5));
    InMux I__4869 (
            .O(N__27723),
            .I(\scaler_2.un3_source_data_0_cry_4 ));
    InMux I__4868 (
            .O(N__27720),
            .I(N__27717));
    LocalMux I__4867 (
            .O(N__27717),
            .I(frame_decoder_CH2data_6));
    CascadeMux I__4866 (
            .O(N__27714),
            .I(N__27711));
    InMux I__4865 (
            .O(N__27711),
            .I(N__27708));
    LocalMux I__4864 (
            .O(N__27708),
            .I(frame_decoder_OFF2data_6));
    InMux I__4863 (
            .O(N__27705),
            .I(\scaler_2.un3_source_data_0_cry_5 ));
    InMux I__4862 (
            .O(N__27702),
            .I(N__27699));
    LocalMux I__4861 (
            .O(N__27699),
            .I(\scaler_2.un3_source_data_0_axb_7 ));
    InMux I__4860 (
            .O(N__27696),
            .I(\scaler_2.un3_source_data_0_cry_6 ));
    InMux I__4859 (
            .O(N__27693),
            .I(N__27690));
    LocalMux I__4858 (
            .O(N__27690),
            .I(N__27687));
    Span4Mux_h I__4857 (
            .O(N__27687),
            .I(N__27684));
    Odrv4 I__4856 (
            .O(N__27684),
            .I(\uart_drone.data_Auxce_0_5 ));
    InMux I__4855 (
            .O(N__27681),
            .I(N__27678));
    LocalMux I__4854 (
            .O(N__27678),
            .I(N__27674));
    InMux I__4853 (
            .O(N__27677),
            .I(N__27670));
    Span4Mux_h I__4852 (
            .O(N__27674),
            .I(N__27666));
    InMux I__4851 (
            .O(N__27673),
            .I(N__27663));
    LocalMux I__4850 (
            .O(N__27670),
            .I(N__27659));
    InMux I__4849 (
            .O(N__27669),
            .I(N__27656));
    Span4Mux_h I__4848 (
            .O(N__27666),
            .I(N__27646));
    LocalMux I__4847 (
            .O(N__27663),
            .I(N__27646));
    InMux I__4846 (
            .O(N__27662),
            .I(N__27643));
    Span4Mux_v I__4845 (
            .O(N__27659),
            .I(N__27640));
    LocalMux I__4844 (
            .O(N__27656),
            .I(N__27637));
    InMux I__4843 (
            .O(N__27655),
            .I(N__27634));
    InMux I__4842 (
            .O(N__27654),
            .I(N__27631));
    InMux I__4841 (
            .O(N__27653),
            .I(N__27628));
    InMux I__4840 (
            .O(N__27652),
            .I(N__27625));
    InMux I__4839 (
            .O(N__27651),
            .I(N__27622));
    Sp12to4 I__4838 (
            .O(N__27646),
            .I(N__27617));
    LocalMux I__4837 (
            .O(N__27643),
            .I(N__27617));
    Sp12to4 I__4836 (
            .O(N__27640),
            .I(N__27610));
    Sp12to4 I__4835 (
            .O(N__27637),
            .I(N__27603));
    LocalMux I__4834 (
            .O(N__27634),
            .I(N__27603));
    LocalMux I__4833 (
            .O(N__27631),
            .I(N__27603));
    LocalMux I__4832 (
            .O(N__27628),
            .I(N__27600));
    LocalMux I__4831 (
            .O(N__27625),
            .I(N__27595));
    LocalMux I__4830 (
            .O(N__27622),
            .I(N__27595));
    Span12Mux_v I__4829 (
            .O(N__27617),
            .I(N__27592));
    InMux I__4828 (
            .O(N__27616),
            .I(N__27587));
    InMux I__4827 (
            .O(N__27615),
            .I(N__27587));
    InMux I__4826 (
            .O(N__27614),
            .I(N__27582));
    InMux I__4825 (
            .O(N__27613),
            .I(N__27582));
    Odrv12 I__4824 (
            .O(N__27610),
            .I(uart_pc_data_0));
    Odrv12 I__4823 (
            .O(N__27603),
            .I(uart_pc_data_0));
    Odrv4 I__4822 (
            .O(N__27600),
            .I(uart_pc_data_0));
    Odrv4 I__4821 (
            .O(N__27595),
            .I(uart_pc_data_0));
    Odrv12 I__4820 (
            .O(N__27592),
            .I(uart_pc_data_0));
    LocalMux I__4819 (
            .O(N__27587),
            .I(uart_pc_data_0));
    LocalMux I__4818 (
            .O(N__27582),
            .I(uart_pc_data_0));
    CEMux I__4817 (
            .O(N__27567),
            .I(N__27564));
    LocalMux I__4816 (
            .O(N__27564),
            .I(N__27561));
    Span4Mux_v I__4815 (
            .O(N__27561),
            .I(N__27558));
    Odrv4 I__4814 (
            .O(N__27558),
            .I(\Commands_frame_decoder.source_offset2data_1_sqmuxa_0 ));
    CascadeMux I__4813 (
            .O(N__27555),
            .I(N__27548));
    InMux I__4812 (
            .O(N__27554),
            .I(N__27544));
    InMux I__4811 (
            .O(N__27553),
            .I(N__27539));
    InMux I__4810 (
            .O(N__27552),
            .I(N__27539));
    InMux I__4809 (
            .O(N__27551),
            .I(N__27536));
    InMux I__4808 (
            .O(N__27548),
            .I(N__27531));
    InMux I__4807 (
            .O(N__27547),
            .I(N__27531));
    LocalMux I__4806 (
            .O(N__27544),
            .I(\uart_pc.N_143 ));
    LocalMux I__4805 (
            .O(N__27539),
            .I(\uart_pc.N_143 ));
    LocalMux I__4804 (
            .O(N__27536),
            .I(\uart_pc.N_143 ));
    LocalMux I__4803 (
            .O(N__27531),
            .I(\uart_pc.N_143 ));
    CascadeMux I__4802 (
            .O(N__27522),
            .I(\uart_pc.N_145_cascade_ ));
    InMux I__4801 (
            .O(N__27519),
            .I(N__27516));
    LocalMux I__4800 (
            .O(N__27516),
            .I(N__27513));
    Span4Mux_h I__4799 (
            .O(N__27513),
            .I(N__27510));
    Odrv4 I__4798 (
            .O(N__27510),
            .I(\uart_drone.data_Auxce_0_0_4 ));
    InMux I__4797 (
            .O(N__27507),
            .I(N__27504));
    LocalMux I__4796 (
            .O(N__27504),
            .I(N__27501));
    Span4Mux_h I__4795 (
            .O(N__27501),
            .I(N__27498));
    Odrv4 I__4794 (
            .O(N__27498),
            .I(\uart_drone.data_Auxce_0_3 ));
    CascadeMux I__4793 (
            .O(N__27495),
            .I(N__27491));
    InMux I__4792 (
            .O(N__27494),
            .I(N__27487));
    InMux I__4791 (
            .O(N__27491),
            .I(N__27482));
    InMux I__4790 (
            .O(N__27490),
            .I(N__27482));
    LocalMux I__4789 (
            .O(N__27487),
            .I(\uart_pc.timer_CountZ1Z_2 ));
    LocalMux I__4788 (
            .O(N__27482),
            .I(\uart_pc.timer_CountZ1Z_2 ));
    InMux I__4787 (
            .O(N__27477),
            .I(N__27474));
    LocalMux I__4786 (
            .O(N__27474),
            .I(\uart_pc.un1_state_2_0_a3_0 ));
    CascadeMux I__4785 (
            .O(N__27471),
            .I(\uart_pc.N_126_li_cascade_ ));
    CascadeMux I__4784 (
            .O(N__27468),
            .I(N__27464));
    CascadeMux I__4783 (
            .O(N__27467),
            .I(N__27459));
    InMux I__4782 (
            .O(N__27464),
            .I(N__27454));
    InMux I__4781 (
            .O(N__27463),
            .I(N__27454));
    InMux I__4780 (
            .O(N__27462),
            .I(N__27449));
    InMux I__4779 (
            .O(N__27459),
            .I(N__27449));
    LocalMux I__4778 (
            .O(N__27454),
            .I(\uart_pc.timer_Count_0_sqmuxa ));
    LocalMux I__4777 (
            .O(N__27449),
            .I(\uart_pc.timer_Count_0_sqmuxa ));
    InMux I__4776 (
            .O(N__27444),
            .I(N__27441));
    LocalMux I__4775 (
            .O(N__27441),
            .I(\uart_pc.timer_Count_RNO_0Z0Z_3 ));
    CascadeMux I__4774 (
            .O(N__27438),
            .I(\uart_pc.timer_Count_0_sqmuxa_cascade_ ));
    InMux I__4773 (
            .O(N__27435),
            .I(N__27432));
    LocalMux I__4772 (
            .O(N__27432),
            .I(\pid_alt.error_i_acumm_preregZ0Z_15 ));
    CascadeMux I__4771 (
            .O(N__27429),
            .I(\pid_alt.m7_e_4_cascade_ ));
    CascadeMux I__4770 (
            .O(N__27426),
            .I(\pid_alt.N_238_cascade_ ));
    InMux I__4769 (
            .O(N__27423),
            .I(N__27420));
    LocalMux I__4768 (
            .O(N__27420),
            .I(\pid_alt.error_i_acumm_preregZ0Z_18 ));
    CascadeMux I__4767 (
            .O(N__27417),
            .I(N__27414));
    InMux I__4766 (
            .O(N__27414),
            .I(N__27411));
    LocalMux I__4765 (
            .O(N__27411),
            .I(\pid_alt.error_i_acumm_preregZ0Z_19 ));
    InMux I__4764 (
            .O(N__27408),
            .I(N__27405));
    LocalMux I__4763 (
            .O(N__27405),
            .I(\pid_alt.error_i_acumm_preregZ0Z_14 ));
    InMux I__4762 (
            .O(N__27402),
            .I(N__27399));
    LocalMux I__4761 (
            .O(N__27399),
            .I(\pid_alt.error_i_acumm_preregZ0Z_17 ));
    InMux I__4760 (
            .O(N__27396),
            .I(N__27393));
    LocalMux I__4759 (
            .O(N__27393),
            .I(\pid_alt.error_i_acumm_preregZ0Z_20 ));
    InMux I__4758 (
            .O(N__27390),
            .I(bfn_11_17_0_));
    InMux I__4757 (
            .O(N__27387),
            .I(\scaler_4.un3_source_data_0_cry_8 ));
    InMux I__4756 (
            .O(N__27384),
            .I(N__27381));
    LocalMux I__4755 (
            .O(N__27381),
            .I(\scaler_4.un3_source_data_0_axb_7 ));
    InMux I__4754 (
            .O(N__27378),
            .I(N__27372));
    InMux I__4753 (
            .O(N__27377),
            .I(N__27372));
    LocalMux I__4752 (
            .O(N__27372),
            .I(frame_decoder_CH4data_7));
    CascadeMux I__4751 (
            .O(N__27369),
            .I(N__27366));
    InMux I__4750 (
            .O(N__27366),
            .I(N__27360));
    InMux I__4749 (
            .O(N__27365),
            .I(N__27360));
    LocalMux I__4748 (
            .O(N__27360),
            .I(N__27357));
    Odrv4 I__4747 (
            .O(N__27357),
            .I(frame_decoder_OFF4data_7));
    InMux I__4746 (
            .O(N__27354),
            .I(N__27351));
    LocalMux I__4745 (
            .O(N__27351),
            .I(\scaler_4.N_1251_i_l_ofxZ0 ));
    InMux I__4744 (
            .O(N__27348),
            .I(N__27345));
    LocalMux I__4743 (
            .O(N__27345),
            .I(N__27342));
    Span4Mux_h I__4742 (
            .O(N__27342),
            .I(N__27338));
    InMux I__4741 (
            .O(N__27341),
            .I(N__27335));
    Span4Mux_v I__4740 (
            .O(N__27338),
            .I(N__27330));
    LocalMux I__4739 (
            .O(N__27335),
            .I(N__27330));
    Odrv4 I__4738 (
            .O(N__27330),
            .I(\Commands_frame_decoder.source_offset4data_1_sqmuxa ));
    CEMux I__4737 (
            .O(N__27327),
            .I(N__27324));
    LocalMux I__4736 (
            .O(N__27324),
            .I(N__27321));
    Span4Mux_v I__4735 (
            .O(N__27321),
            .I(N__27318));
    Odrv4 I__4734 (
            .O(N__27318),
            .I(\Commands_frame_decoder.source_offset4data_1_sqmuxa_0 ));
    InMux I__4733 (
            .O(N__27315),
            .I(N__27312));
    LocalMux I__4732 (
            .O(N__27312),
            .I(\pid_alt.error_i_acumm_preregZ0Z_16 ));
    InMux I__4731 (
            .O(N__27309),
            .I(N__27306));
    LocalMux I__4730 (
            .O(N__27306),
            .I(frame_decoder_CH4data_1));
    CascadeMux I__4729 (
            .O(N__27303),
            .I(N__27300));
    InMux I__4728 (
            .O(N__27300),
            .I(N__27297));
    LocalMux I__4727 (
            .O(N__27297),
            .I(frame_decoder_OFF4data_1));
    InMux I__4726 (
            .O(N__27294),
            .I(\scaler_4.un3_source_data_0_cry_0 ));
    InMux I__4725 (
            .O(N__27291),
            .I(N__27288));
    LocalMux I__4724 (
            .O(N__27288),
            .I(frame_decoder_CH4data_2));
    CascadeMux I__4723 (
            .O(N__27285),
            .I(N__27282));
    InMux I__4722 (
            .O(N__27282),
            .I(N__27279));
    LocalMux I__4721 (
            .O(N__27279),
            .I(N__27276));
    Odrv12 I__4720 (
            .O(N__27276),
            .I(frame_decoder_OFF4data_2));
    InMux I__4719 (
            .O(N__27273),
            .I(\scaler_4.un3_source_data_0_cry_1 ));
    InMux I__4718 (
            .O(N__27270),
            .I(N__27267));
    LocalMux I__4717 (
            .O(N__27267),
            .I(frame_decoder_CH4data_3));
    CascadeMux I__4716 (
            .O(N__27264),
            .I(N__27261));
    InMux I__4715 (
            .O(N__27261),
            .I(N__27258));
    LocalMux I__4714 (
            .O(N__27258),
            .I(frame_decoder_OFF4data_3));
    InMux I__4713 (
            .O(N__27255),
            .I(\scaler_4.un3_source_data_0_cry_2 ));
    InMux I__4712 (
            .O(N__27252),
            .I(N__27249));
    LocalMux I__4711 (
            .O(N__27249),
            .I(N__27246));
    Span4Mux_h I__4710 (
            .O(N__27246),
            .I(N__27243));
    Span4Mux_v I__4709 (
            .O(N__27243),
            .I(N__27240));
    Odrv4 I__4708 (
            .O(N__27240),
            .I(frame_decoder_CH4data_4));
    CascadeMux I__4707 (
            .O(N__27237),
            .I(N__27234));
    InMux I__4706 (
            .O(N__27234),
            .I(N__27231));
    LocalMux I__4705 (
            .O(N__27231),
            .I(frame_decoder_OFF4data_4));
    InMux I__4704 (
            .O(N__27228),
            .I(\scaler_4.un3_source_data_0_cry_3 ));
    InMux I__4703 (
            .O(N__27225),
            .I(N__27222));
    LocalMux I__4702 (
            .O(N__27222),
            .I(frame_decoder_OFF4data_5));
    CascadeMux I__4701 (
            .O(N__27219),
            .I(N__27216));
    InMux I__4700 (
            .O(N__27216),
            .I(N__27213));
    LocalMux I__4699 (
            .O(N__27213),
            .I(N__27210));
    Span4Mux_h I__4698 (
            .O(N__27210),
            .I(N__27207));
    Span4Mux_h I__4697 (
            .O(N__27207),
            .I(N__27204));
    Odrv4 I__4696 (
            .O(N__27204),
            .I(frame_decoder_CH4data_5));
    InMux I__4695 (
            .O(N__27201),
            .I(\scaler_4.un3_source_data_0_cry_4 ));
    InMux I__4694 (
            .O(N__27198),
            .I(N__27195));
    LocalMux I__4693 (
            .O(N__27195),
            .I(frame_decoder_CH4data_6));
    CascadeMux I__4692 (
            .O(N__27192),
            .I(N__27189));
    InMux I__4691 (
            .O(N__27189),
            .I(N__27186));
    LocalMux I__4690 (
            .O(N__27186),
            .I(frame_decoder_OFF4data_6));
    InMux I__4689 (
            .O(N__27183),
            .I(\scaler_4.un3_source_data_0_cry_5 ));
    InMux I__4688 (
            .O(N__27180),
            .I(\scaler_4.un3_source_data_0_cry_6 ));
    CascadeMux I__4687 (
            .O(N__27177),
            .I(N__27174));
    InMux I__4686 (
            .O(N__27174),
            .I(N__27171));
    LocalMux I__4685 (
            .O(N__27171),
            .I(N__27167));
    CascadeMux I__4684 (
            .O(N__27170),
            .I(N__27163));
    Span4Mux_v I__4683 (
            .O(N__27167),
            .I(N__27160));
    InMux I__4682 (
            .O(N__27166),
            .I(N__27157));
    InMux I__4681 (
            .O(N__27163),
            .I(N__27154));
    Span4Mux_v I__4680 (
            .O(N__27160),
            .I(N__27149));
    LocalMux I__4679 (
            .O(N__27157),
            .I(N__27149));
    LocalMux I__4678 (
            .O(N__27154),
            .I(N__27144));
    Span4Mux_h I__4677 (
            .O(N__27149),
            .I(N__27144));
    Odrv4 I__4676 (
            .O(N__27144),
            .I(\pid_alt.pid_preregZ0Z_7 ));
    CascadeMux I__4675 (
            .O(N__27141),
            .I(N__27137));
    InMux I__4674 (
            .O(N__27140),
            .I(N__27133));
    InMux I__4673 (
            .O(N__27137),
            .I(N__27130));
    CascadeMux I__4672 (
            .O(N__27136),
            .I(N__27127));
    LocalMux I__4671 (
            .O(N__27133),
            .I(N__27124));
    LocalMux I__4670 (
            .O(N__27130),
            .I(N__27121));
    InMux I__4669 (
            .O(N__27127),
            .I(N__27118));
    Span4Mux_h I__4668 (
            .O(N__27124),
            .I(N__27115));
    Span4Mux_h I__4667 (
            .O(N__27121),
            .I(N__27110));
    LocalMux I__4666 (
            .O(N__27118),
            .I(N__27110));
    Odrv4 I__4665 (
            .O(N__27115),
            .I(\pid_alt.pid_preregZ0Z_11 ));
    Odrv4 I__4664 (
            .O(N__27110),
            .I(\pid_alt.pid_preregZ0Z_11 ));
    InMux I__4663 (
            .O(N__27105),
            .I(N__27101));
    InMux I__4662 (
            .O(N__27104),
            .I(N__27098));
    LocalMux I__4661 (
            .O(N__27101),
            .I(N__27094));
    LocalMux I__4660 (
            .O(N__27098),
            .I(N__27091));
    InMux I__4659 (
            .O(N__27097),
            .I(N__27088));
    Span4Mux_v I__4658 (
            .O(N__27094),
            .I(N__27081));
    Span4Mux_h I__4657 (
            .O(N__27091),
            .I(N__27081));
    LocalMux I__4656 (
            .O(N__27088),
            .I(N__27081));
    Odrv4 I__4655 (
            .O(N__27081),
            .I(\pid_alt.pid_preregZ0Z_10 ));
    CascadeMux I__4654 (
            .O(N__27078),
            .I(N__27075));
    InMux I__4653 (
            .O(N__27075),
            .I(N__27072));
    LocalMux I__4652 (
            .O(N__27072),
            .I(N__27069));
    Odrv4 I__4651 (
            .O(N__27069),
            .I(\pid_alt.source_pid_1_sqmuxa_0_a2_2_4 ));
    InMux I__4650 (
            .O(N__27066),
            .I(N__27063));
    LocalMux I__4649 (
            .O(N__27063),
            .I(N__27060));
    Span4Mux_v I__4648 (
            .O(N__27060),
            .I(N__27056));
    InMux I__4647 (
            .O(N__27059),
            .I(N__27053));
    Span4Mux_v I__4646 (
            .O(N__27056),
            .I(N__27050));
    LocalMux I__4645 (
            .O(N__27053),
            .I(\Commands_frame_decoder.stateZ0Z_9 ));
    Odrv4 I__4644 (
            .O(N__27050),
            .I(\Commands_frame_decoder.stateZ0Z_9 ));
    InMux I__4643 (
            .O(N__27045),
            .I(N__27036));
    CascadeMux I__4642 (
            .O(N__27044),
            .I(N__27032));
    CascadeMux I__4641 (
            .O(N__27043),
            .I(N__27029));
    InMux I__4640 (
            .O(N__27042),
            .I(N__27023));
    InMux I__4639 (
            .O(N__27041),
            .I(N__27017));
    InMux I__4638 (
            .O(N__27040),
            .I(N__27014));
    InMux I__4637 (
            .O(N__27039),
            .I(N__27011));
    LocalMux I__4636 (
            .O(N__27036),
            .I(N__27005));
    InMux I__4635 (
            .O(N__27035),
            .I(N__27000));
    InMux I__4634 (
            .O(N__27032),
            .I(N__27000));
    InMux I__4633 (
            .O(N__27029),
            .I(N__26993));
    InMux I__4632 (
            .O(N__27028),
            .I(N__26993));
    InMux I__4631 (
            .O(N__27027),
            .I(N__26990));
    CascadeMux I__4630 (
            .O(N__27026),
            .I(N__26986));
    LocalMux I__4629 (
            .O(N__27023),
            .I(N__26983));
    InMux I__4628 (
            .O(N__27022),
            .I(N__26976));
    InMux I__4627 (
            .O(N__27021),
            .I(N__26976));
    InMux I__4626 (
            .O(N__27020),
            .I(N__26976));
    LocalMux I__4625 (
            .O(N__27017),
            .I(N__26973));
    LocalMux I__4624 (
            .O(N__27014),
            .I(N__26969));
    LocalMux I__4623 (
            .O(N__27011),
            .I(N__26966));
    InMux I__4622 (
            .O(N__27010),
            .I(N__26959));
    InMux I__4621 (
            .O(N__27009),
            .I(N__26959));
    InMux I__4620 (
            .O(N__27008),
            .I(N__26959));
    Span4Mux_v I__4619 (
            .O(N__27005),
            .I(N__26954));
    LocalMux I__4618 (
            .O(N__27000),
            .I(N__26954));
    CascadeMux I__4617 (
            .O(N__26999),
            .I(N__26950));
    InMux I__4616 (
            .O(N__26998),
            .I(N__26947));
    LocalMux I__4615 (
            .O(N__26993),
            .I(N__26942));
    LocalMux I__4614 (
            .O(N__26990),
            .I(N__26942));
    InMux I__4613 (
            .O(N__26989),
            .I(N__26937));
    InMux I__4612 (
            .O(N__26986),
            .I(N__26937));
    Span4Mux_v I__4611 (
            .O(N__26983),
            .I(N__26934));
    LocalMux I__4610 (
            .O(N__26976),
            .I(N__26929));
    Span4Mux_v I__4609 (
            .O(N__26973),
            .I(N__26929));
    InMux I__4608 (
            .O(N__26972),
            .I(N__26926));
    Span4Mux_h I__4607 (
            .O(N__26969),
            .I(N__26917));
    Span4Mux_v I__4606 (
            .O(N__26966),
            .I(N__26917));
    LocalMux I__4605 (
            .O(N__26959),
            .I(N__26917));
    Span4Mux_v I__4604 (
            .O(N__26954),
            .I(N__26917));
    InMux I__4603 (
            .O(N__26953),
            .I(N__26912));
    InMux I__4602 (
            .O(N__26950),
            .I(N__26912));
    LocalMux I__4601 (
            .O(N__26947),
            .I(uart_pc_data_rdy));
    Odrv12 I__4600 (
            .O(N__26942),
            .I(uart_pc_data_rdy));
    LocalMux I__4599 (
            .O(N__26937),
            .I(uart_pc_data_rdy));
    Odrv4 I__4598 (
            .O(N__26934),
            .I(uart_pc_data_rdy));
    Odrv4 I__4597 (
            .O(N__26929),
            .I(uart_pc_data_rdy));
    LocalMux I__4596 (
            .O(N__26926),
            .I(uart_pc_data_rdy));
    Odrv4 I__4595 (
            .O(N__26917),
            .I(uart_pc_data_rdy));
    LocalMux I__4594 (
            .O(N__26912),
            .I(uart_pc_data_rdy));
    InMux I__4593 (
            .O(N__26895),
            .I(N__26892));
    LocalMux I__4592 (
            .O(N__26892),
            .I(N__26889));
    Odrv4 I__4591 (
            .O(N__26889),
            .I(frame_decoder_CH3data_2));
    CascadeMux I__4590 (
            .O(N__26886),
            .I(N__26883));
    InMux I__4589 (
            .O(N__26883),
            .I(N__26880));
    LocalMux I__4588 (
            .O(N__26880),
            .I(frame_decoder_OFF3data_2));
    InMux I__4587 (
            .O(N__26877),
            .I(\scaler_3.un3_source_data_0_cry_1 ));
    InMux I__4586 (
            .O(N__26874),
            .I(N__26871));
    LocalMux I__4585 (
            .O(N__26871),
            .I(N__26868));
    Odrv4 I__4584 (
            .O(N__26868),
            .I(frame_decoder_CH3data_3));
    CascadeMux I__4583 (
            .O(N__26865),
            .I(N__26862));
    InMux I__4582 (
            .O(N__26862),
            .I(N__26859));
    LocalMux I__4581 (
            .O(N__26859),
            .I(frame_decoder_OFF3data_3));
    InMux I__4580 (
            .O(N__26856),
            .I(\scaler_3.un3_source_data_0_cry_2 ));
    InMux I__4579 (
            .O(N__26853),
            .I(N__26850));
    LocalMux I__4578 (
            .O(N__26850),
            .I(N__26847));
    Span4Mux_h I__4577 (
            .O(N__26847),
            .I(N__26844));
    Odrv4 I__4576 (
            .O(N__26844),
            .I(frame_decoder_CH3data_4));
    CascadeMux I__4575 (
            .O(N__26841),
            .I(N__26838));
    InMux I__4574 (
            .O(N__26838),
            .I(N__26835));
    LocalMux I__4573 (
            .O(N__26835),
            .I(frame_decoder_OFF3data_4));
    InMux I__4572 (
            .O(N__26832),
            .I(\scaler_3.un3_source_data_0_cry_3 ));
    InMux I__4571 (
            .O(N__26829),
            .I(N__26826));
    LocalMux I__4570 (
            .O(N__26826),
            .I(N__26823));
    Span4Mux_h I__4569 (
            .O(N__26823),
            .I(N__26820));
    Odrv4 I__4568 (
            .O(N__26820),
            .I(frame_decoder_CH3data_5));
    CascadeMux I__4567 (
            .O(N__26817),
            .I(N__26814));
    InMux I__4566 (
            .O(N__26814),
            .I(N__26811));
    LocalMux I__4565 (
            .O(N__26811),
            .I(N__26808));
    Odrv4 I__4564 (
            .O(N__26808),
            .I(frame_decoder_OFF3data_5));
    InMux I__4563 (
            .O(N__26805),
            .I(\scaler_3.un3_source_data_0_cry_4 ));
    InMux I__4562 (
            .O(N__26802),
            .I(N__26799));
    LocalMux I__4561 (
            .O(N__26799),
            .I(N__26796));
    Span4Mux_v I__4560 (
            .O(N__26796),
            .I(N__26793));
    Odrv4 I__4559 (
            .O(N__26793),
            .I(frame_decoder_CH3data_6));
    CascadeMux I__4558 (
            .O(N__26790),
            .I(N__26787));
    InMux I__4557 (
            .O(N__26787),
            .I(N__26784));
    LocalMux I__4556 (
            .O(N__26784),
            .I(frame_decoder_OFF3data_6));
    InMux I__4555 (
            .O(N__26781),
            .I(\scaler_3.un3_source_data_0_cry_5 ));
    InMux I__4554 (
            .O(N__26778),
            .I(N__26775));
    LocalMux I__4553 (
            .O(N__26775),
            .I(N__26772));
    Odrv12 I__4552 (
            .O(N__26772),
            .I(\scaler_3.un3_source_data_0_axb_7 ));
    InMux I__4551 (
            .O(N__26769),
            .I(\scaler_3.un3_source_data_0_cry_6 ));
    InMux I__4550 (
            .O(N__26766),
            .I(N__26763));
    LocalMux I__4549 (
            .O(N__26763),
            .I(N__26760));
    Odrv12 I__4548 (
            .O(N__26760),
            .I(\scaler_3.N_1239_i_l_ofxZ0 ));
    InMux I__4547 (
            .O(N__26757),
            .I(bfn_11_14_0_));
    InMux I__4546 (
            .O(N__26754),
            .I(\scaler_3.un3_source_data_0_cry_8 ));
    CEMux I__4545 (
            .O(N__26751),
            .I(N__26748));
    LocalMux I__4544 (
            .O(N__26748),
            .I(N__26745));
    Sp12to4 I__4543 (
            .O(N__26745),
            .I(N__26741));
    CEMux I__4542 (
            .O(N__26744),
            .I(N__26738));
    Odrv12 I__4541 (
            .O(N__26741),
            .I(\Commands_frame_decoder.source_offset3data_1_sqmuxa_0 ));
    LocalMux I__4540 (
            .O(N__26738),
            .I(\Commands_frame_decoder.source_offset3data_1_sqmuxa_0 ));
    InMux I__4539 (
            .O(N__26733),
            .I(N__26730));
    LocalMux I__4538 (
            .O(N__26730),
            .I(frame_decoder_OFF3data_1));
    CascadeMux I__4537 (
            .O(N__26727),
            .I(N__26724));
    InMux I__4536 (
            .O(N__26724),
            .I(N__26721));
    LocalMux I__4535 (
            .O(N__26721),
            .I(N__26718));
    Span4Mux_v I__4534 (
            .O(N__26718),
            .I(N__26715));
    Odrv4 I__4533 (
            .O(N__26715),
            .I(frame_decoder_CH3data_1));
    InMux I__4532 (
            .O(N__26712),
            .I(\scaler_3.un3_source_data_0_cry_0 ));
    InMux I__4531 (
            .O(N__26709),
            .I(N__26705));
    InMux I__4530 (
            .O(N__26708),
            .I(N__26702));
    LocalMux I__4529 (
            .O(N__26705),
            .I(N__26699));
    LocalMux I__4528 (
            .O(N__26702),
            .I(N__26696));
    Span4Mux_h I__4527 (
            .O(N__26699),
            .I(N__26693));
    Span4Mux_h I__4526 (
            .O(N__26696),
            .I(N__26690));
    Odrv4 I__4525 (
            .O(N__26693),
            .I(frame_decoder_OFF3data_7));
    Odrv4 I__4524 (
            .O(N__26690),
            .I(frame_decoder_OFF3data_7));
    InMux I__4523 (
            .O(N__26685),
            .I(N__26681));
    InMux I__4522 (
            .O(N__26684),
            .I(N__26678));
    LocalMux I__4521 (
            .O(N__26681),
            .I(N__26675));
    LocalMux I__4520 (
            .O(N__26678),
            .I(frame_decoder_CH3data_7));
    Odrv4 I__4519 (
            .O(N__26675),
            .I(frame_decoder_CH3data_7));
    CEMux I__4518 (
            .O(N__26670),
            .I(N__26667));
    LocalMux I__4517 (
            .O(N__26667),
            .I(N__26664));
    Span4Mux_h I__4516 (
            .O(N__26664),
            .I(N__26661));
    Span4Mux_h I__4515 (
            .O(N__26661),
            .I(N__26658));
    Odrv4 I__4514 (
            .O(N__26658),
            .I(\Commands_frame_decoder.source_CH2data_1_sqmuxa_0 ));
    CascadeMux I__4513 (
            .O(N__26655),
            .I(N__26651));
    InMux I__4512 (
            .O(N__26654),
            .I(N__26646));
    InMux I__4511 (
            .O(N__26651),
            .I(N__26639));
    InMux I__4510 (
            .O(N__26650),
            .I(N__26639));
    InMux I__4509 (
            .O(N__26649),
            .I(N__26639));
    LocalMux I__4508 (
            .O(N__26646),
            .I(\Commands_frame_decoder.countZ0Z_0 ));
    LocalMux I__4507 (
            .O(N__26639),
            .I(\Commands_frame_decoder.countZ0Z_0 ));
    InMux I__4506 (
            .O(N__26634),
            .I(N__26629));
    InMux I__4505 (
            .O(N__26633),
            .I(N__26624));
    InMux I__4504 (
            .O(N__26632),
            .I(N__26624));
    LocalMux I__4503 (
            .O(N__26629),
            .I(\Commands_frame_decoder.countZ0Z_1 ));
    LocalMux I__4502 (
            .O(N__26624),
            .I(\Commands_frame_decoder.countZ0Z_1 ));
    SRMux I__4501 (
            .O(N__26619),
            .I(N__26616));
    LocalMux I__4500 (
            .O(N__26616),
            .I(N__26613));
    Span4Mux_v I__4499 (
            .O(N__26613),
            .I(N__26610));
    Sp12to4 I__4498 (
            .O(N__26610),
            .I(N__26607));
    Odrv12 I__4497 (
            .O(N__26607),
            .I(\uart_drone.timer_Count_RNIES9Q1Z0Z_2 ));
    CascadeMux I__4496 (
            .O(N__26604),
            .I(\uart_drone.timer_Count_RNIES9Q1Z0Z_2_cascade_ ));
    CEMux I__4495 (
            .O(N__26601),
            .I(N__26598));
    LocalMux I__4494 (
            .O(N__26598),
            .I(N__26595));
    Span4Mux_h I__4493 (
            .O(N__26595),
            .I(N__26592));
    Span4Mux_h I__4492 (
            .O(N__26592),
            .I(N__26589));
    Odrv4 I__4491 (
            .O(N__26589),
            .I(\uart_drone.data_rdyc_1_0 ));
    InMux I__4490 (
            .O(N__26586),
            .I(N__26581));
    InMux I__4489 (
            .O(N__26585),
            .I(N__26578));
    InMux I__4488 (
            .O(N__26584),
            .I(N__26575));
    LocalMux I__4487 (
            .O(N__26581),
            .I(N__26569));
    LocalMux I__4486 (
            .O(N__26578),
            .I(N__26569));
    LocalMux I__4485 (
            .O(N__26575),
            .I(N__26566));
    InMux I__4484 (
            .O(N__26574),
            .I(N__26563));
    Odrv4 I__4483 (
            .O(N__26569),
            .I(\uart_pc.data_rdyc_1 ));
    Odrv12 I__4482 (
            .O(N__26566),
            .I(\uart_pc.data_rdyc_1 ));
    LocalMux I__4481 (
            .O(N__26563),
            .I(\uart_pc.data_rdyc_1 ));
    InMux I__4480 (
            .O(N__26556),
            .I(N__26553));
    LocalMux I__4479 (
            .O(N__26553),
            .I(\uart_drone.data_Auxce_0_0_0 ));
    InMux I__4478 (
            .O(N__26550),
            .I(N__26547));
    LocalMux I__4477 (
            .O(N__26547),
            .I(\uart_drone.data_Auxce_0_1 ));
    InMux I__4476 (
            .O(N__26544),
            .I(N__26541));
    LocalMux I__4475 (
            .O(N__26541),
            .I(\uart_pc.timer_Count_RNO_0Z0Z_4 ));
    CascadeMux I__4474 (
            .O(N__26538),
            .I(N__26532));
    InMux I__4473 (
            .O(N__26537),
            .I(N__26529));
    InMux I__4472 (
            .O(N__26536),
            .I(N__26526));
    InMux I__4471 (
            .O(N__26535),
            .I(N__26521));
    InMux I__4470 (
            .O(N__26532),
            .I(N__26521));
    LocalMux I__4469 (
            .O(N__26529),
            .I(\uart_pc.timer_CountZ0Z_0 ));
    LocalMux I__4468 (
            .O(N__26526),
            .I(\uart_pc.timer_CountZ0Z_0 ));
    LocalMux I__4467 (
            .O(N__26521),
            .I(\uart_pc.timer_CountZ0Z_0 ));
    CascadeMux I__4466 (
            .O(N__26514),
            .I(\uart_pc.timer_Count_RNO_0Z0Z_1_cascade_ ));
    InMux I__4465 (
            .O(N__26511),
            .I(N__26507));
    InMux I__4464 (
            .O(N__26510),
            .I(N__26504));
    LocalMux I__4463 (
            .O(N__26507),
            .I(\uart_pc.timer_CountZ1Z_1 ));
    LocalMux I__4462 (
            .O(N__26504),
            .I(\uart_pc.timer_CountZ1Z_1 ));
    InMux I__4461 (
            .O(N__26499),
            .I(N__26493));
    InMux I__4460 (
            .O(N__26498),
            .I(N__26493));
    LocalMux I__4459 (
            .O(N__26493),
            .I(N__26490));
    Odrv4 I__4458 (
            .O(N__26490),
            .I(\Commands_frame_decoder.state_ns_0_a4_0_0Z0Z_1 ));
    CascadeMux I__4457 (
            .O(N__26487),
            .I(\Commands_frame_decoder.state_ns_i_a4_2_0_0_cascade_ ));
    InMux I__4456 (
            .O(N__26484),
            .I(N__26477));
    InMux I__4455 (
            .O(N__26483),
            .I(N__26477));
    InMux I__4454 (
            .O(N__26482),
            .I(N__26473));
    LocalMux I__4453 (
            .O(N__26477),
            .I(N__26470));
    InMux I__4452 (
            .O(N__26476),
            .I(N__26467));
    LocalMux I__4451 (
            .O(N__26473),
            .I(N__26459));
    Span4Mux_v I__4450 (
            .O(N__26470),
            .I(N__26459));
    LocalMux I__4449 (
            .O(N__26467),
            .I(N__26459));
    InMux I__4448 (
            .O(N__26466),
            .I(N__26456));
    Span4Mux_h I__4447 (
            .O(N__26459),
            .I(N__26453));
    LocalMux I__4446 (
            .O(N__26456),
            .I(\Commands_frame_decoder.stateZ0Z_12 ));
    Odrv4 I__4445 (
            .O(N__26453),
            .I(\Commands_frame_decoder.stateZ0Z_12 ));
    InMux I__4444 (
            .O(N__26448),
            .I(N__26445));
    LocalMux I__4443 (
            .O(N__26445),
            .I(N__26441));
    InMux I__4442 (
            .O(N__26444),
            .I(N__26438));
    Span4Mux_v I__4441 (
            .O(N__26441),
            .I(N__26433));
    LocalMux I__4440 (
            .O(N__26438),
            .I(N__26433));
    Odrv4 I__4439 (
            .O(N__26433),
            .I(\Commands_frame_decoder.N_330 ));
    InMux I__4438 (
            .O(N__26430),
            .I(N__26427));
    LocalMux I__4437 (
            .O(N__26427),
            .I(N__26424));
    Odrv4 I__4436 (
            .O(N__26424),
            .I(\Commands_frame_decoder.state_ns_i_a4_2_0_0 ));
    InMux I__4435 (
            .O(N__26421),
            .I(N__26418));
    LocalMux I__4434 (
            .O(N__26418),
            .I(\uart_pc_sync.aux_3__0_Z0Z_0 ));
    InMux I__4433 (
            .O(N__26415),
            .I(\uart_pc.un4_timer_Count_1_cry_1 ));
    InMux I__4432 (
            .O(N__26412),
            .I(\uart_pc.un4_timer_Count_1_cry_2 ));
    InMux I__4431 (
            .O(N__26409),
            .I(\uart_pc.un4_timer_Count_1_cry_3 ));
    InMux I__4430 (
            .O(N__26406),
            .I(N__26403));
    LocalMux I__4429 (
            .O(N__26403),
            .I(\uart_pc.timer_Count_RNO_0Z0Z_2 ));
    CEMux I__4428 (
            .O(N__26400),
            .I(N__26397));
    LocalMux I__4427 (
            .O(N__26397),
            .I(N__26393));
    CEMux I__4426 (
            .O(N__26396),
            .I(N__26390));
    Span4Mux_h I__4425 (
            .O(N__26393),
            .I(N__26387));
    LocalMux I__4424 (
            .O(N__26390),
            .I(N__26384));
    Span4Mux_h I__4423 (
            .O(N__26387),
            .I(N__26378));
    Span4Mux_v I__4422 (
            .O(N__26384),
            .I(N__26378));
    CEMux I__4421 (
            .O(N__26383),
            .I(N__26375));
    Span4Mux_v I__4420 (
            .O(N__26378),
            .I(N__26372));
    LocalMux I__4419 (
            .O(N__26375),
            .I(N__26369));
    Span4Mux_v I__4418 (
            .O(N__26372),
            .I(N__26364));
    Span4Mux_v I__4417 (
            .O(N__26369),
            .I(N__26364));
    Odrv4 I__4416 (
            .O(N__26364),
            .I(\Commands_frame_decoder.source_CH4data_1_sqmuxa_0 ));
    InMux I__4415 (
            .O(N__26361),
            .I(N__26358));
    LocalMux I__4414 (
            .O(N__26358),
            .I(N__26355));
    Odrv4 I__4413 (
            .O(N__26355),
            .I(\Commands_frame_decoder.source_CH1data8lt7_0 ));
    InMux I__4412 (
            .O(N__26352),
            .I(N__26349));
    LocalMux I__4411 (
            .O(N__26349),
            .I(N__26346));
    Span4Mux_v I__4410 (
            .O(N__26346),
            .I(N__26342));
    InMux I__4409 (
            .O(N__26345),
            .I(N__26339));
    Span4Mux_h I__4408 (
            .O(N__26342),
            .I(N__26336));
    LocalMux I__4407 (
            .O(N__26339),
            .I(N__26333));
    Odrv4 I__4406 (
            .O(N__26336),
            .I(\pid_alt.error_d_reg_prev_esr_RNIF2611_0Z0Z_7 ));
    Odrv4 I__4405 (
            .O(N__26333),
            .I(\pid_alt.error_d_reg_prev_esr_RNIF2611_0Z0Z_7 ));
    InMux I__4404 (
            .O(N__26328),
            .I(N__26324));
    InMux I__4403 (
            .O(N__26327),
            .I(N__26321));
    LocalMux I__4402 (
            .O(N__26324),
            .I(\pid_alt.error_d_reg_prev_esr_RNICV511Z0Z_6 ));
    LocalMux I__4401 (
            .O(N__26321),
            .I(\pid_alt.error_d_reg_prev_esr_RNICV511Z0Z_6 ));
    InMux I__4400 (
            .O(N__26316),
            .I(N__26312));
    CascadeMux I__4399 (
            .O(N__26315),
            .I(N__26309));
    LocalMux I__4398 (
            .O(N__26312),
            .I(N__26306));
    InMux I__4397 (
            .O(N__26309),
            .I(N__26303));
    Span4Mux_v I__4396 (
            .O(N__26306),
            .I(N__26300));
    LocalMux I__4395 (
            .O(N__26303),
            .I(N__26297));
    Span4Mux_h I__4394 (
            .O(N__26300),
            .I(N__26294));
    Span4Mux_v I__4393 (
            .O(N__26297),
            .I(N__26291));
    Odrv4 I__4392 (
            .O(N__26294),
            .I(\pid_alt.error_d_reg_prev_esr_RNIUI2T2Z0Z_6 ));
    Odrv4 I__4391 (
            .O(N__26291),
            .I(\pid_alt.error_d_reg_prev_esr_RNIUI2T2Z0Z_6 ));
    InMux I__4390 (
            .O(N__26286),
            .I(N__26283));
    LocalMux I__4389 (
            .O(N__26283),
            .I(\pid_alt.error_d_reg_prev_esr_RNIOOKM_0Z0Z_24 ));
    InMux I__4388 (
            .O(N__26280),
            .I(N__26276));
    InMux I__4387 (
            .O(N__26279),
            .I(N__26273));
    LocalMux I__4386 (
            .O(N__26276),
            .I(N__26270));
    LocalMux I__4385 (
            .O(N__26273),
            .I(N__26267));
    Span4Mux_h I__4384 (
            .O(N__26270),
            .I(N__26264));
    Span4Mux_v I__4383 (
            .O(N__26267),
            .I(N__26261));
    Span4Mux_h I__4382 (
            .O(N__26264),
            .I(N__26258));
    Span4Mux_h I__4381 (
            .O(N__26261),
            .I(N__26255));
    Odrv4 I__4380 (
            .O(N__26258),
            .I(\pid_alt.error_d_reg_prev_esr_RNIMMKMZ0Z_23 ));
    Odrv4 I__4379 (
            .O(N__26255),
            .I(\pid_alt.error_d_reg_prev_esr_RNIMMKMZ0Z_23 ));
    CascadeMux I__4378 (
            .O(N__26250),
            .I(N__26247));
    InMux I__4377 (
            .O(N__26247),
            .I(N__26244));
    LocalMux I__4376 (
            .O(N__26244),
            .I(N__26240));
    InMux I__4375 (
            .O(N__26243),
            .I(N__26237));
    Span4Mux_h I__4374 (
            .O(N__26240),
            .I(N__26234));
    LocalMux I__4373 (
            .O(N__26237),
            .I(N__26231));
    Span4Mux_h I__4372 (
            .O(N__26234),
            .I(N__26228));
    Span4Mux_h I__4371 (
            .O(N__26231),
            .I(N__26225));
    Odrv4 I__4370 (
            .O(N__26228),
            .I(\pid_alt.error_d_reg_prev_esr_RNI6BU12Z0Z_22 ));
    Odrv4 I__4369 (
            .O(N__26225),
            .I(\pid_alt.error_d_reg_prev_esr_RNI6BU12Z0Z_22 ));
    CascadeMux I__4368 (
            .O(N__26220),
            .I(N__26217));
    InMux I__4367 (
            .O(N__26217),
            .I(N__26214));
    LocalMux I__4366 (
            .O(N__26214),
            .I(N__26211));
    Span4Mux_h I__4365 (
            .O(N__26211),
            .I(N__26208));
    Odrv4 I__4364 (
            .O(N__26208),
            .I(\pid_alt.error_d_reg_prev_esr_RNIGQS34Z0Z_23 ));
    InMux I__4363 (
            .O(N__26205),
            .I(N__26202));
    LocalMux I__4362 (
            .O(N__26202),
            .I(N__26197));
    InMux I__4361 (
            .O(N__26201),
            .I(N__26194));
    InMux I__4360 (
            .O(N__26200),
            .I(N__26191));
    Span4Mux_v I__4359 (
            .O(N__26197),
            .I(N__26187));
    LocalMux I__4358 (
            .O(N__26194),
            .I(N__26184));
    LocalMux I__4357 (
            .O(N__26191),
            .I(N__26181));
    InMux I__4356 (
            .O(N__26190),
            .I(N__26178));
    Span4Mux_v I__4355 (
            .O(N__26187),
            .I(N__26175));
    Span12Mux_v I__4354 (
            .O(N__26184),
            .I(N__26172));
    Span4Mux_h I__4353 (
            .O(N__26181),
            .I(N__26169));
    LocalMux I__4352 (
            .O(N__26178),
            .I(N__26166));
    Odrv4 I__4351 (
            .O(N__26175),
            .I(uart_drone_data_3));
    Odrv12 I__4350 (
            .O(N__26172),
            .I(uart_drone_data_3));
    Odrv4 I__4349 (
            .O(N__26169),
            .I(uart_drone_data_3));
    Odrv4 I__4348 (
            .O(N__26166),
            .I(uart_drone_data_3));
    InMux I__4347 (
            .O(N__26157),
            .I(N__26154));
    LocalMux I__4346 (
            .O(N__26154),
            .I(N__26151));
    Odrv4 I__4345 (
            .O(N__26151),
            .I(\dron_frame_decoder_1.drone_altitude_11 ));
    CEMux I__4344 (
            .O(N__26148),
            .I(N__26144));
    CEMux I__4343 (
            .O(N__26147),
            .I(N__26141));
    LocalMux I__4342 (
            .O(N__26144),
            .I(N__26138));
    LocalMux I__4341 (
            .O(N__26141),
            .I(N__26135));
    Span4Mux_h I__4340 (
            .O(N__26138),
            .I(N__26132));
    Span4Mux_h I__4339 (
            .O(N__26135),
            .I(N__26129));
    Span4Mux_v I__4338 (
            .O(N__26132),
            .I(N__26126));
    Span4Mux_h I__4337 (
            .O(N__26129),
            .I(N__26123));
    Odrv4 I__4336 (
            .O(N__26126),
            .I(\dron_frame_decoder_1.N_384_0 ));
    Odrv4 I__4335 (
            .O(N__26123),
            .I(\dron_frame_decoder_1.N_384_0 ));
    CascadeMux I__4334 (
            .O(N__26118),
            .I(N__26115));
    InMux I__4333 (
            .O(N__26115),
            .I(N__26111));
    InMux I__4332 (
            .O(N__26114),
            .I(N__26108));
    LocalMux I__4331 (
            .O(N__26111),
            .I(N__26105));
    LocalMux I__4330 (
            .O(N__26108),
            .I(N__26102));
    Span12Mux_v I__4329 (
            .O(N__26105),
            .I(N__26099));
    Span4Mux_h I__4328 (
            .O(N__26102),
            .I(N__26096));
    Odrv12 I__4327 (
            .O(N__26099),
            .I(\pid_alt.error_p_reg_esr_RNIFTRL5Z0Z_3 ));
    Odrv4 I__4326 (
            .O(N__26096),
            .I(\pid_alt.error_p_reg_esr_RNIFTRL5Z0Z_3 ));
    CascadeMux I__4325 (
            .O(N__26091),
            .I(N__26088));
    InMux I__4324 (
            .O(N__26088),
            .I(N__26085));
    LocalMux I__4323 (
            .O(N__26085),
            .I(N__26082));
    Span4Mux_h I__4322 (
            .O(N__26082),
            .I(N__26079));
    Odrv4 I__4321 (
            .O(N__26079),
            .I(\pid_alt.error_d_reg_prev_esr_RNIRFO19Z0Z_3 ));
    InMux I__4320 (
            .O(N__26076),
            .I(N__26070));
    InMux I__4319 (
            .O(N__26075),
            .I(N__26070));
    LocalMux I__4318 (
            .O(N__26070),
            .I(N__26067));
    Span4Mux_v I__4317 (
            .O(N__26067),
            .I(N__26064));
    Span4Mux_h I__4316 (
            .O(N__26064),
            .I(N__26061));
    Odrv4 I__4315 (
            .O(N__26061),
            .I(\pid_alt.error_d_reg_prev_esr_RNI3M511Z0Z_3 ));
    InMux I__4314 (
            .O(N__26058),
            .I(N__26052));
    InMux I__4313 (
            .O(N__26057),
            .I(N__26052));
    LocalMux I__4312 (
            .O(N__26052),
            .I(\pid_alt.error_d_reg_prev_esr_RNI6P511_0Z0Z_4 ));
    CascadeMux I__4311 (
            .O(N__26049),
            .I(N__26045));
    InMux I__4310 (
            .O(N__26048),
            .I(N__26042));
    InMux I__4309 (
            .O(N__26045),
            .I(N__26039));
    LocalMux I__4308 (
            .O(N__26042),
            .I(N__26036));
    LocalMux I__4307 (
            .O(N__26039),
            .I(N__26033));
    Span4Mux_h I__4306 (
            .O(N__26036),
            .I(N__26030));
    Span4Mux_v I__4305 (
            .O(N__26033),
            .I(N__26027));
    Odrv4 I__4304 (
            .O(N__26030),
            .I(\pid_alt.error_d_reg_prev_esr_RNICISB3Z0Z_3 ));
    Odrv4 I__4303 (
            .O(N__26027),
            .I(\pid_alt.error_d_reg_prev_esr_RNICISB3Z0Z_3 ));
    CascadeMux I__4302 (
            .O(N__26022),
            .I(N__26019));
    InMux I__4301 (
            .O(N__26019),
            .I(N__26013));
    InMux I__4300 (
            .O(N__26018),
            .I(N__26013));
    LocalMux I__4299 (
            .O(N__26013),
            .I(\pid_alt.error_d_reg_prevZ0Z_4 ));
    InMux I__4298 (
            .O(N__26010),
            .I(N__26007));
    LocalMux I__4297 (
            .O(N__26007),
            .I(N__26002));
    InMux I__4296 (
            .O(N__26006),
            .I(N__25997));
    InMux I__4295 (
            .O(N__26005),
            .I(N__25997));
    Span4Mux_v I__4294 (
            .O(N__26002),
            .I(N__25992));
    LocalMux I__4293 (
            .O(N__25997),
            .I(N__25992));
    Span4Mux_h I__4292 (
            .O(N__25992),
            .I(N__25989));
    Odrv4 I__4291 (
            .O(N__25989),
            .I(\pid_alt.pid_preregZ0Z_6 ));
    InMux I__4290 (
            .O(N__25986),
            .I(N__25982));
    InMux I__4289 (
            .O(N__25985),
            .I(N__25979));
    LocalMux I__4288 (
            .O(N__25982),
            .I(N__25976));
    LocalMux I__4287 (
            .O(N__25979),
            .I(N__25972));
    Span4Mux_h I__4286 (
            .O(N__25976),
            .I(N__25969));
    InMux I__4285 (
            .O(N__25975),
            .I(N__25966));
    Odrv4 I__4284 (
            .O(N__25972),
            .I(\pid_alt.pid_preregZ0Z_0 ));
    Odrv4 I__4283 (
            .O(N__25969),
            .I(\pid_alt.pid_preregZ0Z_0 ));
    LocalMux I__4282 (
            .O(N__25966),
            .I(\pid_alt.pid_preregZ0Z_0 ));
    InMux I__4281 (
            .O(N__25959),
            .I(N__25955));
    CascadeMux I__4280 (
            .O(N__25958),
            .I(N__25952));
    LocalMux I__4279 (
            .O(N__25955),
            .I(N__25948));
    InMux I__4278 (
            .O(N__25952),
            .I(N__25945));
    InMux I__4277 (
            .O(N__25951),
            .I(N__25942));
    Span4Mux_h I__4276 (
            .O(N__25948),
            .I(N__25937));
    LocalMux I__4275 (
            .O(N__25945),
            .I(N__25937));
    LocalMux I__4274 (
            .O(N__25942),
            .I(\pid_alt.pid_preregZ0Z_1 ));
    Odrv4 I__4273 (
            .O(N__25937),
            .I(\pid_alt.pid_preregZ0Z_1 ));
    InMux I__4272 (
            .O(N__25932),
            .I(N__25929));
    LocalMux I__4271 (
            .O(N__25929),
            .I(N__25924));
    InMux I__4270 (
            .O(N__25928),
            .I(N__25919));
    InMux I__4269 (
            .O(N__25927),
            .I(N__25919));
    Odrv4 I__4268 (
            .O(N__25924),
            .I(\pid_alt.pid_preregZ0Z_2 ));
    LocalMux I__4267 (
            .O(N__25919),
            .I(\pid_alt.pid_preregZ0Z_2 ));
    InMux I__4266 (
            .O(N__25914),
            .I(N__25911));
    LocalMux I__4265 (
            .O(N__25911),
            .I(N__25908));
    Span4Mux_v I__4264 (
            .O(N__25908),
            .I(N__25901));
    InMux I__4263 (
            .O(N__25907),
            .I(N__25892));
    InMux I__4262 (
            .O(N__25906),
            .I(N__25892));
    InMux I__4261 (
            .O(N__25905),
            .I(N__25892));
    InMux I__4260 (
            .O(N__25904),
            .I(N__25892));
    Odrv4 I__4259 (
            .O(N__25901),
            .I(\pid_alt.N_91_1 ));
    LocalMux I__4258 (
            .O(N__25892),
            .I(\pid_alt.N_91_1 ));
    InMux I__4257 (
            .O(N__25887),
            .I(N__25883));
    CascadeMux I__4256 (
            .O(N__25886),
            .I(N__25880));
    LocalMux I__4255 (
            .O(N__25883),
            .I(N__25876));
    InMux I__4254 (
            .O(N__25880),
            .I(N__25871));
    InMux I__4253 (
            .O(N__25879),
            .I(N__25871));
    Odrv12 I__4252 (
            .O(N__25876),
            .I(\pid_alt.pid_preregZ0Z_3 ));
    LocalMux I__4251 (
            .O(N__25871),
            .I(\pid_alt.pid_preregZ0Z_3 ));
    InMux I__4250 (
            .O(N__25866),
            .I(N__25863));
    LocalMux I__4249 (
            .O(N__25863),
            .I(N__25859));
    InMux I__4248 (
            .O(N__25862),
            .I(N__25856));
    Span4Mux_v I__4247 (
            .O(N__25859),
            .I(N__25853));
    LocalMux I__4246 (
            .O(N__25856),
            .I(\Commands_frame_decoder.state_ns_i_a2_1_1Z0Z_0 ));
    Odrv4 I__4245 (
            .O(N__25853),
            .I(\Commands_frame_decoder.state_ns_i_a2_1_1Z0Z_0 ));
    InMux I__4244 (
            .O(N__25848),
            .I(N__25844));
    InMux I__4243 (
            .O(N__25847),
            .I(N__25841));
    LocalMux I__4242 (
            .O(N__25844),
            .I(N__25836));
    LocalMux I__4241 (
            .O(N__25841),
            .I(N__25836));
    Span4Mux_h I__4240 (
            .O(N__25836),
            .I(N__25833));
    Span4Mux_v I__4239 (
            .O(N__25833),
            .I(N__25830));
    Span4Mux_v I__4238 (
            .O(N__25830),
            .I(N__25827));
    Odrv4 I__4237 (
            .O(N__25827),
            .I(\pid_alt.error_p_regZ0Z_5 ));
    InMux I__4236 (
            .O(N__25824),
            .I(N__25820));
    InMux I__4235 (
            .O(N__25823),
            .I(N__25817));
    LocalMux I__4234 (
            .O(N__25820),
            .I(N__25812));
    LocalMux I__4233 (
            .O(N__25817),
            .I(N__25812));
    Odrv4 I__4232 (
            .O(N__25812),
            .I(\pid_alt.error_d_reg_prevZ0Z_5 ));
    InMux I__4231 (
            .O(N__25809),
            .I(N__25803));
    InMux I__4230 (
            .O(N__25808),
            .I(N__25803));
    LocalMux I__4229 (
            .O(N__25803),
            .I(N__25799));
    InMux I__4228 (
            .O(N__25802),
            .I(N__25796));
    Span4Mux_v I__4227 (
            .O(N__25799),
            .I(N__25793));
    LocalMux I__4226 (
            .O(N__25796),
            .I(N__25790));
    Sp12to4 I__4225 (
            .O(N__25793),
            .I(N__25785));
    Span12Mux_v I__4224 (
            .O(N__25790),
            .I(N__25785));
    Odrv12 I__4223 (
            .O(N__25785),
            .I(\pid_alt.error_d_regZ0Z_5 ));
    InMux I__4222 (
            .O(N__25782),
            .I(N__25776));
    InMux I__4221 (
            .O(N__25781),
            .I(N__25776));
    LocalMux I__4220 (
            .O(N__25776),
            .I(N__25773));
    Odrv4 I__4219 (
            .O(N__25773),
            .I(\pid_alt.error_d_reg_prev_esr_RNI9S511Z0Z_5 ));
    CascadeMux I__4218 (
            .O(N__25770),
            .I(N__25766));
    InMux I__4217 (
            .O(N__25769),
            .I(N__25763));
    InMux I__4216 (
            .O(N__25766),
            .I(N__25760));
    LocalMux I__4215 (
            .O(N__25763),
            .I(\uart_drone.data_AuxZ0Z_6 ));
    LocalMux I__4214 (
            .O(N__25760),
            .I(\uart_drone.data_AuxZ0Z_6 ));
    CascadeMux I__4213 (
            .O(N__25755),
            .I(N__25751));
    InMux I__4212 (
            .O(N__25754),
            .I(N__25748));
    InMux I__4211 (
            .O(N__25751),
            .I(N__25745));
    LocalMux I__4210 (
            .O(N__25748),
            .I(\uart_drone.data_AuxZ0Z_7 ));
    LocalMux I__4209 (
            .O(N__25745),
            .I(\uart_drone.data_AuxZ0Z_7 ));
    CEMux I__4208 (
            .O(N__25740),
            .I(N__25737));
    LocalMux I__4207 (
            .O(N__25737),
            .I(N__25734));
    Odrv4 I__4206 (
            .O(N__25734),
            .I(\Commands_frame_decoder.source_CH3data_1_sqmuxa_0 ));
    CascadeMux I__4205 (
            .O(N__25731),
            .I(\Commands_frame_decoder.source_CH3data_1_sqmuxa_cascade_ ));
    InMux I__4204 (
            .O(N__25728),
            .I(N__25724));
    InMux I__4203 (
            .O(N__25727),
            .I(N__25721));
    LocalMux I__4202 (
            .O(N__25724),
            .I(\Commands_frame_decoder.stateZ0Z_5 ));
    LocalMux I__4201 (
            .O(N__25721),
            .I(\Commands_frame_decoder.stateZ0Z_5 ));
    InMux I__4200 (
            .O(N__25716),
            .I(N__25713));
    LocalMux I__4199 (
            .O(N__25713),
            .I(N__25710));
    Odrv4 I__4198 (
            .O(N__25710),
            .I(\Commands_frame_decoder.source_CH4data_1_sqmuxa ));
    CascadeMux I__4197 (
            .O(N__25707),
            .I(\Commands_frame_decoder.source_CH4data_1_sqmuxa_cascade_ ));
    CascadeMux I__4196 (
            .O(N__25704),
            .I(N__25700));
    InMux I__4195 (
            .O(N__25703),
            .I(N__25697));
    InMux I__4194 (
            .O(N__25700),
            .I(N__25694));
    LocalMux I__4193 (
            .O(N__25697),
            .I(\uart_drone.data_AuxZ0Z_0 ));
    LocalMux I__4192 (
            .O(N__25694),
            .I(\uart_drone.data_AuxZ0Z_0 ));
    CascadeMux I__4191 (
            .O(N__25689),
            .I(N__25685));
    InMux I__4190 (
            .O(N__25688),
            .I(N__25682));
    InMux I__4189 (
            .O(N__25685),
            .I(N__25679));
    LocalMux I__4188 (
            .O(N__25682),
            .I(\uart_drone.data_AuxZ0Z_1 ));
    LocalMux I__4187 (
            .O(N__25679),
            .I(\uart_drone.data_AuxZ0Z_1 ));
    CascadeMux I__4186 (
            .O(N__25674),
            .I(N__25670));
    InMux I__4185 (
            .O(N__25673),
            .I(N__25667));
    InMux I__4184 (
            .O(N__25670),
            .I(N__25664));
    LocalMux I__4183 (
            .O(N__25667),
            .I(\uart_drone.data_AuxZ0Z_2 ));
    LocalMux I__4182 (
            .O(N__25664),
            .I(\uart_drone.data_AuxZ0Z_2 ));
    CascadeMux I__4181 (
            .O(N__25659),
            .I(N__25655));
    InMux I__4180 (
            .O(N__25658),
            .I(N__25652));
    InMux I__4179 (
            .O(N__25655),
            .I(N__25649));
    LocalMux I__4178 (
            .O(N__25652),
            .I(\uart_drone.data_AuxZ0Z_3 ));
    LocalMux I__4177 (
            .O(N__25649),
            .I(\uart_drone.data_AuxZ0Z_3 ));
    InMux I__4176 (
            .O(N__25644),
            .I(N__25640));
    InMux I__4175 (
            .O(N__25643),
            .I(N__25637));
    LocalMux I__4174 (
            .O(N__25640),
            .I(\uart_drone.data_AuxZ0Z_4 ));
    LocalMux I__4173 (
            .O(N__25637),
            .I(\uart_drone.data_AuxZ0Z_4 ));
    CascadeMux I__4172 (
            .O(N__25632),
            .I(N__25628));
    InMux I__4171 (
            .O(N__25631),
            .I(N__25625));
    InMux I__4170 (
            .O(N__25628),
            .I(N__25622));
    LocalMux I__4169 (
            .O(N__25625),
            .I(\uart_drone.data_AuxZ0Z_5 ));
    LocalMux I__4168 (
            .O(N__25622),
            .I(\uart_drone.data_AuxZ0Z_5 ));
    InMux I__4167 (
            .O(N__25617),
            .I(N__25612));
    InMux I__4166 (
            .O(N__25616),
            .I(N__25609));
    InMux I__4165 (
            .O(N__25615),
            .I(N__25606));
    LocalMux I__4164 (
            .O(N__25612),
            .I(\Commands_frame_decoder.N_320_0 ));
    LocalMux I__4163 (
            .O(N__25609),
            .I(\Commands_frame_decoder.N_320_0 ));
    LocalMux I__4162 (
            .O(N__25606),
            .I(\Commands_frame_decoder.N_320_0 ));
    InMux I__4161 (
            .O(N__25599),
            .I(N__25596));
    LocalMux I__4160 (
            .O(N__25596),
            .I(\Commands_frame_decoder.state_ns_i_a2_2_1Z0Z_0 ));
    CascadeMux I__4159 (
            .O(N__25593),
            .I(\Commands_frame_decoder.state_ns_0_a4_0_0_2_cascade_ ));
    InMux I__4158 (
            .O(N__25590),
            .I(N__25587));
    LocalMux I__4157 (
            .O(N__25587),
            .I(\Commands_frame_decoder.state_ns_0_a4_0_3_2 ));
    InMux I__4156 (
            .O(N__25584),
            .I(N__25578));
    InMux I__4155 (
            .O(N__25583),
            .I(N__25573));
    InMux I__4154 (
            .O(N__25582),
            .I(N__25573));
    InMux I__4153 (
            .O(N__25581),
            .I(N__25570));
    LocalMux I__4152 (
            .O(N__25578),
            .I(\Commands_frame_decoder.stateZ0Z_1 ));
    LocalMux I__4151 (
            .O(N__25573),
            .I(\Commands_frame_decoder.stateZ0Z_1 ));
    LocalMux I__4150 (
            .O(N__25570),
            .I(\Commands_frame_decoder.stateZ0Z_1 ));
    InMux I__4149 (
            .O(N__25563),
            .I(N__25556));
    InMux I__4148 (
            .O(N__25562),
            .I(N__25556));
    InMux I__4147 (
            .O(N__25561),
            .I(N__25553));
    LocalMux I__4146 (
            .O(N__25556),
            .I(\Commands_frame_decoder.N_364 ));
    LocalMux I__4145 (
            .O(N__25553),
            .I(\Commands_frame_decoder.N_364 ));
    CascadeMux I__4144 (
            .O(N__25548),
            .I(\Commands_frame_decoder.N_360_cascade_ ));
    InMux I__4143 (
            .O(N__25545),
            .I(N__25542));
    LocalMux I__4142 (
            .O(N__25542),
            .I(\Commands_frame_decoder.N_359 ));
    CascadeMux I__4141 (
            .O(N__25539),
            .I(N__25536));
    InMux I__4140 (
            .O(N__25536),
            .I(N__25533));
    LocalMux I__4139 (
            .O(N__25533),
            .I(\Commands_frame_decoder.state_ns_i_0_0 ));
    CascadeMux I__4138 (
            .O(N__25530),
            .I(N__25525));
    InMux I__4137 (
            .O(N__25529),
            .I(N__25519));
    InMux I__4136 (
            .O(N__25528),
            .I(N__25519));
    InMux I__4135 (
            .O(N__25525),
            .I(N__25516));
    InMux I__4134 (
            .O(N__25524),
            .I(N__25513));
    LocalMux I__4133 (
            .O(N__25519),
            .I(\Commands_frame_decoder.stateZ0Z_6 ));
    LocalMux I__4132 (
            .O(N__25516),
            .I(\Commands_frame_decoder.stateZ0Z_6 ));
    LocalMux I__4131 (
            .O(N__25513),
            .I(\Commands_frame_decoder.stateZ0Z_6 ));
    InMux I__4130 (
            .O(N__25506),
            .I(N__25503));
    LocalMux I__4129 (
            .O(N__25503),
            .I(N__25500));
    Span4Mux_v I__4128 (
            .O(N__25500),
            .I(N__25497));
    Span4Mux_v I__4127 (
            .O(N__25497),
            .I(N__25494));
    Sp12to4 I__4126 (
            .O(N__25494),
            .I(N__25490));
    InMux I__4125 (
            .O(N__25493),
            .I(N__25487));
    Span12Mux_s10_h I__4124 (
            .O(N__25490),
            .I(N__25484));
    LocalMux I__4123 (
            .O(N__25487),
            .I(alt_kp_4));
    Odrv12 I__4122 (
            .O(N__25484),
            .I(alt_kp_4));
    InMux I__4121 (
            .O(N__25479),
            .I(N__25475));
    InMux I__4120 (
            .O(N__25478),
            .I(N__25472));
    LocalMux I__4119 (
            .O(N__25475),
            .I(\Commands_frame_decoder.stateZ0Z_4 ));
    LocalMux I__4118 (
            .O(N__25472),
            .I(\Commands_frame_decoder.stateZ0Z_4 ));
    InMux I__4117 (
            .O(N__25467),
            .I(N__25464));
    LocalMux I__4116 (
            .O(N__25464),
            .I(\Commands_frame_decoder.source_CH3data_1_sqmuxa ));
    InMux I__4115 (
            .O(N__25461),
            .I(N__25458));
    LocalMux I__4114 (
            .O(N__25458),
            .I(\uart_pc_sync.aux_2__0_Z0Z_0 ));
    InMux I__4113 (
            .O(N__25455),
            .I(N__25452));
    LocalMux I__4112 (
            .O(N__25452),
            .I(N__25449));
    Odrv4 I__4111 (
            .O(N__25449),
            .I(\uart_pc_sync.aux_0__0_Z0Z_0 ));
    InMux I__4110 (
            .O(N__25446),
            .I(N__25443));
    LocalMux I__4109 (
            .O(N__25443),
            .I(\uart_pc_sync.aux_1__0_Z0Z_0 ));
    SRMux I__4108 (
            .O(N__25440),
            .I(N__25436));
    SRMux I__4107 (
            .O(N__25439),
            .I(N__25433));
    LocalMux I__4106 (
            .O(N__25436),
            .I(\Commands_frame_decoder.un1_state53_iZ0 ));
    LocalMux I__4105 (
            .O(N__25433),
            .I(\Commands_frame_decoder.un1_state53_iZ0 ));
    InMux I__4104 (
            .O(N__25428),
            .I(N__25422));
    InMux I__4103 (
            .O(N__25427),
            .I(N__25417));
    InMux I__4102 (
            .O(N__25426),
            .I(N__25417));
    InMux I__4101 (
            .O(N__25425),
            .I(N__25414));
    LocalMux I__4100 (
            .O(N__25422),
            .I(\Commands_frame_decoder.WDTZ0Z_13 ));
    LocalMux I__4099 (
            .O(N__25417),
            .I(\Commands_frame_decoder.WDTZ0Z_13 ));
    LocalMux I__4098 (
            .O(N__25414),
            .I(\Commands_frame_decoder.WDTZ0Z_13 ));
    InMux I__4097 (
            .O(N__25407),
            .I(N__25401));
    InMux I__4096 (
            .O(N__25406),
            .I(N__25398));
    InMux I__4095 (
            .O(N__25405),
            .I(N__25395));
    InMux I__4094 (
            .O(N__25404),
            .I(N__25392));
    LocalMux I__4093 (
            .O(N__25401),
            .I(\Commands_frame_decoder.WDTZ0Z_12 ));
    LocalMux I__4092 (
            .O(N__25398),
            .I(\Commands_frame_decoder.WDTZ0Z_12 ));
    LocalMux I__4091 (
            .O(N__25395),
            .I(\Commands_frame_decoder.WDTZ0Z_12 ));
    LocalMux I__4090 (
            .O(N__25392),
            .I(\Commands_frame_decoder.WDTZ0Z_12 ));
    InMux I__4089 (
            .O(N__25383),
            .I(N__25377));
    InMux I__4088 (
            .O(N__25382),
            .I(N__25374));
    InMux I__4087 (
            .O(N__25381),
            .I(N__25371));
    InMux I__4086 (
            .O(N__25380),
            .I(N__25368));
    LocalMux I__4085 (
            .O(N__25377),
            .I(\Commands_frame_decoder.WDTZ0Z_11 ));
    LocalMux I__4084 (
            .O(N__25374),
            .I(\Commands_frame_decoder.WDTZ0Z_11 ));
    LocalMux I__4083 (
            .O(N__25371),
            .I(\Commands_frame_decoder.WDTZ0Z_11 ));
    LocalMux I__4082 (
            .O(N__25368),
            .I(\Commands_frame_decoder.WDTZ0Z_11 ));
    InMux I__4081 (
            .O(N__25359),
            .I(N__25355));
    InMux I__4080 (
            .O(N__25358),
            .I(N__25351));
    LocalMux I__4079 (
            .O(N__25355),
            .I(N__25348));
    InMux I__4078 (
            .O(N__25354),
            .I(N__25343));
    LocalMux I__4077 (
            .O(N__25351),
            .I(N__25340));
    Span4Mux_h I__4076 (
            .O(N__25348),
            .I(N__25337));
    InMux I__4075 (
            .O(N__25347),
            .I(N__25334));
    InMux I__4074 (
            .O(N__25346),
            .I(N__25331));
    LocalMux I__4073 (
            .O(N__25343),
            .I(\Commands_frame_decoder.WDTZ0Z_15 ));
    Odrv4 I__4072 (
            .O(N__25340),
            .I(\Commands_frame_decoder.WDTZ0Z_15 ));
    Odrv4 I__4071 (
            .O(N__25337),
            .I(\Commands_frame_decoder.WDTZ0Z_15 ));
    LocalMux I__4070 (
            .O(N__25334),
            .I(\Commands_frame_decoder.WDTZ0Z_15 ));
    LocalMux I__4069 (
            .O(N__25331),
            .I(\Commands_frame_decoder.WDTZ0Z_15 ));
    CascadeMux I__4068 (
            .O(N__25320),
            .I(\Commands_frame_decoder.state_0_sqmuxacf0_1_cascade_ ));
    InMux I__4067 (
            .O(N__25317),
            .I(N__25312));
    InMux I__4066 (
            .O(N__25316),
            .I(N__25309));
    InMux I__4065 (
            .O(N__25315),
            .I(N__25304));
    LocalMux I__4064 (
            .O(N__25312),
            .I(N__25299));
    LocalMux I__4063 (
            .O(N__25309),
            .I(N__25299));
    InMux I__4062 (
            .O(N__25308),
            .I(N__25296));
    InMux I__4061 (
            .O(N__25307),
            .I(N__25293));
    LocalMux I__4060 (
            .O(N__25304),
            .I(\Commands_frame_decoder.WDTZ0Z_14 ));
    Odrv4 I__4059 (
            .O(N__25299),
            .I(\Commands_frame_decoder.WDTZ0Z_14 ));
    LocalMux I__4058 (
            .O(N__25296),
            .I(\Commands_frame_decoder.WDTZ0Z_14 ));
    LocalMux I__4057 (
            .O(N__25293),
            .I(\Commands_frame_decoder.WDTZ0Z_14 ));
    InMux I__4056 (
            .O(N__25284),
            .I(N__25281));
    LocalMux I__4055 (
            .O(N__25281),
            .I(N__25278));
    Odrv4 I__4054 (
            .O(N__25278),
            .I(\Commands_frame_decoder.state_0_sqmuxacf0 ));
    CascadeMux I__4053 (
            .O(N__25275),
            .I(N__25272));
    InMux I__4052 (
            .O(N__25272),
            .I(N__25269));
    LocalMux I__4051 (
            .O(N__25269),
            .I(N__25263));
    InMux I__4050 (
            .O(N__25268),
            .I(N__25256));
    InMux I__4049 (
            .O(N__25267),
            .I(N__25256));
    InMux I__4048 (
            .O(N__25266),
            .I(N__25256));
    Odrv12 I__4047 (
            .O(N__25263),
            .I(\Commands_frame_decoder.preinitZ0 ));
    LocalMux I__4046 (
            .O(N__25256),
            .I(\Commands_frame_decoder.preinitZ0 ));
    InMux I__4045 (
            .O(N__25251),
            .I(N__25248));
    LocalMux I__4044 (
            .O(N__25248),
            .I(N__25245));
    Odrv4 I__4043 (
            .O(N__25245),
            .I(\Commands_frame_decoder.count_1_sqmuxa ));
    InMux I__4042 (
            .O(N__25242),
            .I(N__25239));
    LocalMux I__4041 (
            .O(N__25239),
            .I(N__25235));
    InMux I__4040 (
            .O(N__25238),
            .I(N__25232));
    Odrv4 I__4039 (
            .O(N__25235),
            .I(\Commands_frame_decoder.stateZ0Z_0 ));
    LocalMux I__4038 (
            .O(N__25232),
            .I(\Commands_frame_decoder.stateZ0Z_0 ));
    CascadeMux I__4037 (
            .O(N__25227),
            .I(N__25224));
    InMux I__4036 (
            .O(N__25224),
            .I(N__25221));
    LocalMux I__4035 (
            .O(N__25221),
            .I(\Commands_frame_decoder.state_ns_0_a4_0_1_1 ));
    InMux I__4034 (
            .O(N__25218),
            .I(N__25213));
    InMux I__4033 (
            .O(N__25217),
            .I(N__25210));
    InMux I__4032 (
            .O(N__25216),
            .I(N__25206));
    LocalMux I__4031 (
            .O(N__25213),
            .I(N__25201));
    LocalMux I__4030 (
            .O(N__25210),
            .I(N__25201));
    InMux I__4029 (
            .O(N__25209),
            .I(N__25198));
    LocalMux I__4028 (
            .O(N__25206),
            .I(N__25195));
    Span12Mux_v I__4027 (
            .O(N__25201),
            .I(N__25192));
    LocalMux I__4026 (
            .O(N__25198),
            .I(N__25187));
    Span4Mux_v I__4025 (
            .O(N__25195),
            .I(N__25187));
    Odrv12 I__4024 (
            .O(N__25192),
            .I(uart_drone_data_4));
    Odrv4 I__4023 (
            .O(N__25187),
            .I(uart_drone_data_4));
    InMux I__4022 (
            .O(N__25182),
            .I(N__25179));
    LocalMux I__4021 (
            .O(N__25179),
            .I(drone_altitude_12));
    InMux I__4020 (
            .O(N__25176),
            .I(N__25171));
    InMux I__4019 (
            .O(N__25175),
            .I(N__25168));
    InMux I__4018 (
            .O(N__25174),
            .I(N__25165));
    LocalMux I__4017 (
            .O(N__25171),
            .I(N__25160));
    LocalMux I__4016 (
            .O(N__25168),
            .I(N__25160));
    LocalMux I__4015 (
            .O(N__25165),
            .I(N__25157));
    Span12Mux_v I__4014 (
            .O(N__25160),
            .I(N__25154));
    Span4Mux_v I__4013 (
            .O(N__25157),
            .I(N__25151));
    Odrv12 I__4012 (
            .O(N__25154),
            .I(uart_drone_data_5));
    Odrv4 I__4011 (
            .O(N__25151),
            .I(uart_drone_data_5));
    InMux I__4010 (
            .O(N__25146),
            .I(N__25143));
    LocalMux I__4009 (
            .O(N__25143),
            .I(drone_altitude_13));
    InMux I__4008 (
            .O(N__25140),
            .I(N__25134));
    InMux I__4007 (
            .O(N__25139),
            .I(N__25131));
    InMux I__4006 (
            .O(N__25138),
            .I(N__25128));
    CascadeMux I__4005 (
            .O(N__25137),
            .I(N__25125));
    LocalMux I__4004 (
            .O(N__25134),
            .I(N__25120));
    LocalMux I__4003 (
            .O(N__25131),
            .I(N__25120));
    LocalMux I__4002 (
            .O(N__25128),
            .I(N__25117));
    InMux I__4001 (
            .O(N__25125),
            .I(N__25114));
    Span12Mux_v I__4000 (
            .O(N__25120),
            .I(N__25111));
    Span4Mux_h I__3999 (
            .O(N__25117),
            .I(N__25108));
    LocalMux I__3998 (
            .O(N__25114),
            .I(N__25105));
    Odrv12 I__3997 (
            .O(N__25111),
            .I(uart_drone_data_6));
    Odrv4 I__3996 (
            .O(N__25108),
            .I(uart_drone_data_6));
    Odrv4 I__3995 (
            .O(N__25105),
            .I(uart_drone_data_6));
    InMux I__3994 (
            .O(N__25098),
            .I(N__25095));
    LocalMux I__3993 (
            .O(N__25095),
            .I(drone_altitude_14));
    InMux I__3992 (
            .O(N__25092),
            .I(N__25087));
    InMux I__3991 (
            .O(N__25091),
            .I(N__25084));
    InMux I__3990 (
            .O(N__25090),
            .I(N__25081));
    LocalMux I__3989 (
            .O(N__25087),
            .I(N__25076));
    LocalMux I__3988 (
            .O(N__25084),
            .I(N__25076));
    LocalMux I__3987 (
            .O(N__25081),
            .I(N__25073));
    Span12Mux_v I__3986 (
            .O(N__25076),
            .I(N__25070));
    Span4Mux_h I__3985 (
            .O(N__25073),
            .I(N__25067));
    Odrv12 I__3984 (
            .O(N__25070),
            .I(uart_drone_data_7));
    Odrv4 I__3983 (
            .O(N__25067),
            .I(uart_drone_data_7));
    InMux I__3982 (
            .O(N__25062),
            .I(N__25059));
    LocalMux I__3981 (
            .O(N__25059),
            .I(N__25056));
    Odrv4 I__3980 (
            .O(N__25056),
            .I(drone_altitude_15));
    InMux I__3979 (
            .O(N__25053),
            .I(N__25050));
    LocalMux I__3978 (
            .O(N__25050),
            .I(N__25046));
    InMux I__3977 (
            .O(N__25049),
            .I(N__25043));
    Span4Mux_v I__3976 (
            .O(N__25046),
            .I(N__25037));
    LocalMux I__3975 (
            .O(N__25043),
            .I(N__25037));
    InMux I__3974 (
            .O(N__25042),
            .I(N__25034));
    Span4Mux_v I__3973 (
            .O(N__25037),
            .I(N__25031));
    LocalMux I__3972 (
            .O(N__25034),
            .I(N__25028));
    Span4Mux_v I__3971 (
            .O(N__25031),
            .I(N__25023));
    Span4Mux_h I__3970 (
            .O(N__25028),
            .I(N__25023));
    Odrv4 I__3969 (
            .O(N__25023),
            .I(uart_drone_data_0));
    CascadeMux I__3968 (
            .O(N__25020),
            .I(N__25017));
    InMux I__3967 (
            .O(N__25017),
            .I(N__25014));
    LocalMux I__3966 (
            .O(N__25014),
            .I(\dron_frame_decoder_1.drone_altitude_8 ));
    InMux I__3965 (
            .O(N__25011),
            .I(N__25006));
    InMux I__3964 (
            .O(N__25010),
            .I(N__25003));
    InMux I__3963 (
            .O(N__25009),
            .I(N__24999));
    LocalMux I__3962 (
            .O(N__25006),
            .I(N__24994));
    LocalMux I__3961 (
            .O(N__25003),
            .I(N__24994));
    InMux I__3960 (
            .O(N__25002),
            .I(N__24991));
    LocalMux I__3959 (
            .O(N__24999),
            .I(N__24988));
    Span12Mux_v I__3958 (
            .O(N__24994),
            .I(N__24985));
    LocalMux I__3957 (
            .O(N__24991),
            .I(N__24982));
    Span4Mux_h I__3956 (
            .O(N__24988),
            .I(N__24979));
    Odrv12 I__3955 (
            .O(N__24985),
            .I(uart_drone_data_1));
    Odrv4 I__3954 (
            .O(N__24982),
            .I(uart_drone_data_1));
    Odrv4 I__3953 (
            .O(N__24979),
            .I(uart_drone_data_1));
    InMux I__3952 (
            .O(N__24972),
            .I(N__24969));
    LocalMux I__3951 (
            .O(N__24969),
            .I(\dron_frame_decoder_1.drone_altitude_9 ));
    InMux I__3950 (
            .O(N__24966),
            .I(N__24963));
    LocalMux I__3949 (
            .O(N__24963),
            .I(N__24958));
    CascadeMux I__3948 (
            .O(N__24962),
            .I(N__24954));
    InMux I__3947 (
            .O(N__24961),
            .I(N__24951));
    Span4Mux_s3_v I__3946 (
            .O(N__24958),
            .I(N__24947));
    InMux I__3945 (
            .O(N__24957),
            .I(N__24942));
    InMux I__3944 (
            .O(N__24954),
            .I(N__24942));
    LocalMux I__3943 (
            .O(N__24951),
            .I(N__24939));
    InMux I__3942 (
            .O(N__24950),
            .I(N__24936));
    Span4Mux_v I__3941 (
            .O(N__24947),
            .I(N__24933));
    LocalMux I__3940 (
            .O(N__24942),
            .I(N__24930));
    Span4Mux_v I__3939 (
            .O(N__24939),
            .I(N__24927));
    LocalMux I__3938 (
            .O(N__24936),
            .I(N__24922));
    Span4Mux_v I__3937 (
            .O(N__24933),
            .I(N__24922));
    Span4Mux_h I__3936 (
            .O(N__24930),
            .I(N__24919));
    Odrv4 I__3935 (
            .O(N__24927),
            .I(\pid_alt.stateZ0Z_0 ));
    Odrv4 I__3934 (
            .O(N__24922),
            .I(\pid_alt.stateZ0Z_0 ));
    Odrv4 I__3933 (
            .O(N__24919),
            .I(\pid_alt.stateZ0Z_0 ));
    IoInMux I__3932 (
            .O(N__24912),
            .I(N__24909));
    LocalMux I__3931 (
            .O(N__24909),
            .I(N__24906));
    Span4Mux_s2_v I__3930 (
            .O(N__24906),
            .I(N__24903));
    Odrv4 I__3929 (
            .O(N__24903),
            .I(\pid_alt.state_0_0 ));
    CEMux I__3928 (
            .O(N__24900),
            .I(N__24897));
    LocalMux I__3927 (
            .O(N__24897),
            .I(N__24894));
    Span12Mux_h I__3926 (
            .O(N__24894),
            .I(N__24891));
    Odrv12 I__3925 (
            .O(N__24891),
            .I(\dron_frame_decoder_1.N_392_0 ));
    InMux I__3924 (
            .O(N__24888),
            .I(N__24885));
    LocalMux I__3923 (
            .O(N__24885),
            .I(N__24882));
    Span4Mux_v I__3922 (
            .O(N__24882),
            .I(N__24878));
    InMux I__3921 (
            .O(N__24881),
            .I(N__24875));
    Span4Mux_v I__3920 (
            .O(N__24878),
            .I(N__24870));
    LocalMux I__3919 (
            .O(N__24875),
            .I(N__24870));
    Odrv4 I__3918 (
            .O(N__24870),
            .I(\Commands_frame_decoder.source_offset3data_1_sqmuxa ));
    InMux I__3917 (
            .O(N__24867),
            .I(N__24864));
    LocalMux I__3916 (
            .O(N__24864),
            .I(N__24850));
    InMux I__3915 (
            .O(N__24863),
            .I(N__24845));
    InMux I__3914 (
            .O(N__24862),
            .I(N__24845));
    InMux I__3913 (
            .O(N__24861),
            .I(N__24838));
    InMux I__3912 (
            .O(N__24860),
            .I(N__24838));
    InMux I__3911 (
            .O(N__24859),
            .I(N__24838));
    InMux I__3910 (
            .O(N__24858),
            .I(N__24825));
    InMux I__3909 (
            .O(N__24857),
            .I(N__24825));
    InMux I__3908 (
            .O(N__24856),
            .I(N__24825));
    InMux I__3907 (
            .O(N__24855),
            .I(N__24825));
    InMux I__3906 (
            .O(N__24854),
            .I(N__24825));
    InMux I__3905 (
            .O(N__24853),
            .I(N__24825));
    Odrv12 I__3904 (
            .O(N__24850),
            .I(\Commands_frame_decoder.N_358 ));
    LocalMux I__3903 (
            .O(N__24845),
            .I(\Commands_frame_decoder.N_358 ));
    LocalMux I__3902 (
            .O(N__24838),
            .I(\Commands_frame_decoder.N_358 ));
    LocalMux I__3901 (
            .O(N__24825),
            .I(\Commands_frame_decoder.N_358 ));
    InMux I__3900 (
            .O(N__24816),
            .I(N__24813));
    LocalMux I__3899 (
            .O(N__24813),
            .I(\dron_frame_decoder_1.drone_altitude_4 ));
    CascadeMux I__3898 (
            .O(N__24810),
            .I(N__24807));
    InMux I__3897 (
            .O(N__24807),
            .I(N__24804));
    LocalMux I__3896 (
            .O(N__24804),
            .I(N__24801));
    Odrv4 I__3895 (
            .O(N__24801),
            .I(drone_altitude_i_4));
    InMux I__3894 (
            .O(N__24798),
            .I(N__24795));
    LocalMux I__3893 (
            .O(N__24795),
            .I(\dron_frame_decoder_1.drone_altitude_5 ));
    CascadeMux I__3892 (
            .O(N__24792),
            .I(N__24789));
    InMux I__3891 (
            .O(N__24789),
            .I(N__24786));
    LocalMux I__3890 (
            .O(N__24786),
            .I(N__24783));
    Odrv4 I__3889 (
            .O(N__24783),
            .I(drone_altitude_i_5));
    InMux I__3888 (
            .O(N__24780),
            .I(N__24777));
    LocalMux I__3887 (
            .O(N__24777),
            .I(\dron_frame_decoder_1.drone_altitude_6 ));
    InMux I__3886 (
            .O(N__24774),
            .I(N__24771));
    LocalMux I__3885 (
            .O(N__24771),
            .I(N__24768));
    Odrv4 I__3884 (
            .O(N__24768),
            .I(drone_altitude_i_6));
    InMux I__3883 (
            .O(N__24765),
            .I(N__24762));
    LocalMux I__3882 (
            .O(N__24762),
            .I(\dron_frame_decoder_1.drone_altitude_7 ));
    CascadeMux I__3881 (
            .O(N__24759),
            .I(N__24756));
    InMux I__3880 (
            .O(N__24756),
            .I(N__24753));
    LocalMux I__3879 (
            .O(N__24753),
            .I(N__24750));
    Odrv4 I__3878 (
            .O(N__24750),
            .I(drone_altitude_i_7));
    CascadeMux I__3877 (
            .O(N__24747),
            .I(N__24744));
    InMux I__3876 (
            .O(N__24744),
            .I(N__24741));
    LocalMux I__3875 (
            .O(N__24741),
            .I(N__24738));
    Span4Mux_h I__3874 (
            .O(N__24738),
            .I(N__24735));
    Odrv4 I__3873 (
            .O(N__24735),
            .I(drone_altitude_i_8));
    InMux I__3872 (
            .O(N__24732),
            .I(N__24727));
    InMux I__3871 (
            .O(N__24731),
            .I(N__24724));
    InMux I__3870 (
            .O(N__24730),
            .I(N__24721));
    LocalMux I__3869 (
            .O(N__24727),
            .I(N__24718));
    LocalMux I__3868 (
            .O(N__24724),
            .I(N__24713));
    LocalMux I__3867 (
            .O(N__24721),
            .I(N__24713));
    Span4Mux_h I__3866 (
            .O(N__24718),
            .I(N__24710));
    Odrv12 I__3865 (
            .O(N__24713),
            .I(uart_drone_data_2));
    Odrv4 I__3864 (
            .O(N__24710),
            .I(uart_drone_data_2));
    InMux I__3863 (
            .O(N__24705),
            .I(N__24702));
    LocalMux I__3862 (
            .O(N__24702),
            .I(\dron_frame_decoder_1.drone_altitude_10 ));
    InMux I__3861 (
            .O(N__24699),
            .I(N__24693));
    InMux I__3860 (
            .O(N__24698),
            .I(N__24693));
    LocalMux I__3859 (
            .O(N__24693),
            .I(\pid_alt.error_d_reg_prevZ0Z_24 ));
    InMux I__3858 (
            .O(N__24690),
            .I(N__24681));
    InMux I__3857 (
            .O(N__24689),
            .I(N__24681));
    InMux I__3856 (
            .O(N__24688),
            .I(N__24681));
    LocalMux I__3855 (
            .O(N__24681),
            .I(N__24678));
    Span4Mux_v I__3854 (
            .O(N__24678),
            .I(N__24675));
    Span4Mux_h I__3853 (
            .O(N__24675),
            .I(N__24672));
    Span4Mux_h I__3852 (
            .O(N__24672),
            .I(N__24669));
    Span4Mux_v I__3851 (
            .O(N__24669),
            .I(N__24666));
    Odrv4 I__3850 (
            .O(N__24666),
            .I(\pid_alt.error_d_regZ0Z_24 ));
    InMux I__3849 (
            .O(N__24663),
            .I(N__24654));
    InMux I__3848 (
            .O(N__24662),
            .I(N__24651));
    InMux I__3847 (
            .O(N__24661),
            .I(N__24648));
    InMux I__3846 (
            .O(N__24660),
            .I(N__24643));
    InMux I__3845 (
            .O(N__24659),
            .I(N__24643));
    InMux I__3844 (
            .O(N__24658),
            .I(N__24638));
    InMux I__3843 (
            .O(N__24657),
            .I(N__24638));
    LocalMux I__3842 (
            .O(N__24654),
            .I(N__24623));
    LocalMux I__3841 (
            .O(N__24651),
            .I(N__24623));
    LocalMux I__3840 (
            .O(N__24648),
            .I(N__24623));
    LocalMux I__3839 (
            .O(N__24643),
            .I(N__24623));
    LocalMux I__3838 (
            .O(N__24638),
            .I(N__24623));
    InMux I__3837 (
            .O(N__24637),
            .I(N__24615));
    InMux I__3836 (
            .O(N__24636),
            .I(N__24615));
    InMux I__3835 (
            .O(N__24635),
            .I(N__24615));
    InMux I__3834 (
            .O(N__24634),
            .I(N__24609));
    Span4Mux_v I__3833 (
            .O(N__24623),
            .I(N__24605));
    InMux I__3832 (
            .O(N__24622),
            .I(N__24602));
    LocalMux I__3831 (
            .O(N__24615),
            .I(N__24599));
    InMux I__3830 (
            .O(N__24614),
            .I(N__24596));
    InMux I__3829 (
            .O(N__24613),
            .I(N__24591));
    InMux I__3828 (
            .O(N__24612),
            .I(N__24591));
    LocalMux I__3827 (
            .O(N__24609),
            .I(N__24588));
    InMux I__3826 (
            .O(N__24608),
            .I(N__24585));
    Span4Mux_h I__3825 (
            .O(N__24605),
            .I(N__24580));
    LocalMux I__3824 (
            .O(N__24602),
            .I(N__24580));
    Span4Mux_v I__3823 (
            .O(N__24599),
            .I(N__24573));
    LocalMux I__3822 (
            .O(N__24596),
            .I(N__24573));
    LocalMux I__3821 (
            .O(N__24591),
            .I(N__24573));
    Span4Mux_h I__3820 (
            .O(N__24588),
            .I(N__24568));
    LocalMux I__3819 (
            .O(N__24585),
            .I(N__24568));
    Span4Mux_h I__3818 (
            .O(N__24580),
            .I(N__24565));
    Span4Mux_h I__3817 (
            .O(N__24573),
            .I(N__24560));
    Span4Mux_v I__3816 (
            .O(N__24568),
            .I(N__24560));
    Span4Mux_v I__3815 (
            .O(N__24565),
            .I(N__24557));
    Span4Mux_v I__3814 (
            .O(N__24560),
            .I(N__24554));
    Odrv4 I__3813 (
            .O(N__24557),
            .I(\pid_alt.error_p_regZ0Z_20 ));
    Odrv4 I__3812 (
            .O(N__24554),
            .I(\pid_alt.error_p_regZ0Z_20 ));
    InMux I__3811 (
            .O(N__24549),
            .I(N__24543));
    InMux I__3810 (
            .O(N__24548),
            .I(N__24543));
    LocalMux I__3809 (
            .O(N__24543),
            .I(\pid_alt.error_d_reg_prev_esr_RNIOOKMZ0Z_24 ));
    InMux I__3808 (
            .O(N__24540),
            .I(N__24536));
    InMux I__3807 (
            .O(N__24539),
            .I(N__24533));
    LocalMux I__3806 (
            .O(N__24536),
            .I(N__24530));
    LocalMux I__3805 (
            .O(N__24533),
            .I(N__24527));
    Span4Mux_v I__3804 (
            .O(N__24530),
            .I(N__24524));
    Span4Mux_h I__3803 (
            .O(N__24527),
            .I(N__24521));
    Span4Mux_h I__3802 (
            .O(N__24524),
            .I(N__24516));
    Span4Mux_v I__3801 (
            .O(N__24521),
            .I(N__24516));
    Span4Mux_h I__3800 (
            .O(N__24516),
            .I(N__24513));
    Odrv4 I__3799 (
            .O(N__24513),
            .I(\pid_alt.error_p_regZ0Z_6 ));
    InMux I__3798 (
            .O(N__24510),
            .I(N__24506));
    InMux I__3797 (
            .O(N__24509),
            .I(N__24503));
    LocalMux I__3796 (
            .O(N__24506),
            .I(N__24500));
    LocalMux I__3795 (
            .O(N__24503),
            .I(\pid_alt.error_d_reg_prevZ0Z_6 ));
    Odrv12 I__3794 (
            .O(N__24500),
            .I(\pid_alt.error_d_reg_prevZ0Z_6 ));
    InMux I__3793 (
            .O(N__24495),
            .I(N__24491));
    InMux I__3792 (
            .O(N__24494),
            .I(N__24488));
    LocalMux I__3791 (
            .O(N__24491),
            .I(N__24482));
    LocalMux I__3790 (
            .O(N__24488),
            .I(N__24482));
    InMux I__3789 (
            .O(N__24487),
            .I(N__24479));
    Span4Mux_v I__3788 (
            .O(N__24482),
            .I(N__24474));
    LocalMux I__3787 (
            .O(N__24479),
            .I(N__24474));
    Span4Mux_h I__3786 (
            .O(N__24474),
            .I(N__24471));
    Span4Mux_h I__3785 (
            .O(N__24471),
            .I(N__24468));
    Span4Mux_v I__3784 (
            .O(N__24468),
            .I(N__24465));
    Odrv4 I__3783 (
            .O(N__24465),
            .I(\pid_alt.error_d_regZ0Z_6 ));
    InMux I__3782 (
            .O(N__24462),
            .I(N__24459));
    LocalMux I__3781 (
            .O(N__24459),
            .I(N__24455));
    InMux I__3780 (
            .O(N__24458),
            .I(N__24452));
    Span4Mux_v I__3779 (
            .O(N__24455),
            .I(N__24448));
    LocalMux I__3778 (
            .O(N__24452),
            .I(N__24445));
    InMux I__3777 (
            .O(N__24451),
            .I(N__24442));
    Span4Mux_h I__3776 (
            .O(N__24448),
            .I(N__24439));
    Span4Mux_v I__3775 (
            .O(N__24445),
            .I(N__24436));
    LocalMux I__3774 (
            .O(N__24442),
            .I(N__24433));
    Span4Mux_h I__3773 (
            .O(N__24439),
            .I(N__24430));
    Span4Mux_v I__3772 (
            .O(N__24436),
            .I(N__24425));
    Span4Mux_v I__3771 (
            .O(N__24433),
            .I(N__24425));
    Span4Mux_h I__3770 (
            .O(N__24430),
            .I(N__24422));
    Span4Mux_h I__3769 (
            .O(N__24425),
            .I(N__24419));
    Span4Mux_v I__3768 (
            .O(N__24422),
            .I(N__24415));
    Span4Mux_h I__3767 (
            .O(N__24419),
            .I(N__24412));
    InMux I__3766 (
            .O(N__24418),
            .I(N__24409));
    Odrv4 I__3765 (
            .O(N__24415),
            .I(drone_altitude_0));
    Odrv4 I__3764 (
            .O(N__24412),
            .I(drone_altitude_0));
    LocalMux I__3763 (
            .O(N__24409),
            .I(drone_altitude_0));
    InMux I__3762 (
            .O(N__24402),
            .I(N__24399));
    LocalMux I__3761 (
            .O(N__24399),
            .I(drone_altitude_1));
    InMux I__3760 (
            .O(N__24396),
            .I(N__24393));
    LocalMux I__3759 (
            .O(N__24393),
            .I(drone_altitude_2));
    InMux I__3758 (
            .O(N__24390),
            .I(N__24387));
    LocalMux I__3757 (
            .O(N__24387),
            .I(drone_altitude_3));
    CascadeMux I__3756 (
            .O(N__24384),
            .I(N__24381));
    InMux I__3755 (
            .O(N__24381),
            .I(N__24378));
    LocalMux I__3754 (
            .O(N__24378),
            .I(N__24375));
    Span4Mux_h I__3753 (
            .O(N__24375),
            .I(N__24372));
    Odrv4 I__3752 (
            .O(N__24372),
            .I(\pid_alt.error_d_reg_prev_esr_RNI0BT34Z0Z_25 ));
    InMux I__3751 (
            .O(N__24369),
            .I(N__24363));
    InMux I__3750 (
            .O(N__24368),
            .I(N__24363));
    LocalMux I__3749 (
            .O(N__24363),
            .I(\pid_alt.error_d_reg_prev_esr_RNISSKM_0Z0Z_26 ));
    InMux I__3748 (
            .O(N__24360),
            .I(N__24354));
    InMux I__3747 (
            .O(N__24359),
            .I(N__24354));
    LocalMux I__3746 (
            .O(N__24354),
            .I(\pid_alt.error_d_reg_prev_esr_RNIQQKMZ0Z_25 ));
    CascadeMux I__3745 (
            .O(N__24351),
            .I(N__24348));
    InMux I__3744 (
            .O(N__24348),
            .I(N__24344));
    CascadeMux I__3743 (
            .O(N__24347),
            .I(N__24341));
    LocalMux I__3742 (
            .O(N__24344),
            .I(N__24338));
    InMux I__3741 (
            .O(N__24341),
            .I(N__24335));
    Span4Mux_v I__3740 (
            .O(N__24338),
            .I(N__24332));
    LocalMux I__3739 (
            .O(N__24335),
            .I(N__24329));
    Odrv4 I__3738 (
            .O(N__24332),
            .I(\pid_alt.error_d_reg_prev_esr_RNIINU12Z0Z_25 ));
    Odrv4 I__3737 (
            .O(N__24329),
            .I(\pid_alt.error_d_reg_prev_esr_RNIINU12Z0Z_25 ));
    CascadeMux I__3736 (
            .O(N__24324),
            .I(N__24321));
    InMux I__3735 (
            .O(N__24321),
            .I(N__24318));
    LocalMux I__3734 (
            .O(N__24318),
            .I(N__24315));
    Odrv4 I__3733 (
            .O(N__24315),
            .I(\pid_alt.error_d_reg_prev_esr_RNIO2T34Z0Z_24 ));
    InMux I__3732 (
            .O(N__24312),
            .I(N__24308));
    InMux I__3731 (
            .O(N__24311),
            .I(N__24305));
    LocalMux I__3730 (
            .O(N__24308),
            .I(\pid_alt.error_d_reg_prevZ0Z_25 ));
    LocalMux I__3729 (
            .O(N__24305),
            .I(\pid_alt.error_d_reg_prevZ0Z_25 ));
    InMux I__3728 (
            .O(N__24300),
            .I(N__24295));
    InMux I__3727 (
            .O(N__24299),
            .I(N__24290));
    InMux I__3726 (
            .O(N__24298),
            .I(N__24290));
    LocalMux I__3725 (
            .O(N__24295),
            .I(N__24285));
    LocalMux I__3724 (
            .O(N__24290),
            .I(N__24285));
    Span4Mux_v I__3723 (
            .O(N__24285),
            .I(N__24282));
    Span4Mux_h I__3722 (
            .O(N__24282),
            .I(N__24279));
    Span4Mux_h I__3721 (
            .O(N__24279),
            .I(N__24276));
    Span4Mux_v I__3720 (
            .O(N__24276),
            .I(N__24273));
    Odrv4 I__3719 (
            .O(N__24273),
            .I(\pid_alt.error_d_regZ0Z_25 ));
    InMux I__3718 (
            .O(N__24270),
            .I(N__24267));
    LocalMux I__3717 (
            .O(N__24267),
            .I(\pid_alt.error_d_reg_prev_esr_RNIQQKM_0Z0Z_25 ));
    CascadeMux I__3716 (
            .O(N__24264),
            .I(\pid_alt.error_d_reg_prev_esr_RNIQQKM_0Z0Z_25_cascade_ ));
    CascadeMux I__3715 (
            .O(N__24261),
            .I(N__24257));
    InMux I__3714 (
            .O(N__24260),
            .I(N__24254));
    InMux I__3713 (
            .O(N__24257),
            .I(N__24251));
    LocalMux I__3712 (
            .O(N__24254),
            .I(N__24248));
    LocalMux I__3711 (
            .O(N__24251),
            .I(\pid_alt.error_d_reg_prev_esr_RNIEJU12Z0Z_24 ));
    Odrv4 I__3710 (
            .O(N__24248),
            .I(\pid_alt.error_d_reg_prev_esr_RNIEJU12Z0Z_24 ));
    CascadeMux I__3709 (
            .O(N__24243),
            .I(\pid_alt.error_d_reg_prev_esr_RNIOOKM_0Z0Z_24_cascade_ ));
    CascadeMux I__3708 (
            .O(N__24240),
            .I(N__24236));
    InMux I__3707 (
            .O(N__24239),
            .I(N__24233));
    InMux I__3706 (
            .O(N__24236),
            .I(N__24230));
    LocalMux I__3705 (
            .O(N__24233),
            .I(N__24227));
    LocalMux I__3704 (
            .O(N__24230),
            .I(N__24224));
    Span4Mux_h I__3703 (
            .O(N__24227),
            .I(N__24221));
    Odrv4 I__3702 (
            .O(N__24224),
            .I(\pid_alt.error_d_reg_prev_esr_RNIAFU12Z0Z_23 ));
    Odrv4 I__3701 (
            .O(N__24221),
            .I(\pid_alt.error_d_reg_prev_esr_RNIAFU12Z0Z_23 ));
    InMux I__3700 (
            .O(N__24216),
            .I(N__24213));
    LocalMux I__3699 (
            .O(N__24213),
            .I(N__24210));
    Odrv4 I__3698 (
            .O(N__24210),
            .I(\pid_alt.un9lto29_i_a2_0_and ));
    InMux I__3697 (
            .O(N__24207),
            .I(N__24204));
    LocalMux I__3696 (
            .O(N__24204),
            .I(N__24201));
    Odrv4 I__3695 (
            .O(N__24201),
            .I(\pid_alt.N_96 ));
    CascadeMux I__3694 (
            .O(N__24198),
            .I(N__24192));
    InMux I__3693 (
            .O(N__24197),
            .I(N__24185));
    InMux I__3692 (
            .O(N__24196),
            .I(N__24185));
    InMux I__3691 (
            .O(N__24195),
            .I(N__24185));
    InMux I__3690 (
            .O(N__24192),
            .I(N__24182));
    LocalMux I__3689 (
            .O(N__24185),
            .I(N__24179));
    LocalMux I__3688 (
            .O(N__24182),
            .I(N__24176));
    Span4Mux_h I__3687 (
            .O(N__24179),
            .I(N__24173));
    Odrv12 I__3686 (
            .O(N__24176),
            .I(\pid_alt.pid_preregZ0Z_5 ));
    Odrv4 I__3685 (
            .O(N__24173),
            .I(\pid_alt.pid_preregZ0Z_5 ));
    InMux I__3684 (
            .O(N__24168),
            .I(N__24158));
    InMux I__3683 (
            .O(N__24167),
            .I(N__24158));
    InMux I__3682 (
            .O(N__24166),
            .I(N__24158));
    InMux I__3681 (
            .O(N__24165),
            .I(N__24155));
    LocalMux I__3680 (
            .O(N__24158),
            .I(N__24152));
    LocalMux I__3679 (
            .O(N__24155),
            .I(N__24147));
    Span4Mux_v I__3678 (
            .O(N__24152),
            .I(N__24147));
    Odrv4 I__3677 (
            .O(N__24147),
            .I(\pid_alt.pid_preregZ0Z_4 ));
    InMux I__3676 (
            .O(N__24144),
            .I(N__24141));
    LocalMux I__3675 (
            .O(N__24141),
            .I(N__24138));
    Odrv12 I__3674 (
            .O(N__24138),
            .I(\pid_alt.source_pid_1_sqmuxa_0_a2_0_4 ));
    InMux I__3673 (
            .O(N__24135),
            .I(N__24132));
    LocalMux I__3672 (
            .O(N__24132),
            .I(N__24129));
    Span4Mux_h I__3671 (
            .O(N__24129),
            .I(N__24125));
    InMux I__3670 (
            .O(N__24128),
            .I(N__24122));
    Span4Mux_v I__3669 (
            .O(N__24125),
            .I(N__24119));
    LocalMux I__3668 (
            .O(N__24122),
            .I(N__24116));
    Span4Mux_v I__3667 (
            .O(N__24119),
            .I(N__24113));
    Span12Mux_s9_h I__3666 (
            .O(N__24116),
            .I(N__24110));
    Span4Mux_v I__3665 (
            .O(N__24113),
            .I(N__24107));
    Odrv12 I__3664 (
            .O(N__24110),
            .I(\pid_alt.state_RNIFCSD1Z0Z_0 ));
    Odrv4 I__3663 (
            .O(N__24107),
            .I(\pid_alt.state_RNIFCSD1Z0Z_0 ));
    InMux I__3662 (
            .O(N__24102),
            .I(N__24096));
    InMux I__3661 (
            .O(N__24101),
            .I(N__24089));
    InMux I__3660 (
            .O(N__24100),
            .I(N__24089));
    InMux I__3659 (
            .O(N__24099),
            .I(N__24089));
    LocalMux I__3658 (
            .O(N__24096),
            .I(N__24086));
    LocalMux I__3657 (
            .O(N__24089),
            .I(N__24083));
    Span4Mux_v I__3656 (
            .O(N__24086),
            .I(N__24080));
    Span4Mux_v I__3655 (
            .O(N__24083),
            .I(N__24077));
    Odrv4 I__3654 (
            .O(N__24080),
            .I(\Commands_frame_decoder.source_CH1data8 ));
    Odrv4 I__3653 (
            .O(N__24077),
            .I(\Commands_frame_decoder.source_CH1data8 ));
    InMux I__3652 (
            .O(N__24072),
            .I(N__24066));
    InMux I__3651 (
            .O(N__24071),
            .I(N__24066));
    LocalMux I__3650 (
            .O(N__24066),
            .I(\pid_alt.error_d_reg_prev_esr_RNI6P511Z0Z_4 ));
    InMux I__3649 (
            .O(N__24063),
            .I(N__24057));
    InMux I__3648 (
            .O(N__24062),
            .I(N__24057));
    LocalMux I__3647 (
            .O(N__24057),
            .I(N__24054));
    Span12Mux_v I__3646 (
            .O(N__24054),
            .I(N__24051));
    Odrv12 I__3645 (
            .O(N__24051),
            .I(\pid_alt.error_p_regZ0Z_4 ));
    CascadeMux I__3644 (
            .O(N__24048),
            .I(\pid_alt.un1_reset_0_i_cascade_ ));
    InMux I__3643 (
            .O(N__24045),
            .I(N__24042));
    LocalMux I__3642 (
            .O(N__24042),
            .I(N__24039));
    Span4Mux_h I__3641 (
            .O(N__24039),
            .I(N__24036));
    Odrv4 I__3640 (
            .O(N__24036),
            .I(\pid_alt.pid_preregZ0Z_26 ));
    InMux I__3639 (
            .O(N__24033),
            .I(N__24030));
    LocalMux I__3638 (
            .O(N__24030),
            .I(N__24027));
    Span4Mux_h I__3637 (
            .O(N__24027),
            .I(N__24024));
    Odrv4 I__3636 (
            .O(N__24024),
            .I(\pid_alt.pid_preregZ0Z_25 ));
    CascadeMux I__3635 (
            .O(N__24021),
            .I(N__24018));
    InMux I__3634 (
            .O(N__24018),
            .I(N__24015));
    LocalMux I__3633 (
            .O(N__24015),
            .I(N__24012));
    Span4Mux_v I__3632 (
            .O(N__24012),
            .I(N__24009));
    Odrv4 I__3631 (
            .O(N__24009),
            .I(\pid_alt.pid_preregZ0Z_27 ));
    InMux I__3630 (
            .O(N__24006),
            .I(N__24003));
    LocalMux I__3629 (
            .O(N__24003),
            .I(N__24000));
    Span4Mux_h I__3628 (
            .O(N__24000),
            .I(N__23997));
    Odrv4 I__3627 (
            .O(N__23997),
            .I(\pid_alt.pid_preregZ0Z_24 ));
    InMux I__3626 (
            .O(N__23994),
            .I(N__23991));
    LocalMux I__3625 (
            .O(N__23991),
            .I(N__23987));
    InMux I__3624 (
            .O(N__23990),
            .I(N__23984));
    Odrv4 I__3623 (
            .O(N__23987),
            .I(\pid_alt.un9lto29_i_a2_5_and ));
    LocalMux I__3622 (
            .O(N__23984),
            .I(\pid_alt.un9lto29_i_a2_5_and ));
    InMux I__3621 (
            .O(N__23979),
            .I(N__23976));
    LocalMux I__3620 (
            .O(N__23976),
            .I(N__23969));
    InMux I__3619 (
            .O(N__23975),
            .I(N__23966));
    InMux I__3618 (
            .O(N__23974),
            .I(N__23961));
    InMux I__3617 (
            .O(N__23973),
            .I(N__23961));
    InMux I__3616 (
            .O(N__23972),
            .I(N__23958));
    Span4Mux_v I__3615 (
            .O(N__23969),
            .I(N__23953));
    LocalMux I__3614 (
            .O(N__23966),
            .I(N__23953));
    LocalMux I__3613 (
            .O(N__23961),
            .I(N__23950));
    LocalMux I__3612 (
            .O(N__23958),
            .I(\pid_alt.pid_preregZ0Z_13 ));
    Odrv4 I__3611 (
            .O(N__23953),
            .I(\pid_alt.pid_preregZ0Z_13 ));
    Odrv4 I__3610 (
            .O(N__23950),
            .I(\pid_alt.pid_preregZ0Z_13 ));
    InMux I__3609 (
            .O(N__23943),
            .I(N__23936));
    InMux I__3608 (
            .O(N__23942),
            .I(N__23936));
    InMux I__3607 (
            .O(N__23941),
            .I(N__23933));
    LocalMux I__3606 (
            .O(N__23936),
            .I(N__23930));
    LocalMux I__3605 (
            .O(N__23933),
            .I(\pid_alt.N_124 ));
    Odrv12 I__3604 (
            .O(N__23930),
            .I(\pid_alt.N_124 ));
    InMux I__3603 (
            .O(N__23925),
            .I(N__23922));
    LocalMux I__3602 (
            .O(N__23922),
            .I(N__23917));
    InMux I__3601 (
            .O(N__23921),
            .I(N__23912));
    InMux I__3600 (
            .O(N__23920),
            .I(N__23912));
    Span4Mux_v I__3599 (
            .O(N__23917),
            .I(N__23907));
    LocalMux I__3598 (
            .O(N__23912),
            .I(N__23907));
    Odrv4 I__3597 (
            .O(N__23907),
            .I(\pid_alt.pid_preregZ0Z_8 ));
    CascadeMux I__3596 (
            .O(N__23904),
            .I(N__23901));
    InMux I__3595 (
            .O(N__23901),
            .I(N__23898));
    LocalMux I__3594 (
            .O(N__23898),
            .I(N__23895));
    Odrv4 I__3593 (
            .O(N__23895),
            .I(\pid_alt.N_12_i ));
    InMux I__3592 (
            .O(N__23892),
            .I(N__23888));
    InMux I__3591 (
            .O(N__23891),
            .I(N__23885));
    LocalMux I__3590 (
            .O(N__23888),
            .I(N__23882));
    LocalMux I__3589 (
            .O(N__23885),
            .I(\pid_alt.un9lto29_i_a2_3_and ));
    Odrv4 I__3588 (
            .O(N__23882),
            .I(\pid_alt.un9lto29_i_a2_3_and ));
    CascadeMux I__3587 (
            .O(N__23877),
            .I(N__23874));
    InMux I__3586 (
            .O(N__23874),
            .I(N__23871));
    LocalMux I__3585 (
            .O(N__23871),
            .I(N__23868));
    Odrv4 I__3584 (
            .O(N__23868),
            .I(\pid_alt.source_pid_1_sqmuxa_0_a2_1_0 ));
    InMux I__3583 (
            .O(N__23865),
            .I(N__23861));
    InMux I__3582 (
            .O(N__23864),
            .I(N__23858));
    LocalMux I__3581 (
            .O(N__23861),
            .I(N__23855));
    LocalMux I__3580 (
            .O(N__23858),
            .I(\pid_alt.un9lto29_i_a2_4_and ));
    Odrv4 I__3579 (
            .O(N__23855),
            .I(\pid_alt.un9lto29_i_a2_4_and ));
    InMux I__3578 (
            .O(N__23850),
            .I(N__23847));
    LocalMux I__3577 (
            .O(N__23847),
            .I(N__23844));
    Odrv4 I__3576 (
            .O(N__23844),
            .I(\pid_alt.source_pid_1_sqmuxa_0_a2_0_5 ));
    CascadeMux I__3575 (
            .O(N__23841),
            .I(\pid_alt.N_123_cascade_ ));
    InMux I__3574 (
            .O(N__23838),
            .I(N__23835));
    LocalMux I__3573 (
            .O(N__23835),
            .I(N__23832));
    Span4Mux_h I__3572 (
            .O(N__23832),
            .I(N__23826));
    InMux I__3571 (
            .O(N__23831),
            .I(N__23819));
    InMux I__3570 (
            .O(N__23830),
            .I(N__23819));
    InMux I__3569 (
            .O(N__23829),
            .I(N__23819));
    Odrv4 I__3568 (
            .O(N__23826),
            .I(\pid_alt.pid_preregZ0Z_12 ));
    LocalMux I__3567 (
            .O(N__23819),
            .I(\pid_alt.pid_preregZ0Z_12 ));
    InMux I__3566 (
            .O(N__23814),
            .I(N__23807));
    InMux I__3565 (
            .O(N__23813),
            .I(N__23807));
    InMux I__3564 (
            .O(N__23812),
            .I(N__23804));
    LocalMux I__3563 (
            .O(N__23807),
            .I(\pid_alt.N_123 ));
    LocalMux I__3562 (
            .O(N__23804),
            .I(\pid_alt.N_123 ));
    CascadeMux I__3561 (
            .O(N__23799),
            .I(\pid_alt.N_106_cascade_ ));
    InMux I__3560 (
            .O(N__23796),
            .I(N__23793));
    LocalMux I__3559 (
            .O(N__23793),
            .I(\pid_alt.source_pid_1_sqmuxa_0_a2_0 ));
    InMux I__3558 (
            .O(N__23790),
            .I(N__23787));
    LocalMux I__3557 (
            .O(N__23787),
            .I(\pid_alt.N_100 ));
    CascadeMux I__3556 (
            .O(N__23784),
            .I(\pid_alt.N_91_1_cascade_ ));
    CascadeMux I__3555 (
            .O(N__23781),
            .I(\Commands_frame_decoder.N_358_cascade_ ));
    CascadeMux I__3554 (
            .O(N__23778),
            .I(N__23773));
    CascadeMux I__3553 (
            .O(N__23777),
            .I(N__23770));
    InMux I__3552 (
            .O(N__23776),
            .I(N__23765));
    InMux I__3551 (
            .O(N__23773),
            .I(N__23765));
    InMux I__3550 (
            .O(N__23770),
            .I(N__23762));
    LocalMux I__3549 (
            .O(N__23765),
            .I(\Commands_frame_decoder.stateZ0Z_10 ));
    LocalMux I__3548 (
            .O(N__23762),
            .I(\Commands_frame_decoder.stateZ0Z_10 ));
    InMux I__3547 (
            .O(N__23757),
            .I(N__23754));
    LocalMux I__3546 (
            .O(N__23754),
            .I(N__23750));
    InMux I__3545 (
            .O(N__23753),
            .I(N__23747));
    Span4Mux_v I__3544 (
            .O(N__23750),
            .I(N__23744));
    LocalMux I__3543 (
            .O(N__23747),
            .I(\Commands_frame_decoder.stateZ0Z_3 ));
    Odrv4 I__3542 (
            .O(N__23744),
            .I(\Commands_frame_decoder.stateZ0Z_3 ));
    InMux I__3541 (
            .O(N__23739),
            .I(N__23736));
    LocalMux I__3540 (
            .O(N__23736),
            .I(N__23733));
    Span4Mux_h I__3539 (
            .O(N__23733),
            .I(N__23730));
    Odrv4 I__3538 (
            .O(N__23730),
            .I(\Commands_frame_decoder.source_CH2data_1_sqmuxa ));
    InMux I__3537 (
            .O(N__23727),
            .I(N__23724));
    LocalMux I__3536 (
            .O(N__23724),
            .I(\Commands_frame_decoder.N_327 ));
    CascadeMux I__3535 (
            .O(N__23721),
            .I(N__23718));
    InMux I__3534 (
            .O(N__23718),
            .I(N__23712));
    InMux I__3533 (
            .O(N__23717),
            .I(N__23712));
    LocalMux I__3532 (
            .O(N__23712),
            .I(\Commands_frame_decoder.stateZ0Z_2 ));
    InMux I__3531 (
            .O(N__23709),
            .I(N__23705));
    InMux I__3530 (
            .O(N__23708),
            .I(N__23702));
    LocalMux I__3529 (
            .O(N__23705),
            .I(N__23698));
    LocalMux I__3528 (
            .O(N__23702),
            .I(N__23695));
    InMux I__3527 (
            .O(N__23701),
            .I(N__23692));
    Span4Mux_h I__3526 (
            .O(N__23698),
            .I(N__23687));
    Span4Mux_v I__3525 (
            .O(N__23695),
            .I(N__23687));
    LocalMux I__3524 (
            .O(N__23692),
            .I(\Commands_frame_decoder.stateZ0Z_11 ));
    Odrv4 I__3523 (
            .O(N__23687),
            .I(\Commands_frame_decoder.stateZ0Z_11 ));
    CascadeMux I__3522 (
            .O(N__23682),
            .I(N__23679));
    InMux I__3521 (
            .O(N__23679),
            .I(N__23675));
    InMux I__3520 (
            .O(N__23678),
            .I(N__23672));
    LocalMux I__3519 (
            .O(N__23675),
            .I(\Commands_frame_decoder.stateZ0Z_7 ));
    LocalMux I__3518 (
            .O(N__23672),
            .I(\Commands_frame_decoder.stateZ0Z_7 ));
    InMux I__3517 (
            .O(N__23667),
            .I(N__23664));
    LocalMux I__3516 (
            .O(N__23664),
            .I(N__23660));
    InMux I__3515 (
            .O(N__23663),
            .I(N__23657));
    Span4Mux_v I__3514 (
            .O(N__23660),
            .I(N__23652));
    LocalMux I__3513 (
            .O(N__23657),
            .I(N__23652));
    Odrv4 I__3512 (
            .O(N__23652),
            .I(\Commands_frame_decoder.WDT8lt14_0 ));
    InMux I__3511 (
            .O(N__23649),
            .I(N__23644));
    InMux I__3510 (
            .O(N__23648),
            .I(N__23639));
    InMux I__3509 (
            .O(N__23647),
            .I(N__23639));
    LocalMux I__3508 (
            .O(N__23644),
            .I(\Commands_frame_decoder.WDTZ0Z_8 ));
    LocalMux I__3507 (
            .O(N__23639),
            .I(\Commands_frame_decoder.WDTZ0Z_8 ));
    InMux I__3506 (
            .O(N__23634),
            .I(bfn_9_6_0_));
    CascadeMux I__3505 (
            .O(N__23631),
            .I(N__23626));
    CascadeMux I__3504 (
            .O(N__23630),
            .I(N__23623));
    InMux I__3503 (
            .O(N__23629),
            .I(N__23620));
    InMux I__3502 (
            .O(N__23626),
            .I(N__23615));
    InMux I__3501 (
            .O(N__23623),
            .I(N__23615));
    LocalMux I__3500 (
            .O(N__23620),
            .I(\Commands_frame_decoder.WDTZ0Z_9 ));
    LocalMux I__3499 (
            .O(N__23615),
            .I(\Commands_frame_decoder.WDTZ0Z_9 ));
    InMux I__3498 (
            .O(N__23610),
            .I(\Commands_frame_decoder.un1_WDT_cry_8 ));
    CascadeMux I__3497 (
            .O(N__23607),
            .I(N__23602));
    InMux I__3496 (
            .O(N__23606),
            .I(N__23599));
    InMux I__3495 (
            .O(N__23605),
            .I(N__23594));
    InMux I__3494 (
            .O(N__23602),
            .I(N__23594));
    LocalMux I__3493 (
            .O(N__23599),
            .I(\Commands_frame_decoder.WDTZ0Z_10 ));
    LocalMux I__3492 (
            .O(N__23594),
            .I(\Commands_frame_decoder.WDTZ0Z_10 ));
    InMux I__3491 (
            .O(N__23589),
            .I(\Commands_frame_decoder.un1_WDT_cry_9 ));
    InMux I__3490 (
            .O(N__23586),
            .I(\Commands_frame_decoder.un1_WDT_cry_10 ));
    InMux I__3489 (
            .O(N__23583),
            .I(\Commands_frame_decoder.un1_WDT_cry_11 ));
    InMux I__3488 (
            .O(N__23580),
            .I(\Commands_frame_decoder.un1_WDT_cry_12 ));
    InMux I__3487 (
            .O(N__23577),
            .I(\Commands_frame_decoder.un1_WDT_cry_13 ));
    InMux I__3486 (
            .O(N__23574),
            .I(\Commands_frame_decoder.un1_WDT_cry_14 ));
    InMux I__3485 (
            .O(N__23571),
            .I(N__23568));
    LocalMux I__3484 (
            .O(N__23568),
            .I(uart_input_pc_c));
    InMux I__3483 (
            .O(N__23565),
            .I(N__23561));
    CascadeMux I__3482 (
            .O(N__23564),
            .I(N__23558));
    LocalMux I__3481 (
            .O(N__23561),
            .I(N__23555));
    InMux I__3480 (
            .O(N__23558),
            .I(N__23552));
    Odrv4 I__3479 (
            .O(N__23555),
            .I(\Commands_frame_decoder.state_0_sqmuxa ));
    LocalMux I__3478 (
            .O(N__23552),
            .I(\Commands_frame_decoder.state_0_sqmuxa ));
    InMux I__3477 (
            .O(N__23547),
            .I(N__23544));
    LocalMux I__3476 (
            .O(N__23544),
            .I(\Commands_frame_decoder.WDTZ0Z_0 ));
    InMux I__3475 (
            .O(N__23541),
            .I(N__23538));
    LocalMux I__3474 (
            .O(N__23538),
            .I(\Commands_frame_decoder.WDTZ0Z_1 ));
    InMux I__3473 (
            .O(N__23535),
            .I(\Commands_frame_decoder.un1_WDT_cry_0 ));
    InMux I__3472 (
            .O(N__23532),
            .I(N__23529));
    LocalMux I__3471 (
            .O(N__23529),
            .I(\Commands_frame_decoder.WDTZ0Z_2 ));
    InMux I__3470 (
            .O(N__23526),
            .I(\Commands_frame_decoder.un1_WDT_cry_1 ));
    InMux I__3469 (
            .O(N__23523),
            .I(N__23520));
    LocalMux I__3468 (
            .O(N__23520),
            .I(\Commands_frame_decoder.WDTZ0Z_3 ));
    InMux I__3467 (
            .O(N__23517),
            .I(\Commands_frame_decoder.un1_WDT_cry_2 ));
    InMux I__3466 (
            .O(N__23514),
            .I(N__23509));
    InMux I__3465 (
            .O(N__23513),
            .I(N__23504));
    InMux I__3464 (
            .O(N__23512),
            .I(N__23504));
    LocalMux I__3463 (
            .O(N__23509),
            .I(\Commands_frame_decoder.WDTZ0Z_4 ));
    LocalMux I__3462 (
            .O(N__23504),
            .I(\Commands_frame_decoder.WDTZ0Z_4 ));
    InMux I__3461 (
            .O(N__23499),
            .I(\Commands_frame_decoder.un1_WDT_cry_3 ));
    InMux I__3460 (
            .O(N__23496),
            .I(N__23491));
    InMux I__3459 (
            .O(N__23495),
            .I(N__23486));
    InMux I__3458 (
            .O(N__23494),
            .I(N__23486));
    LocalMux I__3457 (
            .O(N__23491),
            .I(\Commands_frame_decoder.WDTZ0Z_5 ));
    LocalMux I__3456 (
            .O(N__23486),
            .I(\Commands_frame_decoder.WDTZ0Z_5 ));
    InMux I__3455 (
            .O(N__23481),
            .I(\Commands_frame_decoder.un1_WDT_cry_4 ));
    InMux I__3454 (
            .O(N__23478),
            .I(N__23473));
    InMux I__3453 (
            .O(N__23477),
            .I(N__23470));
    InMux I__3452 (
            .O(N__23476),
            .I(N__23467));
    LocalMux I__3451 (
            .O(N__23473),
            .I(\Commands_frame_decoder.WDTZ0Z_6 ));
    LocalMux I__3450 (
            .O(N__23470),
            .I(\Commands_frame_decoder.WDTZ0Z_6 ));
    LocalMux I__3449 (
            .O(N__23467),
            .I(\Commands_frame_decoder.WDTZ0Z_6 ));
    InMux I__3448 (
            .O(N__23460),
            .I(\Commands_frame_decoder.un1_WDT_cry_5 ));
    InMux I__3447 (
            .O(N__23457),
            .I(N__23452));
    InMux I__3446 (
            .O(N__23456),
            .I(N__23449));
    InMux I__3445 (
            .O(N__23455),
            .I(N__23446));
    LocalMux I__3444 (
            .O(N__23452),
            .I(\Commands_frame_decoder.WDTZ0Z_7 ));
    LocalMux I__3443 (
            .O(N__23449),
            .I(\Commands_frame_decoder.WDTZ0Z_7 ));
    LocalMux I__3442 (
            .O(N__23446),
            .I(\Commands_frame_decoder.WDTZ0Z_7 ));
    InMux I__3441 (
            .O(N__23439),
            .I(\Commands_frame_decoder.un1_WDT_cry_6 ));
    CascadeMux I__3440 (
            .O(N__23436),
            .I(N__23433));
    InMux I__3439 (
            .O(N__23433),
            .I(N__23430));
    LocalMux I__3438 (
            .O(N__23430),
            .I(\pid_alt.error_axbZ0Z_1 ));
    CascadeMux I__3437 (
            .O(N__23427),
            .I(N__23424));
    InMux I__3436 (
            .O(N__23424),
            .I(N__23421));
    LocalMux I__3435 (
            .O(N__23421),
            .I(\pid_alt.error_axbZ0Z_12 ));
    CascadeMux I__3434 (
            .O(N__23418),
            .I(N__23415));
    InMux I__3433 (
            .O(N__23415),
            .I(N__23412));
    LocalMux I__3432 (
            .O(N__23412),
            .I(\pid_alt.error_axbZ0Z_13 ));
    CascadeMux I__3431 (
            .O(N__23409),
            .I(N__23406));
    InMux I__3430 (
            .O(N__23406),
            .I(N__23403));
    LocalMux I__3429 (
            .O(N__23403),
            .I(\pid_alt.error_axbZ0Z_14 ));
    CascadeMux I__3428 (
            .O(N__23400),
            .I(N__23397));
    InMux I__3427 (
            .O(N__23397),
            .I(N__23394));
    LocalMux I__3426 (
            .O(N__23394),
            .I(\pid_alt.error_axbZ0Z_2 ));
    InMux I__3425 (
            .O(N__23391),
            .I(N__23388));
    LocalMux I__3424 (
            .O(N__23388),
            .I(N__23385));
    Span4Mux_v I__3423 (
            .O(N__23385),
            .I(N__23382));
    Sp12to4 I__3422 (
            .O(N__23382),
            .I(N__23379));
    Span12Mux_s9_h I__3421 (
            .O(N__23379),
            .I(N__23376));
    Odrv12 I__3420 (
            .O(N__23376),
            .I(alt_ki_0));
    CascadeMux I__3419 (
            .O(N__23373),
            .I(N__23370));
    InMux I__3418 (
            .O(N__23370),
            .I(N__23367));
    LocalMux I__3417 (
            .O(N__23367),
            .I(drone_altitude_i_9));
    InMux I__3416 (
            .O(N__23364),
            .I(N__23360));
    InMux I__3415 (
            .O(N__23363),
            .I(N__23357));
    LocalMux I__3414 (
            .O(N__23360),
            .I(N__23354));
    LocalMux I__3413 (
            .O(N__23357),
            .I(alt_command_0));
    Odrv4 I__3412 (
            .O(N__23354),
            .I(alt_command_0));
    InMux I__3411 (
            .O(N__23349),
            .I(N__23346));
    LocalMux I__3410 (
            .O(N__23346),
            .I(N__23343));
    Span4Mux_h I__3409 (
            .O(N__23343),
            .I(N__23340));
    Span4Mux_h I__3408 (
            .O(N__23340),
            .I(N__23337));
    Odrv4 I__3407 (
            .O(N__23337),
            .I(\pid_alt.O_1_9 ));
    CascadeMux I__3406 (
            .O(N__23334),
            .I(N__23331));
    InMux I__3405 (
            .O(N__23331),
            .I(N__23325));
    InMux I__3404 (
            .O(N__23330),
            .I(N__23325));
    LocalMux I__3403 (
            .O(N__23325),
            .I(\pid_alt.error_d_reg_prevZ0Z_21 ));
    InMux I__3402 (
            .O(N__23322),
            .I(N__23313));
    InMux I__3401 (
            .O(N__23321),
            .I(N__23313));
    InMux I__3400 (
            .O(N__23320),
            .I(N__23313));
    LocalMux I__3399 (
            .O(N__23313),
            .I(N__23310));
    Span4Mux_h I__3398 (
            .O(N__23310),
            .I(N__23307));
    Span4Mux_h I__3397 (
            .O(N__23307),
            .I(N__23304));
    Sp12to4 I__3396 (
            .O(N__23304),
            .I(N__23301));
    Odrv12 I__3395 (
            .O(N__23301),
            .I(\pid_alt.error_d_regZ0Z_21 ));
    InMux I__3394 (
            .O(N__23298),
            .I(N__23295));
    LocalMux I__3393 (
            .O(N__23295),
            .I(\pid_alt.error_d_reg_prev_esr_RNIIIKM_0Z0Z_21 ));
    CascadeMux I__3392 (
            .O(N__23292),
            .I(N__23288));
    InMux I__3391 (
            .O(N__23291),
            .I(N__23285));
    InMux I__3390 (
            .O(N__23288),
            .I(N__23282));
    LocalMux I__3389 (
            .O(N__23285),
            .I(\pid_alt.error_d_reg_prev_esr_RNIS5212Z0Z_19 ));
    LocalMux I__3388 (
            .O(N__23282),
            .I(\pid_alt.error_d_reg_prev_esr_RNIS5212Z0Z_19 ));
    InMux I__3387 (
            .O(N__23277),
            .I(N__23271));
    InMux I__3386 (
            .O(N__23276),
            .I(N__23271));
    LocalMux I__3385 (
            .O(N__23271),
            .I(N__23268));
    Span4Mux_h I__3384 (
            .O(N__23268),
            .I(N__23265));
    Span4Mux_h I__3383 (
            .O(N__23265),
            .I(N__23262));
    Odrv4 I__3382 (
            .O(N__23262),
            .I(\pid_alt.error_d_reg_prev_esr_RNIGGKMZ0Z_20 ));
    CascadeMux I__3381 (
            .O(N__23259),
            .I(\pid_alt.error_d_reg_prev_esr_RNIIIKM_0Z0Z_21_cascade_ ));
    InMux I__3380 (
            .O(N__23256),
            .I(N__23253));
    LocalMux I__3379 (
            .O(N__23253),
            .I(N__23250));
    Span4Mux_h I__3378 (
            .O(N__23250),
            .I(N__23247));
    Odrv4 I__3377 (
            .O(N__23247),
            .I(\pid_alt.error_d_reg_prev_esr_RNIQ8034Z0Z_20 ));
    CascadeMux I__3376 (
            .O(N__23244),
            .I(N__23240));
    InMux I__3375 (
            .O(N__23243),
            .I(N__23237));
    InMux I__3374 (
            .O(N__23240),
            .I(N__23234));
    LocalMux I__3373 (
            .O(N__23237),
            .I(\pid_alt.drone_altitude_i_0 ));
    LocalMux I__3372 (
            .O(N__23234),
            .I(\pid_alt.drone_altitude_i_0 ));
    CascadeMux I__3371 (
            .O(N__23229),
            .I(N__23226));
    InMux I__3370 (
            .O(N__23226),
            .I(N__23223));
    LocalMux I__3369 (
            .O(N__23223),
            .I(\pid_alt.error_axbZ0Z_3 ));
    CascadeMux I__3368 (
            .O(N__23220),
            .I(N__23217));
    InMux I__3367 (
            .O(N__23217),
            .I(N__23214));
    LocalMux I__3366 (
            .O(N__23214),
            .I(drone_altitude_i_10));
    CascadeMux I__3365 (
            .O(N__23211),
            .I(N__23208));
    InMux I__3364 (
            .O(N__23208),
            .I(N__23205));
    LocalMux I__3363 (
            .O(N__23205),
            .I(drone_altitude_i_11));
    InMux I__3362 (
            .O(N__23202),
            .I(N__23199));
    LocalMux I__3361 (
            .O(N__23199),
            .I(N__23196));
    Span4Mux_h I__3360 (
            .O(N__23196),
            .I(N__23192));
    InMux I__3359 (
            .O(N__23195),
            .I(N__23189));
    Odrv4 I__3358 (
            .O(N__23192),
            .I(\pid_alt.error_d_reg_prev_esr_RNIGGKM_0Z0Z_20 ));
    LocalMux I__3357 (
            .O(N__23189),
            .I(\pid_alt.error_d_reg_prev_esr_RNIGGKM_0Z0Z_20 ));
    InMux I__3356 (
            .O(N__23184),
            .I(N__23181));
    LocalMux I__3355 (
            .O(N__23181),
            .I(N__23178));
    Span4Mux_h I__3354 (
            .O(N__23178),
            .I(N__23175));
    Span4Mux_h I__3353 (
            .O(N__23175),
            .I(N__23171));
    InMux I__3352 (
            .O(N__23174),
            .I(N__23168));
    Odrv4 I__3351 (
            .O(N__23171),
            .I(\pid_alt.error_d_reg_prev_esr_RNI86IMZ0Z_19 ));
    LocalMux I__3350 (
            .O(N__23168),
            .I(\pid_alt.error_d_reg_prev_esr_RNI86IMZ0Z_19 ));
    InMux I__3349 (
            .O(N__23163),
            .I(N__23160));
    LocalMux I__3348 (
            .O(N__23160),
            .I(N__23157));
    Odrv12 I__3347 (
            .O(N__23157),
            .I(\dron_frame_decoder_1.state_RNI3T3K1Z0Z_7 ));
    InMux I__3346 (
            .O(N__23154),
            .I(N__23150));
    InMux I__3345 (
            .O(N__23153),
            .I(N__23147));
    LocalMux I__3344 (
            .O(N__23150),
            .I(N__23144));
    LocalMux I__3343 (
            .O(N__23147),
            .I(\pid_alt.error_d_reg_prevZ0Z_26 ));
    Odrv4 I__3342 (
            .O(N__23144),
            .I(\pid_alt.error_d_reg_prevZ0Z_26 ));
    InMux I__3341 (
            .O(N__23139),
            .I(N__23133));
    InMux I__3340 (
            .O(N__23138),
            .I(N__23133));
    LocalMux I__3339 (
            .O(N__23133),
            .I(N__23129));
    InMux I__3338 (
            .O(N__23132),
            .I(N__23126));
    Span4Mux_v I__3337 (
            .O(N__23129),
            .I(N__23123));
    LocalMux I__3336 (
            .O(N__23126),
            .I(N__23120));
    Span4Mux_v I__3335 (
            .O(N__23123),
            .I(N__23117));
    Span4Mux_h I__3334 (
            .O(N__23120),
            .I(N__23114));
    Span4Mux_v I__3333 (
            .O(N__23117),
            .I(N__23111));
    Sp12to4 I__3332 (
            .O(N__23114),
            .I(N__23108));
    Sp12to4 I__3331 (
            .O(N__23111),
            .I(N__23103));
    Span12Mux_v I__3330 (
            .O(N__23108),
            .I(N__23103));
    Odrv12 I__3329 (
            .O(N__23103),
            .I(\pid_alt.error_d_regZ0Z_26 ));
    InMux I__3328 (
            .O(N__23100),
            .I(N__23097));
    LocalMux I__3327 (
            .O(N__23097),
            .I(\pid_alt.error_d_reg_prev_esr_RNIL8611Z0Z_9 ));
    InMux I__3326 (
            .O(N__23094),
            .I(N__23090));
    InMux I__3325 (
            .O(N__23093),
            .I(N__23087));
    LocalMux I__3324 (
            .O(N__23090),
            .I(\pid_alt.error_d_reg_prev_esr_RNIDAHM_0Z0Z_10 ));
    LocalMux I__3323 (
            .O(N__23087),
            .I(\pid_alt.error_d_reg_prev_esr_RNIDAHM_0Z0Z_10 ));
    CascadeMux I__3322 (
            .O(N__23082),
            .I(N__23078));
    CascadeMux I__3321 (
            .O(N__23081),
            .I(N__23075));
    InMux I__3320 (
            .O(N__23078),
            .I(N__23072));
    InMux I__3319 (
            .O(N__23075),
            .I(N__23069));
    LocalMux I__3318 (
            .O(N__23072),
            .I(N__23066));
    LocalMux I__3317 (
            .O(N__23069),
            .I(N__23063));
    Span4Mux_v I__3316 (
            .O(N__23066),
            .I(N__23060));
    Span4Mux_h I__3315 (
            .O(N__23063),
            .I(N__23057));
    Odrv4 I__3314 (
            .O(N__23060),
            .I(\pid_alt.error_d_reg_prev_esr_RNISAR62Z0Z_9 ));
    Odrv4 I__3313 (
            .O(N__23057),
            .I(\pid_alt.error_d_reg_prev_esr_RNISAR62Z0Z_9 ));
    InMux I__3312 (
            .O(N__23052),
            .I(N__23049));
    LocalMux I__3311 (
            .O(N__23049),
            .I(N__23046));
    Span4Mux_v I__3310 (
            .O(N__23046),
            .I(N__23042));
    InMux I__3309 (
            .O(N__23045),
            .I(N__23039));
    Odrv4 I__3308 (
            .O(N__23042),
            .I(\pid_alt.error_d_reg_prev_esr_RNI27U12Z0Z_21 ));
    LocalMux I__3307 (
            .O(N__23039),
            .I(\pid_alt.error_d_reg_prev_esr_RNI27U12Z0Z_21 ));
    InMux I__3306 (
            .O(N__23034),
            .I(N__23031));
    LocalMux I__3305 (
            .O(N__23031),
            .I(\pid_alt.error_d_reg_prev_esr_RNIIIKMZ0Z_21 ));
    InMux I__3304 (
            .O(N__23028),
            .I(N__23022));
    InMux I__3303 (
            .O(N__23027),
            .I(N__23022));
    LocalMux I__3302 (
            .O(N__23022),
            .I(N__23019));
    Span4Mux_h I__3301 (
            .O(N__23019),
            .I(N__23016));
    Odrv4 I__3300 (
            .O(N__23016),
            .I(\pid_alt.error_d_reg_prev_esr_RNIKKKM_0Z0Z_22 ));
    CascadeMux I__3299 (
            .O(N__23013),
            .I(\pid_alt.error_d_reg_prev_esr_RNIIIKMZ0Z_21_cascade_ ));
    CascadeMux I__3298 (
            .O(N__23010),
            .I(N__23007));
    InMux I__3297 (
            .O(N__23007),
            .I(N__23004));
    LocalMux I__3296 (
            .O(N__23004),
            .I(N__23001));
    Odrv4 I__3295 (
            .O(N__23001),
            .I(\pid_alt.error_d_reg_prev_esr_RNI0AS34Z0Z_21 ));
    InMux I__3294 (
            .O(N__22998),
            .I(N__22994));
    InMux I__3293 (
            .O(N__22997),
            .I(N__22991));
    LocalMux I__3292 (
            .O(N__22994),
            .I(N__22988));
    LocalMux I__3291 (
            .O(N__22991),
            .I(\pid_alt.error_d_reg_prev_esr_RNIU2U12Z0Z_20 ));
    Odrv4 I__3290 (
            .O(N__22988),
            .I(\pid_alt.error_d_reg_prev_esr_RNIU2U12Z0Z_20 ));
    CascadeMux I__3289 (
            .O(N__22983),
            .I(\pid_alt.error_d_reg_prev_esr_RNIL8611Z0Z_9_cascade_ ));
    InMux I__3288 (
            .O(N__22980),
            .I(N__22977));
    LocalMux I__3287 (
            .O(N__22977),
            .I(\pid_alt.error_d_reg_prev_esr_RNICI045Z0Z_9 ));
    InMux I__3286 (
            .O(N__22974),
            .I(N__22971));
    LocalMux I__3285 (
            .O(N__22971),
            .I(N__22967));
    InMux I__3284 (
            .O(N__22970),
            .I(N__22964));
    Span4Mux_v I__3283 (
            .O(N__22967),
            .I(N__22959));
    LocalMux I__3282 (
            .O(N__22964),
            .I(N__22959));
    Span4Mux_h I__3281 (
            .O(N__22959),
            .I(N__22956));
    Span4Mux_h I__3280 (
            .O(N__22956),
            .I(N__22953));
    Odrv4 I__3279 (
            .O(N__22953),
            .I(\pid_alt.error_p_regZ0Z_10 ));
    InMux I__3278 (
            .O(N__22950),
            .I(N__22947));
    LocalMux I__3277 (
            .O(N__22947),
            .I(N__22943));
    InMux I__3276 (
            .O(N__22946),
            .I(N__22940));
    Span4Mux_v I__3275 (
            .O(N__22943),
            .I(N__22937));
    LocalMux I__3274 (
            .O(N__22940),
            .I(\pid_alt.error_d_reg_prevZ0Z_10 ));
    Odrv4 I__3273 (
            .O(N__22937),
            .I(\pid_alt.error_d_reg_prevZ0Z_10 ));
    InMux I__3272 (
            .O(N__22932),
            .I(N__22927));
    InMux I__3271 (
            .O(N__22931),
            .I(N__22922));
    InMux I__3270 (
            .O(N__22930),
            .I(N__22922));
    LocalMux I__3269 (
            .O(N__22927),
            .I(N__22919));
    LocalMux I__3268 (
            .O(N__22922),
            .I(N__22916));
    Span4Mux_v I__3267 (
            .O(N__22919),
            .I(N__22913));
    Span4Mux_h I__3266 (
            .O(N__22916),
            .I(N__22910));
    Span4Mux_h I__3265 (
            .O(N__22913),
            .I(N__22907));
    Odrv4 I__3264 (
            .O(N__22910),
            .I(\pid_alt.error_d_regZ0Z_10 ));
    Odrv4 I__3263 (
            .O(N__22907),
            .I(\pid_alt.error_d_regZ0Z_10 ));
    CascadeMux I__3262 (
            .O(N__22902),
            .I(N__22898));
    InMux I__3261 (
            .O(N__22901),
            .I(N__22895));
    InMux I__3260 (
            .O(N__22898),
            .I(N__22892));
    LocalMux I__3259 (
            .O(N__22895),
            .I(\pid_alt.error_d_reg_prev_esr_RNIG75T2Z0Z_8 ));
    LocalMux I__3258 (
            .O(N__22892),
            .I(\pid_alt.error_d_reg_prev_esr_RNIG75T2Z0Z_8 ));
    InMux I__3257 (
            .O(N__22887),
            .I(N__22881));
    InMux I__3256 (
            .O(N__22886),
            .I(N__22881));
    LocalMux I__3255 (
            .O(N__22881),
            .I(N__22878));
    Span4Mux_h I__3254 (
            .O(N__22878),
            .I(N__22875));
    Span4Mux_v I__3253 (
            .O(N__22875),
            .I(N__22872));
    Span4Mux_h I__3252 (
            .O(N__22872),
            .I(N__22869));
    Odrv4 I__3251 (
            .O(N__22869),
            .I(\pid_alt.error_p_regZ0Z_9 ));
    CascadeMux I__3250 (
            .O(N__22866),
            .I(N__22863));
    InMux I__3249 (
            .O(N__22863),
            .I(N__22857));
    InMux I__3248 (
            .O(N__22862),
            .I(N__22857));
    LocalMux I__3247 (
            .O(N__22857),
            .I(\pid_alt.error_d_reg_prevZ0Z_9 ));
    InMux I__3246 (
            .O(N__22854),
            .I(N__22845));
    InMux I__3245 (
            .O(N__22853),
            .I(N__22845));
    InMux I__3244 (
            .O(N__22852),
            .I(N__22845));
    LocalMux I__3243 (
            .O(N__22845),
            .I(N__22842));
    Span4Mux_v I__3242 (
            .O(N__22842),
            .I(N__22839));
    Span4Mux_h I__3241 (
            .O(N__22839),
            .I(N__22836));
    Span4Mux_h I__3240 (
            .O(N__22836),
            .I(N__22833));
    Odrv4 I__3239 (
            .O(N__22833),
            .I(\pid_alt.error_d_regZ0Z_9 ));
    InMux I__3238 (
            .O(N__22830),
            .I(N__22827));
    LocalMux I__3237 (
            .O(N__22827),
            .I(\pid_alt.error_d_reg_prev_esr_RNIL8611_0Z0Z_9 ));
    InMux I__3236 (
            .O(N__22824),
            .I(N__22818));
    InMux I__3235 (
            .O(N__22823),
            .I(N__22818));
    LocalMux I__3234 (
            .O(N__22818),
            .I(N__22815));
    Span4Mux_h I__3233 (
            .O(N__22815),
            .I(N__22812));
    Odrv4 I__3232 (
            .O(N__22812),
            .I(\pid_alt.error_d_reg_prev_esr_RNII5611Z0Z_8 ));
    InMux I__3231 (
            .O(N__22809),
            .I(N__22805));
    CascadeMux I__3230 (
            .O(N__22808),
            .I(N__22802));
    LocalMux I__3229 (
            .O(N__22805),
            .I(N__22799));
    InMux I__3228 (
            .O(N__22802),
            .I(N__22796));
    Span4Mux_v I__3227 (
            .O(N__22799),
            .I(N__22793));
    LocalMux I__3226 (
            .O(N__22796),
            .I(N__22790));
    Span4Mux_v I__3225 (
            .O(N__22793),
            .I(N__22785));
    Span4Mux_v I__3224 (
            .O(N__22790),
            .I(N__22785));
    Odrv4 I__3223 (
            .O(N__22785),
            .I(\pid_alt.error_d_reg_prev_esr_RNI7T3T2Z0Z_7 ));
    CascadeMux I__3222 (
            .O(N__22782),
            .I(\pid_alt.error_d_reg_prev_esr_RNIL8611_0Z0Z_9_cascade_ ));
    InMux I__3221 (
            .O(N__22779),
            .I(N__22776));
    LocalMux I__3220 (
            .O(N__22776),
            .I(\pid_alt.error_d_reg_prev_esr_RNIN49Q5Z0Z_8 ));
    CascadeMux I__3219 (
            .O(N__22773),
            .I(N__22769));
    CascadeMux I__3218 (
            .O(N__22772),
            .I(N__22766));
    InMux I__3217 (
            .O(N__22769),
            .I(N__22763));
    InMux I__3216 (
            .O(N__22766),
            .I(N__22760));
    LocalMux I__3215 (
            .O(N__22763),
            .I(N__22755));
    LocalMux I__3214 (
            .O(N__22760),
            .I(N__22755));
    Odrv4 I__3213 (
            .O(N__22755),
            .I(\pid_alt.error_d_reg_prev_esr_RNIL81T2Z0Z_5 ));
    InMux I__3212 (
            .O(N__22752),
            .I(N__22749));
    LocalMux I__3211 (
            .O(N__22749),
            .I(N__22746));
    Span4Mux_h I__3210 (
            .O(N__22746),
            .I(N__22743));
    Odrv4 I__3209 (
            .O(N__22743),
            .I(\pid_alt.error_d_reg_prev_esr_RNIJR3Q5Z0Z_6 ));
    CascadeMux I__3208 (
            .O(N__22740),
            .I(N__22736));
    InMux I__3207 (
            .O(N__22739),
            .I(N__22733));
    InMux I__3206 (
            .O(N__22736),
            .I(N__22730));
    LocalMux I__3205 (
            .O(N__22733),
            .I(N__22727));
    LocalMux I__3204 (
            .O(N__22730),
            .I(N__22724));
    Span4Mux_v I__3203 (
            .O(N__22727),
            .I(N__22719));
    Span4Mux_h I__3202 (
            .O(N__22724),
            .I(N__22719));
    Odrv4 I__3201 (
            .O(N__22719),
            .I(\pid_alt.pid_preregZ0Z_29 ));
    InMux I__3200 (
            .O(N__22716),
            .I(N__22710));
    InMux I__3199 (
            .O(N__22715),
            .I(N__22710));
    LocalMux I__3198 (
            .O(N__22710),
            .I(\pid_alt.pid_preregZ0Z_14 ));
    InMux I__3197 (
            .O(N__22707),
            .I(N__22704));
    LocalMux I__3196 (
            .O(N__22704),
            .I(\pid_alt.error_d_reg_prev_esr_RNICV511_0Z0Z_6 ));
    CascadeMux I__3195 (
            .O(N__22701),
            .I(\pid_alt.error_d_reg_prev_esr_RNICV511_0Z0Z_6_cascade_ ));
    InMux I__3194 (
            .O(N__22698),
            .I(N__22695));
    LocalMux I__3193 (
            .O(N__22695),
            .I(\pid_alt.error_d_reg_prev_esr_RNI171A6Z0Z_5 ));
    CascadeMux I__3192 (
            .O(N__22692),
            .I(N__22688));
    InMux I__3191 (
            .O(N__22691),
            .I(N__22685));
    InMux I__3190 (
            .O(N__22688),
            .I(N__22682));
    LocalMux I__3189 (
            .O(N__22685),
            .I(\pid_alt.error_d_reg_prev_esr_RNICUVC3Z0Z_4 ));
    LocalMux I__3188 (
            .O(N__22682),
            .I(\pid_alt.error_d_reg_prev_esr_RNICUVC3Z0Z_4 ));
    InMux I__3187 (
            .O(N__22677),
            .I(N__22674));
    LocalMux I__3186 (
            .O(N__22674),
            .I(\pid_alt.error_d_reg_prev_esr_RNI9S511_0Z0Z_5 ));
    CascadeMux I__3185 (
            .O(N__22671),
            .I(\pid_alt.error_d_reg_prev_esr_RNI9S511_0Z0Z_5_cascade_ ));
    InMux I__3184 (
            .O(N__22668),
            .I(N__22665));
    LocalMux I__3183 (
            .O(N__22665),
            .I(\pid_alt.error_d_reg_prev_esr_RNIOGSO6Z0Z_4 ));
    CascadeMux I__3182 (
            .O(N__22662),
            .I(N__22659));
    InMux I__3181 (
            .O(N__22659),
            .I(N__22656));
    LocalMux I__3180 (
            .O(N__22656),
            .I(\pid_alt.N_232_i ));
    InMux I__3179 (
            .O(N__22653),
            .I(bfn_8_12_0_));
    InMux I__3178 (
            .O(N__22650),
            .I(N__22644));
    InMux I__3177 (
            .O(N__22649),
            .I(N__22641));
    InMux I__3176 (
            .O(N__22648),
            .I(N__22636));
    InMux I__3175 (
            .O(N__22647),
            .I(N__22636));
    LocalMux I__3174 (
            .O(N__22644),
            .I(\dron_frame_decoder_1.stateZ0Z_0 ));
    LocalMux I__3173 (
            .O(N__22641),
            .I(\dron_frame_decoder_1.stateZ0Z_0 ));
    LocalMux I__3172 (
            .O(N__22636),
            .I(\dron_frame_decoder_1.stateZ0Z_0 ));
    InMux I__3171 (
            .O(N__22629),
            .I(N__22626));
    LocalMux I__3170 (
            .O(N__22626),
            .I(\dron_frame_decoder_1.state_ns_i_i_a2_2_0_0 ));
    InMux I__3169 (
            .O(N__22623),
            .I(N__22620));
    LocalMux I__3168 (
            .O(N__22620),
            .I(N__22617));
    Odrv4 I__3167 (
            .O(N__22617),
            .I(\pid_alt.pid_preregZ0Z_22 ));
    InMux I__3166 (
            .O(N__22614),
            .I(N__22611));
    LocalMux I__3165 (
            .O(N__22611),
            .I(N__22608));
    Odrv4 I__3164 (
            .O(N__22608),
            .I(\pid_alt.pid_preregZ0Z_21 ));
    CascadeMux I__3163 (
            .O(N__22605),
            .I(N__22602));
    InMux I__3162 (
            .O(N__22602),
            .I(N__22599));
    LocalMux I__3161 (
            .O(N__22599),
            .I(N__22596));
    Odrv4 I__3160 (
            .O(N__22596),
            .I(\pid_alt.pid_preregZ0Z_23 ));
    InMux I__3159 (
            .O(N__22593),
            .I(N__22590));
    LocalMux I__3158 (
            .O(N__22590),
            .I(N__22587));
    Odrv4 I__3157 (
            .O(N__22587),
            .I(\pid_alt.pid_preregZ0Z_20 ));
    InMux I__3156 (
            .O(N__22584),
            .I(N__22581));
    LocalMux I__3155 (
            .O(N__22581),
            .I(N__22578));
    Odrv4 I__3154 (
            .O(N__22578),
            .I(\pid_alt.source_pid10lt4_0 ));
    InMux I__3153 (
            .O(N__22575),
            .I(N__22572));
    LocalMux I__3152 (
            .O(N__22572),
            .I(N__22569));
    Odrv4 I__3151 (
            .O(N__22569),
            .I(\pid_alt.un9lto29_i_a2_2_and ));
    InMux I__3150 (
            .O(N__22566),
            .I(N__22562));
    InMux I__3149 (
            .O(N__22565),
            .I(N__22559));
    LocalMux I__3148 (
            .O(N__22562),
            .I(N__22556));
    LocalMux I__3147 (
            .O(N__22559),
            .I(N__22553));
    Odrv12 I__3146 (
            .O(N__22556),
            .I(\pid_alt.pid_preregZ0Z_28 ));
    Odrv4 I__3145 (
            .O(N__22553),
            .I(\pid_alt.pid_preregZ0Z_28 ));
    CascadeMux I__3144 (
            .O(N__22548),
            .I(N__22545));
    InMux I__3143 (
            .O(N__22545),
            .I(N__22539));
    InMux I__3142 (
            .O(N__22544),
            .I(N__22539));
    LocalMux I__3141 (
            .O(N__22539),
            .I(N__22536));
    Odrv4 I__3140 (
            .O(N__22536),
            .I(\pid_alt.pid_preregZ0Z_15 ));
    InMux I__3139 (
            .O(N__22533),
            .I(N__22522));
    InMux I__3138 (
            .O(N__22532),
            .I(N__22522));
    InMux I__3137 (
            .O(N__22531),
            .I(N__22522));
    InMux I__3136 (
            .O(N__22530),
            .I(N__22517));
    InMux I__3135 (
            .O(N__22529),
            .I(N__22517));
    LocalMux I__3134 (
            .O(N__22522),
            .I(N__22509));
    LocalMux I__3133 (
            .O(N__22517),
            .I(N__22509));
    InMux I__3132 (
            .O(N__22516),
            .I(N__22502));
    InMux I__3131 (
            .O(N__22515),
            .I(N__22502));
    InMux I__3130 (
            .O(N__22514),
            .I(N__22502));
    Span4Mux_v I__3129 (
            .O(N__22509),
            .I(N__22497));
    LocalMux I__3128 (
            .O(N__22502),
            .I(N__22497));
    Odrv4 I__3127 (
            .O(N__22497),
            .I(\dron_frame_decoder_1.WDT_RNIPI9R2Z0Z_15 ));
    InMux I__3126 (
            .O(N__22494),
            .I(N__22485));
    InMux I__3125 (
            .O(N__22493),
            .I(N__22485));
    InMux I__3124 (
            .O(N__22492),
            .I(N__22485));
    LocalMux I__3123 (
            .O(N__22485),
            .I(\dron_frame_decoder_1.stateZ0Z_7 ));
    CEMux I__3122 (
            .O(N__22482),
            .I(N__22478));
    CEMux I__3121 (
            .O(N__22481),
            .I(N__22475));
    LocalMux I__3120 (
            .O(N__22478),
            .I(N__22467));
    LocalMux I__3119 (
            .O(N__22475),
            .I(N__22467));
    CEMux I__3118 (
            .O(N__22474),
            .I(N__22464));
    CEMux I__3117 (
            .O(N__22473),
            .I(N__22461));
    CEMux I__3116 (
            .O(N__22472),
            .I(N__22458));
    Span4Mux_v I__3115 (
            .O(N__22467),
            .I(N__22451));
    LocalMux I__3114 (
            .O(N__22464),
            .I(N__22451));
    LocalMux I__3113 (
            .O(N__22461),
            .I(N__22451));
    LocalMux I__3112 (
            .O(N__22458),
            .I(N__22448));
    Span4Mux_v I__3111 (
            .O(N__22451),
            .I(N__22443));
    Span4Mux_v I__3110 (
            .O(N__22448),
            .I(N__22443));
    Span4Mux_v I__3109 (
            .O(N__22443),
            .I(N__22440));
    Span4Mux_h I__3108 (
            .O(N__22440),
            .I(N__22437));
    Span4Mux_v I__3107 (
            .O(N__22437),
            .I(N__22434));
    Odrv4 I__3106 (
            .O(N__22434),
            .I(\Commands_frame_decoder.state_RNIF38SZ0Z_6 ));
    CascadeMux I__3105 (
            .O(N__22431),
            .I(N__22428));
    InMux I__3104 (
            .O(N__22428),
            .I(N__22425));
    LocalMux I__3103 (
            .O(N__22425),
            .I(N__22422));
    Odrv4 I__3102 (
            .O(N__22422),
            .I(\Commands_frame_decoder.N_354 ));
    InMux I__3101 (
            .O(N__22419),
            .I(N__22416));
    LocalMux I__3100 (
            .O(N__22416),
            .I(\Commands_frame_decoder.source_offset2data_1_sqmuxa ));
    InMux I__3099 (
            .O(N__22413),
            .I(N__22407));
    InMux I__3098 (
            .O(N__22412),
            .I(N__22407));
    LocalMux I__3097 (
            .O(N__22407),
            .I(\Commands_frame_decoder.stateZ0Z_8 ));
    CascadeMux I__3096 (
            .O(N__22404),
            .I(N__22401));
    InMux I__3095 (
            .O(N__22401),
            .I(N__22398));
    LocalMux I__3094 (
            .O(N__22398),
            .I(\dron_frame_decoder_1.un1_sink_data_valid_5_i_0 ));
    CascadeMux I__3093 (
            .O(N__22395),
            .I(\dron_frame_decoder_1.un1_sink_data_valid_5_i_0_cascade_ ));
    InMux I__3092 (
            .O(N__22392),
            .I(N__22386));
    InMux I__3091 (
            .O(N__22391),
            .I(N__22383));
    InMux I__3090 (
            .O(N__22390),
            .I(N__22378));
    InMux I__3089 (
            .O(N__22389),
            .I(N__22378));
    LocalMux I__3088 (
            .O(N__22386),
            .I(\dron_frame_decoder_1.stateZ0Z_5 ));
    LocalMux I__3087 (
            .O(N__22383),
            .I(\dron_frame_decoder_1.stateZ0Z_5 ));
    LocalMux I__3086 (
            .O(N__22378),
            .I(\dron_frame_decoder_1.stateZ0Z_5 ));
    CascadeMux I__3085 (
            .O(N__22371),
            .I(N__22368));
    InMux I__3084 (
            .O(N__22368),
            .I(N__22363));
    InMux I__3083 (
            .O(N__22367),
            .I(N__22358));
    InMux I__3082 (
            .O(N__22366),
            .I(N__22358));
    LocalMux I__3081 (
            .O(N__22363),
            .I(\dron_frame_decoder_1.stateZ0Z_4 ));
    LocalMux I__3080 (
            .O(N__22358),
            .I(\dron_frame_decoder_1.stateZ0Z_4 ));
    CascadeMux I__3079 (
            .O(N__22353),
            .I(\Commands_frame_decoder.WDT8lt12_0_cascade_ ));
    InMux I__3078 (
            .O(N__22350),
            .I(N__22347));
    LocalMux I__3077 (
            .O(N__22347),
            .I(\Commands_frame_decoder.state_0_sqmuxacf1 ));
    InMux I__3076 (
            .O(N__22344),
            .I(N__22341));
    LocalMux I__3075 (
            .O(N__22341),
            .I(\Commands_frame_decoder.WDT_RNII19A1Z0Z_4 ));
    InMux I__3074 (
            .O(N__22338),
            .I(N__22335));
    LocalMux I__3073 (
            .O(N__22335),
            .I(N__22332));
    Odrv4 I__3072 (
            .O(N__22332),
            .I(\uart_drone_sync.aux_2__0__0_0 ));
    InMux I__3071 (
            .O(N__22329),
            .I(N__22326));
    LocalMux I__3070 (
            .O(N__22326),
            .I(\uart_drone_sync.aux_3__0__0_0 ));
    SRMux I__3069 (
            .O(N__22323),
            .I(N__22319));
    SRMux I__3068 (
            .O(N__22322),
            .I(N__22316));
    LocalMux I__3067 (
            .O(N__22319),
            .I(N__22313));
    LocalMux I__3066 (
            .O(N__22316),
            .I(N__22310));
    Span4Mux_h I__3065 (
            .O(N__22313),
            .I(N__22307));
    Span4Mux_h I__3064 (
            .O(N__22310),
            .I(N__22304));
    Odrv4 I__3063 (
            .O(N__22307),
            .I(\dron_frame_decoder_1.source_data_valid_2_sqmuxa_iZ0 ));
    Odrv4 I__3062 (
            .O(N__22304),
            .I(\dron_frame_decoder_1.source_data_valid_2_sqmuxa_iZ0 ));
    CascadeMux I__3061 (
            .O(N__22299),
            .I(\Commands_frame_decoder.source_offset2data_1_sqmuxa_cascade_ ));
    CascadeMux I__3060 (
            .O(N__22296),
            .I(\Commands_frame_decoder.N_322_0_cascade_ ));
    IoInMux I__3059 (
            .O(N__22293),
            .I(N__22290));
    LocalMux I__3058 (
            .O(N__22290),
            .I(N__22287));
    Span4Mux_s1_v I__3057 (
            .O(N__22287),
            .I(N__22284));
    Odrv4 I__3056 (
            .O(N__22284),
            .I(\pid_alt.N_410_0 ));
    InMux I__3055 (
            .O(N__22281),
            .I(N__22278));
    LocalMux I__3054 (
            .O(N__22278),
            .I(\uart_drone_sync.aux_1__0__0_0 ));
    InMux I__3053 (
            .O(N__22275),
            .I(N__22272));
    LocalMux I__3052 (
            .O(N__22272),
            .I(N__22269));
    Odrv4 I__3051 (
            .O(N__22269),
            .I(uart_input_drone_c));
    InMux I__3050 (
            .O(N__22266),
            .I(N__22263));
    LocalMux I__3049 (
            .O(N__22263),
            .I(\uart_drone_sync.aux_0__0__0_0 ));
    CascadeMux I__3048 (
            .O(N__22260),
            .I(\Commands_frame_decoder.WDT8lto13_1_cascade_ ));
    InMux I__3047 (
            .O(N__22257),
            .I(N__22254));
    LocalMux I__3046 (
            .O(N__22254),
            .I(\Commands_frame_decoder.WDT_RNI2VDI1Z0Z_10 ));
    CascadeMux I__3045 (
            .O(N__22251),
            .I(\Commands_frame_decoder.WDT8lto9_3_cascade_ ));
    InMux I__3044 (
            .O(N__22248),
            .I(N__22244));
    InMux I__3043 (
            .O(N__22247),
            .I(N__22240));
    LocalMux I__3042 (
            .O(N__22244),
            .I(N__22237));
    InMux I__3041 (
            .O(N__22243),
            .I(N__22234));
    LocalMux I__3040 (
            .O(N__22240),
            .I(N__22231));
    Span12Mux_s6_h I__3039 (
            .O(N__22237),
            .I(N__22228));
    LocalMux I__3038 (
            .O(N__22234),
            .I(N__22225));
    Span4Mux_v I__3037 (
            .O(N__22231),
            .I(N__22222));
    Span12Mux_h I__3036 (
            .O(N__22228),
            .I(N__22217));
    Span12Mux_s7_h I__3035 (
            .O(N__22225),
            .I(N__22217));
    Span4Mux_h I__3034 (
            .O(N__22222),
            .I(N__22214));
    Odrv12 I__3033 (
            .O(N__22217),
            .I(\pid_alt.error_13 ));
    Odrv4 I__3032 (
            .O(N__22214),
            .I(\pid_alt.error_13 ));
    InMux I__3031 (
            .O(N__22209),
            .I(\pid_alt.error_cry_12 ));
    InMux I__3030 (
            .O(N__22206),
            .I(N__22203));
    LocalMux I__3029 (
            .O(N__22203),
            .I(N__22200));
    Span4Mux_s2_h I__3028 (
            .O(N__22200),
            .I(N__22197));
    Span4Mux_h I__3027 (
            .O(N__22197),
            .I(N__22193));
    InMux I__3026 (
            .O(N__22196),
            .I(N__22190));
    Span4Mux_h I__3025 (
            .O(N__22193),
            .I(N__22186));
    LocalMux I__3024 (
            .O(N__22190),
            .I(N__22183));
    InMux I__3023 (
            .O(N__22189),
            .I(N__22180));
    Span4Mux_h I__3022 (
            .O(N__22186),
            .I(N__22177));
    Span4Mux_s3_h I__3021 (
            .O(N__22183),
            .I(N__22174));
    LocalMux I__3020 (
            .O(N__22180),
            .I(N__22171));
    Span4Mux_h I__3019 (
            .O(N__22177),
            .I(N__22166));
    Span4Mux_h I__3018 (
            .O(N__22174),
            .I(N__22166));
    Span4Mux_s3_h I__3017 (
            .O(N__22171),
            .I(N__22163));
    Span4Mux_v I__3016 (
            .O(N__22166),
            .I(N__22158));
    Span4Mux_h I__3015 (
            .O(N__22163),
            .I(N__22158));
    Odrv4 I__3014 (
            .O(N__22158),
            .I(\pid_alt.error_14 ));
    InMux I__3013 (
            .O(N__22155),
            .I(\pid_alt.error_cry_13 ));
    InMux I__3012 (
            .O(N__22152),
            .I(\pid_alt.error_cry_14 ));
    InMux I__3011 (
            .O(N__22149),
            .I(N__22146));
    LocalMux I__3010 (
            .O(N__22146),
            .I(N__22143));
    Span4Mux_s2_h I__3009 (
            .O(N__22143),
            .I(N__22140));
    Span4Mux_h I__3008 (
            .O(N__22140),
            .I(N__22136));
    InMux I__3007 (
            .O(N__22139),
            .I(N__22133));
    Span4Mux_h I__3006 (
            .O(N__22136),
            .I(N__22129));
    LocalMux I__3005 (
            .O(N__22133),
            .I(N__22126));
    InMux I__3004 (
            .O(N__22132),
            .I(N__22123));
    Span4Mux_h I__3003 (
            .O(N__22129),
            .I(N__22120));
    Span4Mux_s3_h I__3002 (
            .O(N__22126),
            .I(N__22117));
    LocalMux I__3001 (
            .O(N__22123),
            .I(N__22114));
    Span4Mux_h I__3000 (
            .O(N__22120),
            .I(N__22109));
    Span4Mux_h I__2999 (
            .O(N__22117),
            .I(N__22109));
    Span4Mux_s3_h I__2998 (
            .O(N__22114),
            .I(N__22106));
    Span4Mux_v I__2997 (
            .O(N__22109),
            .I(N__22101));
    Span4Mux_h I__2996 (
            .O(N__22106),
            .I(N__22101));
    Odrv4 I__2995 (
            .O(N__22101),
            .I(\pid_alt.error_15 ));
    InMux I__2994 (
            .O(N__22098),
            .I(N__22095));
    LocalMux I__2993 (
            .O(N__22095),
            .I(alt_command_4));
    InMux I__2992 (
            .O(N__22092),
            .I(N__22089));
    LocalMux I__2991 (
            .O(N__22089),
            .I(N__22086));
    Odrv4 I__2990 (
            .O(N__22086),
            .I(alt_command_5));
    InMux I__2989 (
            .O(N__22083),
            .I(N__22080));
    LocalMux I__2988 (
            .O(N__22080),
            .I(N__22077));
    Odrv4 I__2987 (
            .O(N__22077),
            .I(alt_command_6));
    InMux I__2986 (
            .O(N__22074),
            .I(N__22071));
    LocalMux I__2985 (
            .O(N__22071),
            .I(alt_command_7));
    CascadeMux I__2984 (
            .O(N__22068),
            .I(N__22065));
    InMux I__2983 (
            .O(N__22065),
            .I(N__22062));
    LocalMux I__2982 (
            .O(N__22062),
            .I(N__22059));
    Span4Mux_v I__2981 (
            .O(N__22059),
            .I(N__22056));
    Odrv4 I__2980 (
            .O(N__22056),
            .I(\pid_alt.error_d_reg_prev_esr_RNIOTU12Z0Z_27 ));
    CascadeMux I__2979 (
            .O(N__22053),
            .I(N__22048));
    InMux I__2978 (
            .O(N__22052),
            .I(N__22044));
    InMux I__2977 (
            .O(N__22051),
            .I(N__22041));
    InMux I__2976 (
            .O(N__22048),
            .I(N__22038));
    InMux I__2975 (
            .O(N__22047),
            .I(N__22035));
    LocalMux I__2974 (
            .O(N__22044),
            .I(N__22030));
    LocalMux I__2973 (
            .O(N__22041),
            .I(N__22030));
    LocalMux I__2972 (
            .O(N__22038),
            .I(\pid_alt.error_d_reg_prev_esr_RNIUUKMZ0Z_27 ));
    LocalMux I__2971 (
            .O(N__22035),
            .I(\pid_alt.error_d_reg_prev_esr_RNIUUKMZ0Z_27 ));
    Odrv12 I__2970 (
            .O(N__22030),
            .I(\pid_alt.error_d_reg_prev_esr_RNIUUKMZ0Z_27 ));
    InMux I__2969 (
            .O(N__22023),
            .I(N__22019));
    InMux I__2968 (
            .O(N__22022),
            .I(N__22016));
    LocalMux I__2967 (
            .O(N__22019),
            .I(N__22010));
    LocalMux I__2966 (
            .O(N__22016),
            .I(N__22010));
    InMux I__2965 (
            .O(N__22015),
            .I(N__22005));
    Span4Mux_v I__2964 (
            .O(N__22010),
            .I(N__22002));
    InMux I__2963 (
            .O(N__22009),
            .I(N__21997));
    InMux I__2962 (
            .O(N__22008),
            .I(N__21997));
    LocalMux I__2961 (
            .O(N__22005),
            .I(\pid_alt.un1_pid_prereg_296_1 ));
    Odrv4 I__2960 (
            .O(N__22002),
            .I(\pid_alt.un1_pid_prereg_296_1 ));
    LocalMux I__2959 (
            .O(N__21997),
            .I(\pid_alt.un1_pid_prereg_296_1 ));
    InMux I__2958 (
            .O(N__21990),
            .I(N__21987));
    LocalMux I__2957 (
            .O(N__21987),
            .I(N__21984));
    Span4Mux_v I__2956 (
            .O(N__21984),
            .I(N__21981));
    Odrv4 I__2955 (
            .O(N__21981),
            .I(\pid_alt.error_d_reg_prev_esr_RNIOTU12_0Z0Z_27 ));
    InMux I__2954 (
            .O(N__21978),
            .I(N__21974));
    InMux I__2953 (
            .O(N__21977),
            .I(N__21971));
    LocalMux I__2952 (
            .O(N__21974),
            .I(N__21968));
    LocalMux I__2951 (
            .O(N__21971),
            .I(alt_command_1));
    Odrv4 I__2950 (
            .O(N__21968),
            .I(alt_command_1));
    InMux I__2949 (
            .O(N__21963),
            .I(N__21960));
    LocalMux I__2948 (
            .O(N__21960),
            .I(N__21957));
    Span4Mux_s2_h I__2947 (
            .O(N__21957),
            .I(N__21954));
    Span4Mux_h I__2946 (
            .O(N__21954),
            .I(N__21950));
    InMux I__2945 (
            .O(N__21953),
            .I(N__21947));
    Span4Mux_h I__2944 (
            .O(N__21950),
            .I(N__21943));
    LocalMux I__2943 (
            .O(N__21947),
            .I(N__21940));
    InMux I__2942 (
            .O(N__21946),
            .I(N__21937));
    Span4Mux_h I__2941 (
            .O(N__21943),
            .I(N__21934));
    Span4Mux_s3_h I__2940 (
            .O(N__21940),
            .I(N__21931));
    LocalMux I__2939 (
            .O(N__21937),
            .I(N__21928));
    Span4Mux_h I__2938 (
            .O(N__21934),
            .I(N__21923));
    Span4Mux_h I__2937 (
            .O(N__21931),
            .I(N__21923));
    Span4Mux_s3_h I__2936 (
            .O(N__21928),
            .I(N__21920));
    Span4Mux_v I__2935 (
            .O(N__21923),
            .I(N__21915));
    Span4Mux_h I__2934 (
            .O(N__21920),
            .I(N__21915));
    Odrv4 I__2933 (
            .O(N__21915),
            .I(\pid_alt.error_5 ));
    InMux I__2932 (
            .O(N__21912),
            .I(\pid_alt.error_cry_4 ));
    CascadeMux I__2931 (
            .O(N__21909),
            .I(N__21905));
    CascadeMux I__2930 (
            .O(N__21908),
            .I(N__21902));
    InMux I__2929 (
            .O(N__21905),
            .I(N__21899));
    InMux I__2928 (
            .O(N__21902),
            .I(N__21896));
    LocalMux I__2927 (
            .O(N__21899),
            .I(alt_command_2));
    LocalMux I__2926 (
            .O(N__21896),
            .I(alt_command_2));
    InMux I__2925 (
            .O(N__21891),
            .I(N__21886));
    InMux I__2924 (
            .O(N__21890),
            .I(N__21883));
    InMux I__2923 (
            .O(N__21889),
            .I(N__21880));
    LocalMux I__2922 (
            .O(N__21886),
            .I(N__21877));
    LocalMux I__2921 (
            .O(N__21883),
            .I(N__21874));
    LocalMux I__2920 (
            .O(N__21880),
            .I(N__21871));
    Span12Mux_s6_h I__2919 (
            .O(N__21877),
            .I(N__21868));
    Span4Mux_s3_h I__2918 (
            .O(N__21874),
            .I(N__21865));
    Span12Mux_s7_h I__2917 (
            .O(N__21871),
            .I(N__21860));
    Span12Mux_h I__2916 (
            .O(N__21868),
            .I(N__21860));
    Span4Mux_h I__2915 (
            .O(N__21865),
            .I(N__21857));
    Odrv12 I__2914 (
            .O(N__21860),
            .I(\pid_alt.error_6 ));
    Odrv4 I__2913 (
            .O(N__21857),
            .I(\pid_alt.error_6 ));
    InMux I__2912 (
            .O(N__21852),
            .I(\pid_alt.error_cry_5 ));
    InMux I__2911 (
            .O(N__21849),
            .I(N__21845));
    InMux I__2910 (
            .O(N__21848),
            .I(N__21842));
    LocalMux I__2909 (
            .O(N__21845),
            .I(alt_command_3));
    LocalMux I__2908 (
            .O(N__21842),
            .I(alt_command_3));
    InMux I__2907 (
            .O(N__21837),
            .I(N__21834));
    LocalMux I__2906 (
            .O(N__21834),
            .I(N__21831));
    Span4Mux_s2_h I__2905 (
            .O(N__21831),
            .I(N__21827));
    InMux I__2904 (
            .O(N__21830),
            .I(N__21824));
    Span4Mux_h I__2903 (
            .O(N__21827),
            .I(N__21821));
    LocalMux I__2902 (
            .O(N__21824),
            .I(N__21817));
    Span4Mux_h I__2901 (
            .O(N__21821),
            .I(N__21814));
    InMux I__2900 (
            .O(N__21820),
            .I(N__21811));
    Span4Mux_s3_h I__2899 (
            .O(N__21817),
            .I(N__21808));
    Span4Mux_h I__2898 (
            .O(N__21814),
            .I(N__21805));
    LocalMux I__2897 (
            .O(N__21811),
            .I(N__21802));
    Span4Mux_h I__2896 (
            .O(N__21808),
            .I(N__21799));
    Span4Mux_h I__2895 (
            .O(N__21805),
            .I(N__21796));
    Span4Mux_s3_h I__2894 (
            .O(N__21802),
            .I(N__21793));
    Span4Mux_v I__2893 (
            .O(N__21799),
            .I(N__21786));
    Span4Mux_v I__2892 (
            .O(N__21796),
            .I(N__21786));
    Span4Mux_h I__2891 (
            .O(N__21793),
            .I(N__21786));
    Odrv4 I__2890 (
            .O(N__21786),
            .I(\pid_alt.error_7 ));
    InMux I__2889 (
            .O(N__21783),
            .I(\pid_alt.error_cry_6 ));
    InMux I__2888 (
            .O(N__21780),
            .I(N__21777));
    LocalMux I__2887 (
            .O(N__21777),
            .I(N__21774));
    Span4Mux_s2_h I__2886 (
            .O(N__21774),
            .I(N__21771));
    Span4Mux_h I__2885 (
            .O(N__21771),
            .I(N__21767));
    InMux I__2884 (
            .O(N__21770),
            .I(N__21764));
    Span4Mux_h I__2883 (
            .O(N__21767),
            .I(N__21760));
    LocalMux I__2882 (
            .O(N__21764),
            .I(N__21757));
    InMux I__2881 (
            .O(N__21763),
            .I(N__21754));
    Span4Mux_h I__2880 (
            .O(N__21760),
            .I(N__21751));
    Span4Mux_s3_h I__2879 (
            .O(N__21757),
            .I(N__21748));
    LocalMux I__2878 (
            .O(N__21754),
            .I(N__21745));
    Span4Mux_h I__2877 (
            .O(N__21751),
            .I(N__21740));
    Span4Mux_h I__2876 (
            .O(N__21748),
            .I(N__21740));
    Span4Mux_s3_h I__2875 (
            .O(N__21745),
            .I(N__21737));
    Span4Mux_v I__2874 (
            .O(N__21740),
            .I(N__21732));
    Span4Mux_h I__2873 (
            .O(N__21737),
            .I(N__21732));
    Odrv4 I__2872 (
            .O(N__21732),
            .I(\pid_alt.error_8 ));
    InMux I__2871 (
            .O(N__21729),
            .I(bfn_7_20_0_));
    InMux I__2870 (
            .O(N__21726),
            .I(N__21723));
    LocalMux I__2869 (
            .O(N__21723),
            .I(N__21720));
    Span4Mux_s2_h I__2868 (
            .O(N__21720),
            .I(N__21717));
    Span4Mux_h I__2867 (
            .O(N__21717),
            .I(N__21713));
    InMux I__2866 (
            .O(N__21716),
            .I(N__21710));
    Span4Mux_h I__2865 (
            .O(N__21713),
            .I(N__21706));
    LocalMux I__2864 (
            .O(N__21710),
            .I(N__21703));
    InMux I__2863 (
            .O(N__21709),
            .I(N__21700));
    Span4Mux_h I__2862 (
            .O(N__21706),
            .I(N__21697));
    Span4Mux_s3_h I__2861 (
            .O(N__21703),
            .I(N__21694));
    LocalMux I__2860 (
            .O(N__21700),
            .I(N__21691));
    Span4Mux_h I__2859 (
            .O(N__21697),
            .I(N__21686));
    Span4Mux_h I__2858 (
            .O(N__21694),
            .I(N__21686));
    Span4Mux_s3_h I__2857 (
            .O(N__21691),
            .I(N__21683));
    Span4Mux_v I__2856 (
            .O(N__21686),
            .I(N__21678));
    Span4Mux_h I__2855 (
            .O(N__21683),
            .I(N__21678));
    Odrv4 I__2854 (
            .O(N__21678),
            .I(\pid_alt.error_9 ));
    InMux I__2853 (
            .O(N__21675),
            .I(\pid_alt.error_cry_8 ));
    InMux I__2852 (
            .O(N__21672),
            .I(N__21669));
    LocalMux I__2851 (
            .O(N__21669),
            .I(N__21665));
    InMux I__2850 (
            .O(N__21668),
            .I(N__21661));
    Span4Mux_v I__2849 (
            .O(N__21665),
            .I(N__21658));
    InMux I__2848 (
            .O(N__21664),
            .I(N__21655));
    LocalMux I__2847 (
            .O(N__21661),
            .I(N__21652));
    Span4Mux_v I__2846 (
            .O(N__21658),
            .I(N__21647));
    LocalMux I__2845 (
            .O(N__21655),
            .I(N__21647));
    Span12Mux_s10_v I__2844 (
            .O(N__21652),
            .I(N__21644));
    Span4Mux_h I__2843 (
            .O(N__21647),
            .I(N__21641));
    Span12Mux_h I__2842 (
            .O(N__21644),
            .I(N__21638));
    Span4Mux_h I__2841 (
            .O(N__21641),
            .I(N__21635));
    Odrv12 I__2840 (
            .O(N__21638),
            .I(\pid_alt.error_10 ));
    Odrv4 I__2839 (
            .O(N__21635),
            .I(\pid_alt.error_10 ));
    InMux I__2838 (
            .O(N__21630),
            .I(\pid_alt.error_cry_9 ));
    InMux I__2837 (
            .O(N__21627),
            .I(N__21624));
    LocalMux I__2836 (
            .O(N__21624),
            .I(N__21621));
    Span4Mux_s1_h I__2835 (
            .O(N__21621),
            .I(N__21617));
    InMux I__2834 (
            .O(N__21620),
            .I(N__21613));
    Sp12to4 I__2833 (
            .O(N__21617),
            .I(N__21610));
    InMux I__2832 (
            .O(N__21616),
            .I(N__21607));
    LocalMux I__2831 (
            .O(N__21613),
            .I(N__21604));
    Span12Mux_s10_v I__2830 (
            .O(N__21610),
            .I(N__21601));
    LocalMux I__2829 (
            .O(N__21607),
            .I(N__21598));
    Span4Mux_s3_h I__2828 (
            .O(N__21604),
            .I(N__21595));
    Span12Mux_h I__2827 (
            .O(N__21601),
            .I(N__21590));
    Span12Mux_s10_v I__2826 (
            .O(N__21598),
            .I(N__21590));
    Span4Mux_h I__2825 (
            .O(N__21595),
            .I(N__21587));
    Odrv12 I__2824 (
            .O(N__21590),
            .I(\pid_alt.error_11 ));
    Odrv4 I__2823 (
            .O(N__21587),
            .I(\pid_alt.error_11 ));
    InMux I__2822 (
            .O(N__21582),
            .I(\pid_alt.error_cry_10 ));
    InMux I__2821 (
            .O(N__21579),
            .I(N__21576));
    LocalMux I__2820 (
            .O(N__21576),
            .I(N__21573));
    Span4Mux_v I__2819 (
            .O(N__21573),
            .I(N__21570));
    Span4Mux_h I__2818 (
            .O(N__21570),
            .I(N__21566));
    InMux I__2817 (
            .O(N__21569),
            .I(N__21563));
    Span4Mux_h I__2816 (
            .O(N__21566),
            .I(N__21559));
    LocalMux I__2815 (
            .O(N__21563),
            .I(N__21556));
    InMux I__2814 (
            .O(N__21562),
            .I(N__21553));
    Span4Mux_h I__2813 (
            .O(N__21559),
            .I(N__21550));
    Span4Mux_v I__2812 (
            .O(N__21556),
            .I(N__21547));
    LocalMux I__2811 (
            .O(N__21553),
            .I(N__21544));
    Span4Mux_h I__2810 (
            .O(N__21550),
            .I(N__21541));
    Span4Mux_v I__2809 (
            .O(N__21547),
            .I(N__21536));
    Span4Mux_v I__2808 (
            .O(N__21544),
            .I(N__21536));
    Span4Mux_v I__2807 (
            .O(N__21541),
            .I(N__21531));
    Span4Mux_h I__2806 (
            .O(N__21536),
            .I(N__21531));
    Odrv4 I__2805 (
            .O(N__21531),
            .I(\pid_alt.error_12 ));
    InMux I__2804 (
            .O(N__21528),
            .I(\pid_alt.error_cry_11 ));
    InMux I__2803 (
            .O(N__21525),
            .I(N__21516));
    InMux I__2802 (
            .O(N__21524),
            .I(N__21516));
    InMux I__2801 (
            .O(N__21523),
            .I(N__21516));
    LocalMux I__2800 (
            .O(N__21516),
            .I(N__21513));
    Span4Mux_h I__2799 (
            .O(N__21513),
            .I(N__21510));
    Span4Mux_h I__2798 (
            .O(N__21510),
            .I(N__21507));
    Span4Mux_v I__2797 (
            .O(N__21507),
            .I(N__21504));
    Span4Mux_v I__2796 (
            .O(N__21504),
            .I(N__21501));
    Odrv4 I__2795 (
            .O(N__21501),
            .I(\pid_alt.error_d_regZ0Z_27 ));
    CascadeMux I__2794 (
            .O(N__21498),
            .I(N__21495));
    InMux I__2793 (
            .O(N__21495),
            .I(N__21489));
    InMux I__2792 (
            .O(N__21494),
            .I(N__21489));
    LocalMux I__2791 (
            .O(N__21489),
            .I(\pid_alt.error_d_reg_prevZ0Z_27 ));
    InMux I__2790 (
            .O(N__21486),
            .I(N__21482));
    InMux I__2789 (
            .O(N__21485),
            .I(N__21479));
    LocalMux I__2788 (
            .O(N__21482),
            .I(N__21476));
    LocalMux I__2787 (
            .O(N__21479),
            .I(N__21473));
    Span4Mux_v I__2786 (
            .O(N__21476),
            .I(N__21469));
    Span4Mux_v I__2785 (
            .O(N__21473),
            .I(N__21466));
    InMux I__2784 (
            .O(N__21472),
            .I(N__21463));
    Span4Mux_h I__2783 (
            .O(N__21469),
            .I(N__21460));
    Span4Mux_v I__2782 (
            .O(N__21466),
            .I(N__21455));
    LocalMux I__2781 (
            .O(N__21463),
            .I(N__21455));
    Sp12to4 I__2780 (
            .O(N__21460),
            .I(N__21452));
    Span4Mux_h I__2779 (
            .O(N__21455),
            .I(N__21449));
    Span12Mux_h I__2778 (
            .O(N__21452),
            .I(N__21446));
    Span4Mux_h I__2777 (
            .O(N__21449),
            .I(N__21443));
    Odrv12 I__2776 (
            .O(N__21446),
            .I(\pid_alt.error_1 ));
    Odrv4 I__2775 (
            .O(N__21443),
            .I(\pid_alt.error_1 ));
    InMux I__2774 (
            .O(N__21438),
            .I(\pid_alt.error_cry_0 ));
    InMux I__2773 (
            .O(N__21435),
            .I(N__21431));
    InMux I__2772 (
            .O(N__21434),
            .I(N__21427));
    LocalMux I__2771 (
            .O(N__21431),
            .I(N__21424));
    InMux I__2770 (
            .O(N__21430),
            .I(N__21421));
    LocalMux I__2769 (
            .O(N__21427),
            .I(N__21418));
    Span4Mux_v I__2768 (
            .O(N__21424),
            .I(N__21415));
    LocalMux I__2767 (
            .O(N__21421),
            .I(N__21412));
    Span12Mux_s11_v I__2766 (
            .O(N__21418),
            .I(N__21409));
    Span4Mux_v I__2765 (
            .O(N__21415),
            .I(N__21404));
    Span4Mux_v I__2764 (
            .O(N__21412),
            .I(N__21404));
    Span12Mux_h I__2763 (
            .O(N__21409),
            .I(N__21401));
    Span4Mux_h I__2762 (
            .O(N__21404),
            .I(N__21398));
    Odrv12 I__2761 (
            .O(N__21401),
            .I(\pid_alt.error_2 ));
    Odrv4 I__2760 (
            .O(N__21398),
            .I(\pid_alt.error_2 ));
    InMux I__2759 (
            .O(N__21393),
            .I(\pid_alt.error_cry_1 ));
    InMux I__2758 (
            .O(N__21390),
            .I(N__21387));
    LocalMux I__2757 (
            .O(N__21387),
            .I(N__21384));
    Span4Mux_v I__2756 (
            .O(N__21384),
            .I(N__21380));
    InMux I__2755 (
            .O(N__21383),
            .I(N__21376));
    Span4Mux_h I__2754 (
            .O(N__21380),
            .I(N__21373));
    InMux I__2753 (
            .O(N__21379),
            .I(N__21370));
    LocalMux I__2752 (
            .O(N__21376),
            .I(N__21367));
    Sp12to4 I__2751 (
            .O(N__21373),
            .I(N__21364));
    LocalMux I__2750 (
            .O(N__21370),
            .I(N__21361));
    Span4Mux_v I__2749 (
            .O(N__21367),
            .I(N__21358));
    Span12Mux_h I__2748 (
            .O(N__21364),
            .I(N__21355));
    Span12Mux_s11_v I__2747 (
            .O(N__21361),
            .I(N__21352));
    Span4Mux_h I__2746 (
            .O(N__21358),
            .I(N__21349));
    Odrv12 I__2745 (
            .O(N__21355),
            .I(\pid_alt.error_3 ));
    Odrv12 I__2744 (
            .O(N__21352),
            .I(\pid_alt.error_3 ));
    Odrv4 I__2743 (
            .O(N__21349),
            .I(\pid_alt.error_3 ));
    InMux I__2742 (
            .O(N__21342),
            .I(\pid_alt.error_cry_2 ));
    InMux I__2741 (
            .O(N__21339),
            .I(N__21336));
    LocalMux I__2740 (
            .O(N__21336),
            .I(N__21333));
    Span4Mux_s2_h I__2739 (
            .O(N__21333),
            .I(N__21330));
    Span4Mux_h I__2738 (
            .O(N__21330),
            .I(N__21326));
    InMux I__2737 (
            .O(N__21329),
            .I(N__21323));
    Span4Mux_h I__2736 (
            .O(N__21326),
            .I(N__21319));
    LocalMux I__2735 (
            .O(N__21323),
            .I(N__21316));
    InMux I__2734 (
            .O(N__21322),
            .I(N__21313));
    Span4Mux_h I__2733 (
            .O(N__21319),
            .I(N__21310));
    Span4Mux_s3_h I__2732 (
            .O(N__21316),
            .I(N__21307));
    LocalMux I__2731 (
            .O(N__21313),
            .I(N__21304));
    Span4Mux_h I__2730 (
            .O(N__21310),
            .I(N__21299));
    Span4Mux_h I__2729 (
            .O(N__21307),
            .I(N__21299));
    Span4Mux_s3_h I__2728 (
            .O(N__21304),
            .I(N__21296));
    Span4Mux_v I__2727 (
            .O(N__21299),
            .I(N__21291));
    Span4Mux_h I__2726 (
            .O(N__21296),
            .I(N__21291));
    Odrv4 I__2725 (
            .O(N__21291),
            .I(\pid_alt.error_4 ));
    InMux I__2724 (
            .O(N__21288),
            .I(\pid_alt.error_cry_3 ));
    InMux I__2723 (
            .O(N__21285),
            .I(\pid_alt.un1_pid_prereg_0_cry_28 ));
    InMux I__2722 (
            .O(N__21282),
            .I(\pid_alt.un1_pid_prereg_0_cry_29 ));
    InMux I__2721 (
            .O(N__21279),
            .I(N__21276));
    LocalMux I__2720 (
            .O(N__21276),
            .I(\pid_alt.error_d_reg_prev_esr_RNI8JT34Z0Z_26 ));
    CascadeMux I__2719 (
            .O(N__21273),
            .I(\pid_alt.error_d_reg_prev_esr_RNISSKMZ0Z_26_cascade_ ));
    InMux I__2718 (
            .O(N__21270),
            .I(N__21267));
    LocalMux I__2717 (
            .O(N__21267),
            .I(N__21264));
    Odrv4 I__2716 (
            .O(N__21264),
            .I(\pid_alt.error_d_reg_prev_esr_RNIMRU12Z0Z_26 ));
    InMux I__2715 (
            .O(N__21261),
            .I(N__21257));
    InMux I__2714 (
            .O(N__21260),
            .I(N__21254));
    LocalMux I__2713 (
            .O(N__21257),
            .I(\pid_alt.error_d_reg_prev_esr_RNISSKMZ0Z_26 ));
    LocalMux I__2712 (
            .O(N__21254),
            .I(\pid_alt.error_d_reg_prev_esr_RNISSKMZ0Z_26 ));
    CascadeMux I__2711 (
            .O(N__21249),
            .I(\pid_alt.un1_pid_prereg_296_1_cascade_ ));
    CascadeMux I__2710 (
            .O(N__21246),
            .I(N__21243));
    InMux I__2709 (
            .O(N__21243),
            .I(N__21240));
    LocalMux I__2708 (
            .O(N__21240),
            .I(\pid_alt.error_d_reg_prev_esr_RNIKQJO2Z0Z_26 ));
    InMux I__2707 (
            .O(N__21237),
            .I(N__21234));
    LocalMux I__2706 (
            .O(N__21234),
            .I(N__21231));
    Odrv12 I__2705 (
            .O(N__21231),
            .I(\pid_alt.error_d_reg_prev_esr_RNIK3024Z0Z_19 ));
    CascadeMux I__2704 (
            .O(N__21228),
            .I(N__21224));
    CascadeMux I__2703 (
            .O(N__21227),
            .I(N__21221));
    InMux I__2702 (
            .O(N__21224),
            .I(N__21218));
    InMux I__2701 (
            .O(N__21221),
            .I(N__21215));
    LocalMux I__2700 (
            .O(N__21218),
            .I(N__21212));
    LocalMux I__2699 (
            .O(N__21215),
            .I(\pid_alt.error_d_reg_prev_esr_RNIOTT02Z0Z_18 ));
    Odrv4 I__2698 (
            .O(N__21212),
            .I(\pid_alt.error_d_reg_prev_esr_RNIOTT02Z0Z_18 ));
    InMux I__2697 (
            .O(N__21207),
            .I(\pid_alt.un1_pid_prereg_0_cry_19 ));
    InMux I__2696 (
            .O(N__21204),
            .I(\pid_alt.un1_pid_prereg_0_cry_20 ));
    InMux I__2695 (
            .O(N__21201),
            .I(\pid_alt.un1_pid_prereg_0_cry_21 ));
    CascadeMux I__2694 (
            .O(N__21198),
            .I(N__21195));
    InMux I__2693 (
            .O(N__21195),
            .I(N__21192));
    LocalMux I__2692 (
            .O(N__21192),
            .I(N__21189));
    Span4Mux_v I__2691 (
            .O(N__21189),
            .I(N__21186));
    Odrv4 I__2690 (
            .O(N__21186),
            .I(\pid_alt.error_d_reg_prev_esr_RNI8IS34Z0Z_22 ));
    InMux I__2689 (
            .O(N__21183),
            .I(bfn_7_16_0_));
    InMux I__2688 (
            .O(N__21180),
            .I(\pid_alt.un1_pid_prereg_0_cry_23 ));
    InMux I__2687 (
            .O(N__21177),
            .I(\pid_alt.un1_pid_prereg_0_cry_24 ));
    InMux I__2686 (
            .O(N__21174),
            .I(\pid_alt.un1_pid_prereg_0_cry_25 ));
    InMux I__2685 (
            .O(N__21171),
            .I(\pid_alt.un1_pid_prereg_0_cry_26 ));
    InMux I__2684 (
            .O(N__21168),
            .I(\pid_alt.un1_pid_prereg_0_cry_27 ));
    InMux I__2683 (
            .O(N__21165),
            .I(N__21162));
    LocalMux I__2682 (
            .O(N__21162),
            .I(N__21159));
    Odrv4 I__2681 (
            .O(N__21159),
            .I(\pid_alt.error_d_reg_prev_esr_RNIP92N4Z0Z_11 ));
    CascadeMux I__2680 (
            .O(N__21156),
            .I(N__21153));
    InMux I__2679 (
            .O(N__21153),
            .I(N__21150));
    LocalMux I__2678 (
            .O(N__21150),
            .I(N__21147));
    Odrv4 I__2677 (
            .O(N__21147),
            .I(\pid_alt.error_d_reg_prev_esr_RNIOFGB2Z0Z_10 ));
    InMux I__2676 (
            .O(N__21144),
            .I(\pid_alt.un1_pid_prereg_0_cry_11 ));
    InMux I__2675 (
            .O(N__21141),
            .I(N__21138));
    LocalMux I__2674 (
            .O(N__21138),
            .I(N__21135));
    Span4Mux_v I__2673 (
            .O(N__21135),
            .I(N__21132));
    Span4Mux_h I__2672 (
            .O(N__21132),
            .I(N__21129));
    Odrv4 I__2671 (
            .O(N__21129),
            .I(\pid_alt.error_d_reg_prev_esr_RNIT4AF4Z0Z_12 ));
    CascadeMux I__2670 (
            .O(N__21126),
            .I(N__21123));
    InMux I__2669 (
            .O(N__21123),
            .I(N__21120));
    LocalMux I__2668 (
            .O(N__21120),
            .I(N__21116));
    InMux I__2667 (
            .O(N__21119),
            .I(N__21113));
    Span4Mux_h I__2666 (
            .O(N__21116),
            .I(N__21110));
    LocalMux I__2665 (
            .O(N__21113),
            .I(\pid_alt.error_d_reg_prev_esr_RNI1QHB2Z0Z_11 ));
    Odrv4 I__2664 (
            .O(N__21110),
            .I(\pid_alt.error_d_reg_prev_esr_RNI1QHB2Z0Z_11 ));
    InMux I__2663 (
            .O(N__21105),
            .I(\pid_alt.un1_pid_prereg_0_cry_12 ));
    InMux I__2662 (
            .O(N__21102),
            .I(N__21099));
    LocalMux I__2661 (
            .O(N__21099),
            .I(N__21096));
    Span4Mux_h I__2660 (
            .O(N__21096),
            .I(N__21093));
    Odrv4 I__2659 (
            .O(N__21093),
            .I(\pid_alt.error_d_reg_prev_esr_RNICQF44Z0Z_13 ));
    CascadeMux I__2658 (
            .O(N__21090),
            .I(N__21087));
    InMux I__2657 (
            .O(N__21087),
            .I(N__21083));
    InMux I__2656 (
            .O(N__21086),
            .I(N__21080));
    LocalMux I__2655 (
            .O(N__21083),
            .I(N__21077));
    LocalMux I__2654 (
            .O(N__21080),
            .I(N__21074));
    Span4Mux_v I__2653 (
            .O(N__21077),
            .I(N__21071));
    Odrv4 I__2652 (
            .O(N__21074),
            .I(\pid_alt.error_d_reg_prev_esr_RNISAO32Z0Z_12 ));
    Odrv4 I__2651 (
            .O(N__21071),
            .I(\pid_alt.error_d_reg_prev_esr_RNISAO32Z0Z_12 ));
    InMux I__2650 (
            .O(N__21066),
            .I(\pid_alt.un1_pid_prereg_0_cry_13 ));
    InMux I__2649 (
            .O(N__21063),
            .I(N__21060));
    LocalMux I__2648 (
            .O(N__21060),
            .I(N__21057));
    Span4Mux_h I__2647 (
            .O(N__21057),
            .I(N__21054));
    Odrv4 I__2646 (
            .O(N__21054),
            .I(\pid_alt.error_d_reg_prev_esr_RNI88G14Z0Z_14 ));
    CascadeMux I__2645 (
            .O(N__21051),
            .I(N__21048));
    InMux I__2644 (
            .O(N__21048),
            .I(N__21044));
    CascadeMux I__2643 (
            .O(N__21047),
            .I(N__21041));
    LocalMux I__2642 (
            .O(N__21044),
            .I(N__21038));
    InMux I__2641 (
            .O(N__21041),
            .I(N__21035));
    Span4Mux_h I__2640 (
            .O(N__21038),
            .I(N__21032));
    LocalMux I__2639 (
            .O(N__21035),
            .I(\pid_alt.error_d_reg_prev_esr_RNIGFN02Z0Z_13 ));
    Odrv4 I__2638 (
            .O(N__21032),
            .I(\pid_alt.error_d_reg_prev_esr_RNIGFN02Z0Z_13 ));
    InMux I__2637 (
            .O(N__21027),
            .I(bfn_7_15_0_));
    InMux I__2636 (
            .O(N__21024),
            .I(N__21021));
    LocalMux I__2635 (
            .O(N__21021),
            .I(N__21018));
    Odrv4 I__2634 (
            .O(N__21018),
            .I(\pid_alt.error_d_reg_prev_esr_RNIOQI14Z0Z_15 ));
    CascadeMux I__2633 (
            .O(N__21015),
            .I(N__21012));
    InMux I__2632 (
            .O(N__21012),
            .I(N__21008));
    InMux I__2631 (
            .O(N__21011),
            .I(N__21005));
    LocalMux I__2630 (
            .O(N__21008),
            .I(N__21002));
    LocalMux I__2629 (
            .O(N__21005),
            .I(N__20999));
    Span4Mux_h I__2628 (
            .O(N__21002),
            .I(N__20996));
    Odrv4 I__2627 (
            .O(N__20999),
            .I(\pid_alt.error_d_reg_prev_esr_RNIOOO02Z0Z_14 ));
    Odrv4 I__2626 (
            .O(N__20996),
            .I(\pid_alt.error_d_reg_prev_esr_RNIOOO02Z0Z_14 ));
    InMux I__2625 (
            .O(N__20991),
            .I(N__20988));
    LocalMux I__2624 (
            .O(N__20988),
            .I(N__20985));
    Odrv4 I__2623 (
            .O(N__20985),
            .I(\pid_alt.pid_preregZ0Z_16 ));
    InMux I__2622 (
            .O(N__20982),
            .I(\pid_alt.un1_pid_prereg_0_cry_15 ));
    InMux I__2621 (
            .O(N__20979),
            .I(N__20976));
    LocalMux I__2620 (
            .O(N__20976),
            .I(N__20973));
    Odrv4 I__2619 (
            .O(N__20973),
            .I(\pid_alt.error_d_reg_prev_esr_RNI8DL14Z0Z_16 ));
    CascadeMux I__2618 (
            .O(N__20970),
            .I(N__20967));
    InMux I__2617 (
            .O(N__20967),
            .I(N__20963));
    InMux I__2616 (
            .O(N__20966),
            .I(N__20960));
    LocalMux I__2615 (
            .O(N__20963),
            .I(N__20957));
    LocalMux I__2614 (
            .O(N__20960),
            .I(\pid_alt.error_d_reg_prev_esr_RNI02Q02Z0Z_15 ));
    Odrv12 I__2613 (
            .O(N__20957),
            .I(\pid_alt.error_d_reg_prev_esr_RNI02Q02Z0Z_15 ));
    InMux I__2612 (
            .O(N__20952),
            .I(N__20949));
    LocalMux I__2611 (
            .O(N__20949),
            .I(N__20946));
    Odrv4 I__2610 (
            .O(N__20946),
            .I(\pid_alt.pid_preregZ0Z_17 ));
    InMux I__2609 (
            .O(N__20943),
            .I(\pid_alt.un1_pid_prereg_0_cry_16 ));
    InMux I__2608 (
            .O(N__20940),
            .I(N__20937));
    LocalMux I__2607 (
            .O(N__20937),
            .I(N__20934));
    Odrv12 I__2606 (
            .O(N__20934),
            .I(\pid_alt.error_d_reg_prev_esr_RNIOVN14Z0Z_17 ));
    CascadeMux I__2605 (
            .O(N__20931),
            .I(N__20927));
    CascadeMux I__2604 (
            .O(N__20930),
            .I(N__20924));
    InMux I__2603 (
            .O(N__20927),
            .I(N__20921));
    InMux I__2602 (
            .O(N__20924),
            .I(N__20918));
    LocalMux I__2601 (
            .O(N__20921),
            .I(N__20915));
    LocalMux I__2600 (
            .O(N__20918),
            .I(\pid_alt.error_d_reg_prev_esr_RNI8BR02Z0Z_16 ));
    Odrv4 I__2599 (
            .O(N__20915),
            .I(\pid_alt.error_d_reg_prev_esr_RNI8BR02Z0Z_16 ));
    InMux I__2598 (
            .O(N__20910),
            .I(N__20907));
    LocalMux I__2597 (
            .O(N__20907),
            .I(N__20904));
    Odrv4 I__2596 (
            .O(N__20904),
            .I(\pid_alt.pid_preregZ0Z_18 ));
    InMux I__2595 (
            .O(N__20901),
            .I(\pid_alt.un1_pid_prereg_0_cry_17 ));
    InMux I__2594 (
            .O(N__20898),
            .I(N__20895));
    LocalMux I__2593 (
            .O(N__20895),
            .I(N__20892));
    Odrv4 I__2592 (
            .O(N__20892),
            .I(\pid_alt.error_d_reg_prev_esr_RNI8IQ14Z0Z_18 ));
    CascadeMux I__2591 (
            .O(N__20889),
            .I(N__20885));
    CascadeMux I__2590 (
            .O(N__20888),
            .I(N__20882));
    InMux I__2589 (
            .O(N__20885),
            .I(N__20879));
    InMux I__2588 (
            .O(N__20882),
            .I(N__20876));
    LocalMux I__2587 (
            .O(N__20879),
            .I(N__20873));
    LocalMux I__2586 (
            .O(N__20876),
            .I(\pid_alt.error_d_reg_prev_esr_RNIGKS02Z0Z_17 ));
    Odrv4 I__2585 (
            .O(N__20873),
            .I(\pid_alt.error_d_reg_prev_esr_RNIGKS02Z0Z_17 ));
    CascadeMux I__2584 (
            .O(N__20868),
            .I(N__20865));
    InMux I__2583 (
            .O(N__20865),
            .I(N__20862));
    LocalMux I__2582 (
            .O(N__20862),
            .I(N__20859));
    Odrv4 I__2581 (
            .O(N__20859),
            .I(\pid_alt.pid_preregZ0Z_19 ));
    InMux I__2580 (
            .O(N__20856),
            .I(\pid_alt.un1_pid_prereg_0_cry_18 ));
    InMux I__2579 (
            .O(N__20853),
            .I(N__20850));
    LocalMux I__2578 (
            .O(N__20850),
            .I(N__20847));
    Odrv4 I__2577 (
            .O(N__20847),
            .I(\pid_alt.error_d_reg_prev_esr_RNILDG87Z0Z_2 ));
    InMux I__2576 (
            .O(N__20844),
            .I(\pid_alt.un1_pid_prereg_0_cry_2 ));
    InMux I__2575 (
            .O(N__20841),
            .I(\pid_alt.un1_pid_prereg_0_cry_3 ));
    InMux I__2574 (
            .O(N__20838),
            .I(\pid_alt.un1_pid_prereg_0_cry_4 ));
    InMux I__2573 (
            .O(N__20835),
            .I(\pid_alt.un1_pid_prereg_0_cry_5 ));
    InMux I__2572 (
            .O(N__20832),
            .I(bfn_7_14_0_));
    InMux I__2571 (
            .O(N__20829),
            .I(N__20826));
    LocalMux I__2570 (
            .O(N__20826),
            .I(N__20823));
    Span4Mux_h I__2569 (
            .O(N__20823),
            .I(N__20820));
    Odrv4 I__2568 (
            .O(N__20820),
            .I(\pid_alt.error_d_reg_prev_esr_RNI5G6Q5Z0Z_7 ));
    InMux I__2567 (
            .O(N__20817),
            .I(\pid_alt.un1_pid_prereg_0_cry_7 ));
    InMux I__2566 (
            .O(N__20814),
            .I(\pid_alt.un1_pid_prereg_0_cry_8 ));
    InMux I__2565 (
            .O(N__20811),
            .I(\pid_alt.un1_pid_prereg_0_cry_9 ));
    InMux I__2564 (
            .O(N__20808),
            .I(N__20805));
    LocalMux I__2563 (
            .O(N__20805),
            .I(N__20802));
    Odrv4 I__2562 (
            .O(N__20802),
            .I(\pid_alt.error_d_reg_prev_esr_RNIKQBI4Z0Z_10 ));
    InMux I__2561 (
            .O(N__20799),
            .I(\pid_alt.un1_pid_prereg_0_cry_10 ));
    InMux I__2560 (
            .O(N__20796),
            .I(N__20793));
    LocalMux I__2559 (
            .O(N__20793),
            .I(N__20790));
    Odrv12 I__2558 (
            .O(N__20790),
            .I(\pid_alt.error_d_reg_esr_RNITF511_2Z0Z_1 ));
    InMux I__2557 (
            .O(N__20787),
            .I(N__20784));
    LocalMux I__2556 (
            .O(N__20784),
            .I(N__20779));
    InMux I__2555 (
            .O(N__20783),
            .I(N__20774));
    InMux I__2554 (
            .O(N__20782),
            .I(N__20771));
    Span4Mux_h I__2553 (
            .O(N__20779),
            .I(N__20768));
    InMux I__2552 (
            .O(N__20778),
            .I(N__20765));
    InMux I__2551 (
            .O(N__20777),
            .I(N__20762));
    LocalMux I__2550 (
            .O(N__20774),
            .I(N__20757));
    LocalMux I__2549 (
            .O(N__20771),
            .I(N__20757));
    Span4Mux_h I__2548 (
            .O(N__20768),
            .I(N__20754));
    LocalMux I__2547 (
            .O(N__20765),
            .I(N__20749));
    LocalMux I__2546 (
            .O(N__20762),
            .I(N__20749));
    Span4Mux_h I__2545 (
            .O(N__20757),
            .I(N__20746));
    Odrv4 I__2544 (
            .O(N__20754),
            .I(\pid_alt.error_p_regZ0Z_0 ));
    Odrv4 I__2543 (
            .O(N__20749),
            .I(\pid_alt.error_p_regZ0Z_0 ));
    Odrv4 I__2542 (
            .O(N__20746),
            .I(\pid_alt.error_p_regZ0Z_0 ));
    InMux I__2541 (
            .O(N__20739),
            .I(N__20735));
    InMux I__2540 (
            .O(N__20738),
            .I(N__20731));
    LocalMux I__2539 (
            .O(N__20735),
            .I(N__20728));
    InMux I__2538 (
            .O(N__20734),
            .I(N__20725));
    LocalMux I__2537 (
            .O(N__20731),
            .I(N__20719));
    Span4Mux_v I__2536 (
            .O(N__20728),
            .I(N__20714));
    LocalMux I__2535 (
            .O(N__20725),
            .I(N__20714));
    InMux I__2534 (
            .O(N__20724),
            .I(N__20711));
    InMux I__2533 (
            .O(N__20723),
            .I(N__20708));
    InMux I__2532 (
            .O(N__20722),
            .I(N__20705));
    Span4Mux_h I__2531 (
            .O(N__20719),
            .I(N__20702));
    Span4Mux_v I__2530 (
            .O(N__20714),
            .I(N__20699));
    LocalMux I__2529 (
            .O(N__20711),
            .I(N__20694));
    LocalMux I__2528 (
            .O(N__20708),
            .I(N__20694));
    LocalMux I__2527 (
            .O(N__20705),
            .I(N__20691));
    Odrv4 I__2526 (
            .O(N__20702),
            .I(\pid_alt.error_d_regZ0Z_0 ));
    Odrv4 I__2525 (
            .O(N__20699),
            .I(\pid_alt.error_d_regZ0Z_0 ));
    Odrv4 I__2524 (
            .O(N__20694),
            .I(\pid_alt.error_d_regZ0Z_0 ));
    Odrv12 I__2523 (
            .O(N__20691),
            .I(\pid_alt.error_d_regZ0Z_0 ));
    InMux I__2522 (
            .O(N__20682),
            .I(N__20678));
    CascadeMux I__2521 (
            .O(N__20681),
            .I(N__20674));
    LocalMux I__2520 (
            .O(N__20678),
            .I(N__20671));
    InMux I__2519 (
            .O(N__20677),
            .I(N__20668));
    InMux I__2518 (
            .O(N__20674),
            .I(N__20665));
    Odrv4 I__2517 (
            .O(N__20671),
            .I(\dron_frame_decoder_1.stateZ0Z_1 ));
    LocalMux I__2516 (
            .O(N__20668),
            .I(\dron_frame_decoder_1.stateZ0Z_1 ));
    LocalMux I__2515 (
            .O(N__20665),
            .I(\dron_frame_decoder_1.stateZ0Z_1 ));
    InMux I__2514 (
            .O(N__20658),
            .I(N__20655));
    LocalMux I__2513 (
            .O(N__20655),
            .I(N__20652));
    Odrv4 I__2512 (
            .O(N__20652),
            .I(\dron_frame_decoder_1.state_RNO_1Z0Z_0 ));
    CascadeMux I__2511 (
            .O(N__20649),
            .I(N__20646));
    InMux I__2510 (
            .O(N__20646),
            .I(N__20643));
    LocalMux I__2509 (
            .O(N__20643),
            .I(N__20639));
    InMux I__2508 (
            .O(N__20642),
            .I(N__20636));
    Span4Mux_v I__2507 (
            .O(N__20639),
            .I(N__20631));
    LocalMux I__2506 (
            .O(N__20636),
            .I(N__20631));
    Span4Mux_h I__2505 (
            .O(N__20631),
            .I(N__20628));
    Span4Mux_v I__2504 (
            .O(N__20628),
            .I(N__20625));
    Odrv4 I__2503 (
            .O(N__20625),
            .I(\pid_alt.error_d_reg_prev_i_0 ));
    InMux I__2502 (
            .O(N__20622),
            .I(N__20619));
    LocalMux I__2501 (
            .O(N__20619),
            .I(N__20616));
    Span4Mux_h I__2500 (
            .O(N__20616),
            .I(N__20613));
    Odrv4 I__2499 (
            .O(N__20613),
            .I(\pid_alt.error_p_reg_esr_RNI3SMI1Z0Z_0 ));
    InMux I__2498 (
            .O(N__20610),
            .I(\pid_alt.un1_pid_prereg_un1_pid_prereg_0_cry_0_c_THRU_CO ));
    InMux I__2497 (
            .O(N__20607),
            .I(N__20604));
    LocalMux I__2496 (
            .O(N__20604),
            .I(\pid_alt.error_p_reg_esr_RNIFPN33Z0Z_0 ));
    InMux I__2495 (
            .O(N__20601),
            .I(\pid_alt.un1_pid_prereg_0_cry_0 ));
    InMux I__2494 (
            .O(N__20598),
            .I(N__20595));
    LocalMux I__2493 (
            .O(N__20595),
            .I(N__20592));
    Odrv12 I__2492 (
            .O(N__20592),
            .I(\pid_alt.error_d_reg_prev_esr_RNIF0465Z0Z_2 ));
    InMux I__2491 (
            .O(N__20589),
            .I(\pid_alt.un1_pid_prereg_0_cry_1 ));
    CascadeMux I__2490 (
            .O(N__20586),
            .I(\Commands_frame_decoder.source_CH2data_1_sqmuxa_cascade_ ));
    CascadeMux I__2489 (
            .O(N__20583),
            .I(\dron_frame_decoder_1.state_ns_0_i_a2_1_0Z0Z_3_cascade_ ));
    InMux I__2488 (
            .O(N__20580),
            .I(N__20577));
    LocalMux I__2487 (
            .O(N__20577),
            .I(\dron_frame_decoder_1.N_188_4 ));
    CascadeMux I__2486 (
            .O(N__20574),
            .I(\dron_frame_decoder_1.state_ns_0_i_a2_1Z0Z_3_cascade_ ));
    CascadeMux I__2485 (
            .O(N__20571),
            .I(\dron_frame_decoder_1.state_RNO_0Z0Z_0_cascade_ ));
    CascadeMux I__2484 (
            .O(N__20568),
            .I(\dron_frame_decoder_1.state_ns_0_i_a2_0_0_1Z0Z_1_cascade_ ));
    InMux I__2483 (
            .O(N__20565),
            .I(N__20562));
    LocalMux I__2482 (
            .O(N__20562),
            .I(\dron_frame_decoder_1.state_ns_0_i_a2_0_1 ));
    CascadeMux I__2481 (
            .O(N__20559),
            .I(N__20556));
    InMux I__2480 (
            .O(N__20556),
            .I(N__20552));
    InMux I__2479 (
            .O(N__20555),
            .I(N__20549));
    LocalMux I__2478 (
            .O(N__20552),
            .I(N__20546));
    LocalMux I__2477 (
            .O(N__20549),
            .I(\dron_frame_decoder_1.state_ns_0_i_a2_1Z0Z_3 ));
    Odrv4 I__2476 (
            .O(N__20546),
            .I(\dron_frame_decoder_1.state_ns_0_i_a2_1Z0Z_3 ));
    CascadeMux I__2475 (
            .O(N__20541),
            .I(\dron_frame_decoder_1.state_ns_0_i_a2_0_1_cascade_ ));
    InMux I__2474 (
            .O(N__20538),
            .I(\dron_frame_decoder_1.un1_WDT_cry_11 ));
    CascadeMux I__2473 (
            .O(N__20535),
            .I(N__20532));
    InMux I__2472 (
            .O(N__20532),
            .I(N__20528));
    CascadeMux I__2471 (
            .O(N__20531),
            .I(N__20524));
    LocalMux I__2470 (
            .O(N__20528),
            .I(N__20520));
    InMux I__2469 (
            .O(N__20527),
            .I(N__20515));
    InMux I__2468 (
            .O(N__20524),
            .I(N__20515));
    InMux I__2467 (
            .O(N__20523),
            .I(N__20512));
    Span4Mux_v I__2466 (
            .O(N__20520),
            .I(N__20507));
    LocalMux I__2465 (
            .O(N__20515),
            .I(N__20507));
    LocalMux I__2464 (
            .O(N__20512),
            .I(\dron_frame_decoder_1.WDTZ0Z_13 ));
    Odrv4 I__2463 (
            .O(N__20507),
            .I(\dron_frame_decoder_1.WDTZ0Z_13 ));
    InMux I__2462 (
            .O(N__20502),
            .I(\dron_frame_decoder_1.un1_WDT_cry_12 ));
    InMux I__2461 (
            .O(N__20499),
            .I(N__20496));
    LocalMux I__2460 (
            .O(N__20496),
            .I(N__20491));
    InMux I__2459 (
            .O(N__20495),
            .I(N__20488));
    InMux I__2458 (
            .O(N__20494),
            .I(N__20485));
    Span4Mux_v I__2457 (
            .O(N__20491),
            .I(N__20480));
    LocalMux I__2456 (
            .O(N__20488),
            .I(N__20480));
    LocalMux I__2455 (
            .O(N__20485),
            .I(\dron_frame_decoder_1.WDTZ0Z_14 ));
    Odrv4 I__2454 (
            .O(N__20480),
            .I(\dron_frame_decoder_1.WDTZ0Z_14 ));
    InMux I__2453 (
            .O(N__20475),
            .I(\dron_frame_decoder_1.un1_WDT_cry_13 ));
    InMux I__2452 (
            .O(N__20472),
            .I(\dron_frame_decoder_1.un1_WDT_cry_14 ));
    CascadeMux I__2451 (
            .O(N__20469),
            .I(N__20466));
    InMux I__2450 (
            .O(N__20466),
            .I(N__20462));
    InMux I__2449 (
            .O(N__20465),
            .I(N__20459));
    LocalMux I__2448 (
            .O(N__20462),
            .I(N__20455));
    LocalMux I__2447 (
            .O(N__20459),
            .I(N__20452));
    InMux I__2446 (
            .O(N__20458),
            .I(N__20449));
    Span4Mux_v I__2445 (
            .O(N__20455),
            .I(N__20444));
    Span4Mux_v I__2444 (
            .O(N__20452),
            .I(N__20444));
    LocalMux I__2443 (
            .O(N__20449),
            .I(\dron_frame_decoder_1.WDTZ0Z_15 ));
    Odrv4 I__2442 (
            .O(N__20444),
            .I(\dron_frame_decoder_1.WDTZ0Z_15 ));
    CascadeMux I__2441 (
            .O(N__20439),
            .I(N__20435));
    InMux I__2440 (
            .O(N__20438),
            .I(N__20430));
    InMux I__2439 (
            .O(N__20435),
            .I(N__20430));
    LocalMux I__2438 (
            .O(N__20430),
            .I(\dron_frame_decoder_1.stateZ0Z_3 ));
    CascadeMux I__2437 (
            .O(N__20427),
            .I(N__20424));
    InMux I__2436 (
            .O(N__20424),
            .I(N__20418));
    InMux I__2435 (
            .O(N__20423),
            .I(N__20418));
    LocalMux I__2434 (
            .O(N__20418),
            .I(\dron_frame_decoder_1.stateZ0Z_2 ));
    CascadeMux I__2433 (
            .O(N__20415),
            .I(\dron_frame_decoder_1.N_188_4_cascade_ ));
    InMux I__2432 (
            .O(N__20412),
            .I(N__20409));
    LocalMux I__2431 (
            .O(N__20409),
            .I(\dron_frame_decoder_1.state_ns_0_i_a2_0_0_3 ));
    InMux I__2430 (
            .O(N__20406),
            .I(N__20403));
    LocalMux I__2429 (
            .O(N__20403),
            .I(N__20399));
    InMux I__2428 (
            .O(N__20402),
            .I(N__20396));
    Span4Mux_v I__2427 (
            .O(N__20399),
            .I(N__20393));
    LocalMux I__2426 (
            .O(N__20396),
            .I(\dron_frame_decoder_1.WDTZ0Z_4 ));
    Odrv4 I__2425 (
            .O(N__20393),
            .I(\dron_frame_decoder_1.WDTZ0Z_4 ));
    InMux I__2424 (
            .O(N__20388),
            .I(\dron_frame_decoder_1.un1_WDT_cry_3 ));
    InMux I__2423 (
            .O(N__20385),
            .I(N__20382));
    LocalMux I__2422 (
            .O(N__20382),
            .I(N__20378));
    InMux I__2421 (
            .O(N__20381),
            .I(N__20375));
    Span4Mux_v I__2420 (
            .O(N__20378),
            .I(N__20372));
    LocalMux I__2419 (
            .O(N__20375),
            .I(\dron_frame_decoder_1.WDTZ0Z_5 ));
    Odrv4 I__2418 (
            .O(N__20372),
            .I(\dron_frame_decoder_1.WDTZ0Z_5 ));
    InMux I__2417 (
            .O(N__20367),
            .I(\dron_frame_decoder_1.un1_WDT_cry_4 ));
    InMux I__2416 (
            .O(N__20364),
            .I(N__20361));
    LocalMux I__2415 (
            .O(N__20361),
            .I(N__20357));
    InMux I__2414 (
            .O(N__20360),
            .I(N__20354));
    Span4Mux_h I__2413 (
            .O(N__20357),
            .I(N__20351));
    LocalMux I__2412 (
            .O(N__20354),
            .I(\dron_frame_decoder_1.WDTZ0Z_6 ));
    Odrv4 I__2411 (
            .O(N__20351),
            .I(\dron_frame_decoder_1.WDTZ0Z_6 ));
    InMux I__2410 (
            .O(N__20346),
            .I(\dron_frame_decoder_1.un1_WDT_cry_5 ));
    InMux I__2409 (
            .O(N__20343),
            .I(N__20340));
    LocalMux I__2408 (
            .O(N__20340),
            .I(N__20336));
    InMux I__2407 (
            .O(N__20339),
            .I(N__20333));
    Span4Mux_h I__2406 (
            .O(N__20336),
            .I(N__20330));
    LocalMux I__2405 (
            .O(N__20333),
            .I(\dron_frame_decoder_1.WDTZ0Z_7 ));
    Odrv4 I__2404 (
            .O(N__20330),
            .I(\dron_frame_decoder_1.WDTZ0Z_7 ));
    InMux I__2403 (
            .O(N__20325),
            .I(\dron_frame_decoder_1.un1_WDT_cry_6 ));
    InMux I__2402 (
            .O(N__20322),
            .I(N__20318));
    InMux I__2401 (
            .O(N__20321),
            .I(N__20315));
    LocalMux I__2400 (
            .O(N__20318),
            .I(N__20312));
    LocalMux I__2399 (
            .O(N__20315),
            .I(\dron_frame_decoder_1.WDTZ0Z_8 ));
    Odrv4 I__2398 (
            .O(N__20312),
            .I(\dron_frame_decoder_1.WDTZ0Z_8 ));
    InMux I__2397 (
            .O(N__20307),
            .I(bfn_7_8_0_));
    CascadeMux I__2396 (
            .O(N__20304),
            .I(N__20301));
    InMux I__2395 (
            .O(N__20301),
            .I(N__20297));
    InMux I__2394 (
            .O(N__20300),
            .I(N__20294));
    LocalMux I__2393 (
            .O(N__20297),
            .I(N__20291));
    LocalMux I__2392 (
            .O(N__20294),
            .I(\dron_frame_decoder_1.WDTZ0Z_9 ));
    Odrv4 I__2391 (
            .O(N__20291),
            .I(\dron_frame_decoder_1.WDTZ0Z_9 ));
    InMux I__2390 (
            .O(N__20286),
            .I(\dron_frame_decoder_1.un1_WDT_cry_8 ));
    InMux I__2389 (
            .O(N__20283),
            .I(N__20279));
    InMux I__2388 (
            .O(N__20282),
            .I(N__20276));
    LocalMux I__2387 (
            .O(N__20279),
            .I(N__20273));
    LocalMux I__2386 (
            .O(N__20276),
            .I(\dron_frame_decoder_1.WDTZ0Z_10 ));
    Odrv4 I__2385 (
            .O(N__20273),
            .I(\dron_frame_decoder_1.WDTZ0Z_10 ));
    InMux I__2384 (
            .O(N__20268),
            .I(\dron_frame_decoder_1.un1_WDT_cry_9 ));
    InMux I__2383 (
            .O(N__20265),
            .I(N__20258));
    InMux I__2382 (
            .O(N__20264),
            .I(N__20258));
    InMux I__2381 (
            .O(N__20263),
            .I(N__20255));
    LocalMux I__2380 (
            .O(N__20258),
            .I(N__20252));
    LocalMux I__2379 (
            .O(N__20255),
            .I(\dron_frame_decoder_1.WDTZ0Z_11 ));
    Odrv4 I__2378 (
            .O(N__20252),
            .I(\dron_frame_decoder_1.WDTZ0Z_11 ));
    InMux I__2377 (
            .O(N__20247),
            .I(\dron_frame_decoder_1.un1_WDT_cry_10 ));
    InMux I__2376 (
            .O(N__20244),
            .I(N__20237));
    InMux I__2375 (
            .O(N__20243),
            .I(N__20237));
    InMux I__2374 (
            .O(N__20242),
            .I(N__20234));
    LocalMux I__2373 (
            .O(N__20237),
            .I(N__20231));
    LocalMux I__2372 (
            .O(N__20234),
            .I(\dron_frame_decoder_1.WDTZ0Z_12 ));
    Odrv4 I__2371 (
            .O(N__20231),
            .I(\dron_frame_decoder_1.WDTZ0Z_12 ));
    InMux I__2370 (
            .O(N__20226),
            .I(N__20223));
    LocalMux I__2369 (
            .O(N__20223),
            .I(\pid_alt.error_d_reg_prev_esr_RNIKKKMZ0Z_22 ));
    InMux I__2368 (
            .O(N__20220),
            .I(N__20217));
    LocalMux I__2367 (
            .O(N__20217),
            .I(\pid_alt.error_d_reg_prev_esr_RNIMMKM_0Z0Z_23 ));
    CascadeMux I__2366 (
            .O(N__20214),
            .I(\pid_alt.error_d_reg_prev_esr_RNIKKKMZ0Z_22_cascade_ ));
    InMux I__2365 (
            .O(N__20211),
            .I(N__20208));
    LocalMux I__2364 (
            .O(N__20208),
            .I(N__20203));
    InMux I__2363 (
            .O(N__20207),
            .I(N__20198));
    InMux I__2362 (
            .O(N__20206),
            .I(N__20198));
    Span12Mux_s5_h I__2361 (
            .O(N__20203),
            .I(N__20193));
    LocalMux I__2360 (
            .O(N__20198),
            .I(N__20193));
    Span12Mux_v I__2359 (
            .O(N__20193),
            .I(N__20190));
    Odrv12 I__2358 (
            .O(N__20190),
            .I(\pid_alt.error_d_regZ0Z_23 ));
    InMux I__2357 (
            .O(N__20187),
            .I(N__20183));
    InMux I__2356 (
            .O(N__20186),
            .I(N__20180));
    LocalMux I__2355 (
            .O(N__20183),
            .I(\pid_alt.error_d_reg_prevZ0Z_23 ));
    LocalMux I__2354 (
            .O(N__20180),
            .I(\pid_alt.error_d_reg_prevZ0Z_23 ));
    InMux I__2353 (
            .O(N__20175),
            .I(N__20172));
    LocalMux I__2352 (
            .O(N__20172),
            .I(N__20169));
    Span4Mux_v I__2351 (
            .O(N__20169),
            .I(N__20166));
    Span4Mux_h I__2350 (
            .O(N__20166),
            .I(N__20163));
    Odrv4 I__2349 (
            .O(N__20163),
            .I(\pid_alt.O_1_8 ));
    CascadeMux I__2348 (
            .O(N__20160),
            .I(N__20156));
    InMux I__2347 (
            .O(N__20159),
            .I(N__20153));
    InMux I__2346 (
            .O(N__20156),
            .I(N__20150));
    LocalMux I__2345 (
            .O(N__20153),
            .I(N__20145));
    LocalMux I__2344 (
            .O(N__20150),
            .I(N__20145));
    Span4Mux_h I__2343 (
            .O(N__20145),
            .I(N__20142));
    Odrv4 I__2342 (
            .O(N__20142),
            .I(\dron_frame_decoder_1.WDT10_0_i ));
    InMux I__2341 (
            .O(N__20139),
            .I(N__20136));
    LocalMux I__2340 (
            .O(N__20136),
            .I(\dron_frame_decoder_1.WDTZ0Z_0 ));
    InMux I__2339 (
            .O(N__20133),
            .I(N__20130));
    LocalMux I__2338 (
            .O(N__20130),
            .I(\dron_frame_decoder_1.WDTZ0Z_1 ));
    InMux I__2337 (
            .O(N__20127),
            .I(\dron_frame_decoder_1.un1_WDT_cry_0 ));
    InMux I__2336 (
            .O(N__20124),
            .I(N__20121));
    LocalMux I__2335 (
            .O(N__20121),
            .I(\dron_frame_decoder_1.WDTZ0Z_2 ));
    InMux I__2334 (
            .O(N__20118),
            .I(\dron_frame_decoder_1.un1_WDT_cry_1 ));
    InMux I__2333 (
            .O(N__20115),
            .I(N__20112));
    LocalMux I__2332 (
            .O(N__20112),
            .I(\dron_frame_decoder_1.WDTZ0Z_3 ));
    InMux I__2331 (
            .O(N__20109),
            .I(\dron_frame_decoder_1.un1_WDT_cry_2 ));
    CascadeMux I__2330 (
            .O(N__20106),
            .I(\pid_alt.error_d_reg_prev_esr_RNISPHM_0Z0Z_15_cascade_ ));
    InMux I__2329 (
            .O(N__20103),
            .I(N__20097));
    InMux I__2328 (
            .O(N__20102),
            .I(N__20097));
    LocalMux I__2327 (
            .O(N__20097),
            .I(\pid_alt.error_d_reg_prev_esr_RNIPMHMZ0Z_14 ));
    InMux I__2326 (
            .O(N__20094),
            .I(N__20088));
    InMux I__2325 (
            .O(N__20093),
            .I(N__20088));
    LocalMux I__2324 (
            .O(N__20088),
            .I(N__20085));
    Span4Mux_h I__2323 (
            .O(N__20085),
            .I(N__20082));
    Span4Mux_v I__2322 (
            .O(N__20082),
            .I(N__20079));
    Odrv4 I__2321 (
            .O(N__20079),
            .I(\pid_alt.error_p_regZ0Z_14 ));
    CascadeMux I__2320 (
            .O(N__20076),
            .I(\pid_alt.error_d_reg_prev_esr_RNIPMHM_0Z0Z_14_cascade_ ));
    InMux I__2319 (
            .O(N__20073),
            .I(N__20064));
    InMux I__2318 (
            .O(N__20072),
            .I(N__20064));
    InMux I__2317 (
            .O(N__20071),
            .I(N__20064));
    LocalMux I__2316 (
            .O(N__20064),
            .I(N__20061));
    Span12Mux_s6_h I__2315 (
            .O(N__20061),
            .I(N__20058));
    Span12Mux_v I__2314 (
            .O(N__20058),
            .I(N__20055));
    Odrv12 I__2313 (
            .O(N__20055),
            .I(\pid_alt.error_d_regZ0Z_14 ));
    CascadeMux I__2312 (
            .O(N__20052),
            .I(N__20049));
    InMux I__2311 (
            .O(N__20049),
            .I(N__20043));
    InMux I__2310 (
            .O(N__20048),
            .I(N__20043));
    LocalMux I__2309 (
            .O(N__20043),
            .I(\pid_alt.error_d_reg_prevZ0Z_14 ));
    InMux I__2308 (
            .O(N__20040),
            .I(N__20034));
    InMux I__2307 (
            .O(N__20039),
            .I(N__20034));
    LocalMux I__2306 (
            .O(N__20034),
            .I(N__20031));
    Span4Mux_h I__2305 (
            .O(N__20031),
            .I(N__20028));
    Odrv4 I__2304 (
            .O(N__20028),
            .I(\pid_alt.error_d_reg_prev_esr_RNIMJHMZ0Z_13 ));
    InMux I__2303 (
            .O(N__20025),
            .I(N__20022));
    LocalMux I__2302 (
            .O(N__20022),
            .I(\pid_alt.error_d_reg_prev_esr_RNIPMHM_0Z0Z_14 ));
    CascadeMux I__2301 (
            .O(N__20019),
            .I(\pid_alt.error_d_reg_prev_esr_RNIMMKM_0Z0Z_23_cascade_ ));
    InMux I__2300 (
            .O(N__20016),
            .I(N__20012));
    InMux I__2299 (
            .O(N__20015),
            .I(N__20009));
    LocalMux I__2298 (
            .O(N__20012),
            .I(\pid_alt.error_d_reg_prevZ0Z_22 ));
    LocalMux I__2297 (
            .O(N__20009),
            .I(\pid_alt.error_d_reg_prevZ0Z_22 ));
    InMux I__2296 (
            .O(N__20004),
            .I(N__19998));
    InMux I__2295 (
            .O(N__20003),
            .I(N__19998));
    LocalMux I__2294 (
            .O(N__19998),
            .I(N__19994));
    InMux I__2293 (
            .O(N__19997),
            .I(N__19991));
    Span4Mux_v I__2292 (
            .O(N__19994),
            .I(N__19986));
    LocalMux I__2291 (
            .O(N__19991),
            .I(N__19986));
    Span4Mux_h I__2290 (
            .O(N__19986),
            .I(N__19983));
    Span4Mux_v I__2289 (
            .O(N__19983),
            .I(N__19980));
    Span4Mux_v I__2288 (
            .O(N__19980),
            .I(N__19977));
    Odrv4 I__2287 (
            .O(N__19977),
            .I(\pid_alt.error_d_regZ0Z_22 ));
    InMux I__2286 (
            .O(N__19974),
            .I(N__19968));
    InMux I__2285 (
            .O(N__19973),
            .I(N__19968));
    LocalMux I__2284 (
            .O(N__19968),
            .I(N__19965));
    Span4Mux_h I__2283 (
            .O(N__19965),
            .I(N__19962));
    Odrv4 I__2282 (
            .O(N__19962),
            .I(\pid_alt.error_p_regZ0Z_7 ));
    InMux I__2281 (
            .O(N__19959),
            .I(N__19953));
    InMux I__2280 (
            .O(N__19958),
            .I(N__19953));
    LocalMux I__2279 (
            .O(N__19953),
            .I(\pid_alt.error_d_reg_prevZ0Z_7 ));
    InMux I__2278 (
            .O(N__19950),
            .I(N__19941));
    InMux I__2277 (
            .O(N__19949),
            .I(N__19941));
    InMux I__2276 (
            .O(N__19948),
            .I(N__19941));
    LocalMux I__2275 (
            .O(N__19941),
            .I(N__19938));
    Span4Mux_v I__2274 (
            .O(N__19938),
            .I(N__19935));
    Span4Mux_h I__2273 (
            .O(N__19935),
            .I(N__19932));
    Odrv4 I__2272 (
            .O(N__19932),
            .I(\pid_alt.error_d_regZ0Z_7 ));
    InMux I__2271 (
            .O(N__19929),
            .I(N__19925));
    InMux I__2270 (
            .O(N__19928),
            .I(N__19922));
    LocalMux I__2269 (
            .O(N__19925),
            .I(N__19919));
    LocalMux I__2268 (
            .O(N__19922),
            .I(N__19916));
    Span4Mux_v I__2267 (
            .O(N__19919),
            .I(N__19913));
    Span4Mux_h I__2266 (
            .O(N__19916),
            .I(N__19910));
    Odrv4 I__2265 (
            .O(N__19913),
            .I(\pid_alt.error_p_regZ0Z_8 ));
    Odrv4 I__2264 (
            .O(N__19910),
            .I(\pid_alt.error_p_regZ0Z_8 ));
    InMux I__2263 (
            .O(N__19905),
            .I(N__19898));
    InMux I__2262 (
            .O(N__19904),
            .I(N__19898));
    InMux I__2261 (
            .O(N__19903),
            .I(N__19895));
    LocalMux I__2260 (
            .O(N__19898),
            .I(N__19890));
    LocalMux I__2259 (
            .O(N__19895),
            .I(N__19890));
    Span4Mux_v I__2258 (
            .O(N__19890),
            .I(N__19887));
    Span4Mux_h I__2257 (
            .O(N__19887),
            .I(N__19884));
    Odrv4 I__2256 (
            .O(N__19884),
            .I(\pid_alt.error_d_regZ0Z_8 ));
    InMux I__2255 (
            .O(N__19881),
            .I(N__19877));
    InMux I__2254 (
            .O(N__19880),
            .I(N__19874));
    LocalMux I__2253 (
            .O(N__19877),
            .I(\pid_alt.error_d_reg_prevZ0Z_8 ));
    LocalMux I__2252 (
            .O(N__19874),
            .I(\pid_alt.error_d_reg_prevZ0Z_8 ));
    InMux I__2251 (
            .O(N__19869),
            .I(N__19863));
    InMux I__2250 (
            .O(N__19868),
            .I(N__19863));
    LocalMux I__2249 (
            .O(N__19863),
            .I(N__19860));
    Odrv4 I__2248 (
            .O(N__19860),
            .I(\pid_alt.error_d_reg_prev_esr_RNISPHMZ0Z_15 ));
    InMux I__2247 (
            .O(N__19857),
            .I(N__19854));
    LocalMux I__2246 (
            .O(N__19854),
            .I(\pid_alt.error_d_reg_prevZ0Z_0 ));
    InMux I__2245 (
            .O(N__19851),
            .I(N__19847));
    InMux I__2244 (
            .O(N__19850),
            .I(N__19844));
    LocalMux I__2243 (
            .O(N__19847),
            .I(\pid_alt.error_d_reg_prevZ0Z_15 ));
    LocalMux I__2242 (
            .O(N__19844),
            .I(\pid_alt.error_d_reg_prevZ0Z_15 ));
    InMux I__2241 (
            .O(N__19839),
            .I(N__19835));
    InMux I__2240 (
            .O(N__19838),
            .I(N__19832));
    LocalMux I__2239 (
            .O(N__19835),
            .I(N__19827));
    LocalMux I__2238 (
            .O(N__19832),
            .I(N__19827));
    Span4Mux_v I__2237 (
            .O(N__19827),
            .I(N__19824));
    Span4Mux_h I__2236 (
            .O(N__19824),
            .I(N__19821));
    Odrv4 I__2235 (
            .O(N__19821),
            .I(\pid_alt.error_p_regZ0Z_15 ));
    InMux I__2234 (
            .O(N__19818),
            .I(N__19813));
    InMux I__2233 (
            .O(N__19817),
            .I(N__19810));
    InMux I__2232 (
            .O(N__19816),
            .I(N__19807));
    LocalMux I__2231 (
            .O(N__19813),
            .I(N__19800));
    LocalMux I__2230 (
            .O(N__19810),
            .I(N__19800));
    LocalMux I__2229 (
            .O(N__19807),
            .I(N__19800));
    Span12Mux_v I__2228 (
            .O(N__19800),
            .I(N__19797));
    Odrv12 I__2227 (
            .O(N__19797),
            .I(\pid_alt.error_d_regZ0Z_15 ));
    InMux I__2226 (
            .O(N__19794),
            .I(N__19791));
    LocalMux I__2225 (
            .O(N__19791),
            .I(\pid_alt.error_d_reg_prev_esr_RNISPHM_0Z0Z_15 ));
    CascadeMux I__2224 (
            .O(N__19788),
            .I(\pid_alt.error_d_reg_prev_esr_RNIVSHMZ0Z_16_cascade_ ));
    InMux I__2223 (
            .O(N__19785),
            .I(N__19779));
    InMux I__2222 (
            .O(N__19784),
            .I(N__19779));
    LocalMux I__2221 (
            .O(N__19779),
            .I(N__19776));
    Span4Mux_h I__2220 (
            .O(N__19776),
            .I(N__19773));
    Span4Mux_v I__2219 (
            .O(N__19773),
            .I(N__19770));
    Odrv4 I__2218 (
            .O(N__19770),
            .I(\pid_alt.error_p_regZ0Z_16 ));
    CascadeMux I__2217 (
            .O(N__19767),
            .I(N__19764));
    InMux I__2216 (
            .O(N__19764),
            .I(N__19758));
    InMux I__2215 (
            .O(N__19763),
            .I(N__19758));
    LocalMux I__2214 (
            .O(N__19758),
            .I(\pid_alt.error_d_reg_prevZ0Z_16 ));
    InMux I__2213 (
            .O(N__19755),
            .I(N__19746));
    InMux I__2212 (
            .O(N__19754),
            .I(N__19746));
    InMux I__2211 (
            .O(N__19753),
            .I(N__19746));
    LocalMux I__2210 (
            .O(N__19746),
            .I(N__19743));
    Span4Mux_v I__2209 (
            .O(N__19743),
            .I(N__19740));
    Span4Mux_v I__2208 (
            .O(N__19740),
            .I(N__19737));
    Span4Mux_h I__2207 (
            .O(N__19737),
            .I(N__19734));
    Odrv4 I__2206 (
            .O(N__19734),
            .I(\pid_alt.error_d_regZ0Z_16 ));
    InMux I__2205 (
            .O(N__19731),
            .I(N__19728));
    LocalMux I__2204 (
            .O(N__19728),
            .I(\pid_alt.error_d_reg_prev_esr_RNIVSHM_0Z0Z_16 ));
    CascadeMux I__2203 (
            .O(N__19725),
            .I(\pid_alt.error_d_reg_prev_esr_RNIVSHM_0Z0Z_16_cascade_ ));
    CascadeMux I__2202 (
            .O(N__19722),
            .I(\pid_alt.error_d_reg_prev_esr_RNII5611_0Z0Z_8_cascade_ ));
    InMux I__2201 (
            .O(N__19719),
            .I(N__19716));
    LocalMux I__2200 (
            .O(N__19716),
            .I(\pid_alt.error_d_reg_prev_esr_RNIF2611Z0Z_7 ));
    InMux I__2199 (
            .O(N__19713),
            .I(N__19710));
    LocalMux I__2198 (
            .O(N__19710),
            .I(\pid_alt.error_d_reg_prev_esr_RNII5611_0Z0Z_8 ));
    CascadeMux I__2197 (
            .O(N__19707),
            .I(\pid_alt.error_d_reg_prev_esr_RNIF2611Z0Z_7_cascade_ ));
    InMux I__2196 (
            .O(N__19704),
            .I(N__19698));
    InMux I__2195 (
            .O(N__19703),
            .I(N__19698));
    LocalMux I__2194 (
            .O(N__19698),
            .I(N__19695));
    Span4Mux_h I__2193 (
            .O(N__19695),
            .I(N__19692));
    Span4Mux_v I__2192 (
            .O(N__19692),
            .I(N__19689));
    Odrv4 I__2191 (
            .O(N__19689),
            .I(\pid_alt.error_p_regZ0Z_11 ));
    CascadeMux I__2190 (
            .O(N__19686),
            .I(N__19683));
    InMux I__2189 (
            .O(N__19683),
            .I(N__19677));
    InMux I__2188 (
            .O(N__19682),
            .I(N__19677));
    LocalMux I__2187 (
            .O(N__19677),
            .I(\pid_alt.error_d_reg_prevZ0Z_11 ));
    InMux I__2186 (
            .O(N__19674),
            .I(N__19665));
    InMux I__2185 (
            .O(N__19673),
            .I(N__19665));
    InMux I__2184 (
            .O(N__19672),
            .I(N__19665));
    LocalMux I__2183 (
            .O(N__19665),
            .I(N__19661));
    CascadeMux I__2182 (
            .O(N__19664),
            .I(N__19658));
    Span4Mux_v I__2181 (
            .O(N__19661),
            .I(N__19655));
    InMux I__2180 (
            .O(N__19658),
            .I(N__19652));
    Span4Mux_h I__2179 (
            .O(N__19655),
            .I(N__19649));
    LocalMux I__2178 (
            .O(N__19652),
            .I(\pid_alt.error_d_regZ0Z_11 ));
    Odrv4 I__2177 (
            .O(N__19649),
            .I(\pid_alt.error_d_regZ0Z_11 ));
    InMux I__2176 (
            .O(N__19644),
            .I(N__19641));
    LocalMux I__2175 (
            .O(N__19641),
            .I(\pid_alt.error_d_reg_prev_esr_RNI7E8R_0Z0Z_11 ));
    InMux I__2174 (
            .O(N__19638),
            .I(N__19632));
    InMux I__2173 (
            .O(N__19637),
            .I(N__19632));
    LocalMux I__2172 (
            .O(N__19632),
            .I(\pid_alt.error_d_reg_prev_esr_RNIDAHMZ0Z_10 ));
    CascadeMux I__2171 (
            .O(N__19629),
            .I(\pid_alt.error_d_reg_prev_esr_RNI7E8R_0Z0Z_11_cascade_ ));
    InMux I__2170 (
            .O(N__19626),
            .I(N__19623));
    LocalMux I__2169 (
            .O(N__19623),
            .I(N__19620));
    Odrv4 I__2168 (
            .O(N__19620),
            .I(\pid_alt.error_d_reg_prev_esr_RNIJGHM_0Z0Z_12 ));
    InMux I__2167 (
            .O(N__19617),
            .I(N__19614));
    LocalMux I__2166 (
            .O(N__19614),
            .I(N__19610));
    InMux I__2165 (
            .O(N__19613),
            .I(N__19607));
    Odrv4 I__2164 (
            .O(N__19610),
            .I(\pid_alt.error_d_reg_prev_esr_RNI7E8RZ0Z_11 ));
    LocalMux I__2163 (
            .O(N__19607),
            .I(\pid_alt.error_d_reg_prev_esr_RNI7E8RZ0Z_11 ));
    CascadeMux I__2162 (
            .O(N__19602),
            .I(\pid_alt.error_d_reg_prev_esr_RNIOFGB2Z0Z_10_cascade_ ));
    InMux I__2161 (
            .O(N__19599),
            .I(N__19596));
    LocalMux I__2160 (
            .O(N__19596),
            .I(\pid_alt.error_d_reg_prev_esr_RNIVSHMZ0Z_16 ));
    InMux I__2159 (
            .O(N__19593),
            .I(N__19587));
    InMux I__2158 (
            .O(N__19592),
            .I(N__19587));
    LocalMux I__2157 (
            .O(N__19587),
            .I(N__19584));
    Span12Mux_h I__2156 (
            .O(N__19584),
            .I(N__19581));
    Odrv12 I__2155 (
            .O(N__19581),
            .I(\pid_alt.error_d_reg_prev_esr_RNI20IM_0Z0Z_17 ));
    CascadeMux I__2154 (
            .O(N__19578),
            .I(\dron_frame_decoder_1.WDT10lto9_3_cascade_ ));
    CascadeMux I__2153 (
            .O(N__19575),
            .I(\dron_frame_decoder_1.WDT10lt12_0_cascade_ ));
    InMux I__2152 (
            .O(N__19572),
            .I(N__19569));
    LocalMux I__2151 (
            .O(N__19569),
            .I(\dron_frame_decoder_1.WDT10_0_i_1 ));
    InMux I__2150 (
            .O(N__19566),
            .I(N__19563));
    LocalMux I__2149 (
            .O(N__19563),
            .I(\dron_frame_decoder_1.WDT10lt12_0 ));
    InMux I__2148 (
            .O(N__19560),
            .I(N__19557));
    LocalMux I__2147 (
            .O(N__19557),
            .I(\dron_frame_decoder_1.WDT10lt14_0 ));
    CEMux I__2146 (
            .O(N__19554),
            .I(N__19551));
    LocalMux I__2145 (
            .O(N__19551),
            .I(\pid_alt.state_1_0_0 ));
    InMux I__2144 (
            .O(N__19548),
            .I(N__19542));
    InMux I__2143 (
            .O(N__19547),
            .I(N__19542));
    LocalMux I__2142 (
            .O(N__19542),
            .I(N__19539));
    Span4Mux_v I__2141 (
            .O(N__19539),
            .I(N__19536));
    Odrv4 I__2140 (
            .O(N__19536),
            .I(\pid_alt.error_p_regZ0Z_12 ));
    InMux I__2139 (
            .O(N__19533),
            .I(N__19527));
    InMux I__2138 (
            .O(N__19532),
            .I(N__19527));
    LocalMux I__2137 (
            .O(N__19527),
            .I(\pid_alt.error_d_reg_prevZ0Z_12 ));
    InMux I__2136 (
            .O(N__19524),
            .I(N__19515));
    InMux I__2135 (
            .O(N__19523),
            .I(N__19515));
    InMux I__2134 (
            .O(N__19522),
            .I(N__19515));
    LocalMux I__2133 (
            .O(N__19515),
            .I(N__19512));
    Span4Mux_h I__2132 (
            .O(N__19512),
            .I(N__19509));
    Sp12to4 I__2131 (
            .O(N__19509),
            .I(N__19506));
    Odrv12 I__2130 (
            .O(N__19506),
            .I(\pid_alt.error_d_regZ0Z_12 ));
    CascadeMux I__2129 (
            .O(N__19503),
            .I(\pid_alt.error_d_reg_prev_esr_RNIJGHM_0Z0Z_12_cascade_ ));
    InMux I__2128 (
            .O(N__19500),
            .I(N__19495));
    InMux I__2127 (
            .O(N__19499),
            .I(N__19490));
    InMux I__2126 (
            .O(N__19498),
            .I(N__19490));
    LocalMux I__2125 (
            .O(N__19495),
            .I(N__19485));
    LocalMux I__2124 (
            .O(N__19490),
            .I(N__19485));
    Span4Mux_h I__2123 (
            .O(N__19485),
            .I(N__19482));
    Sp12to4 I__2122 (
            .O(N__19482),
            .I(N__19479));
    Odrv12 I__2121 (
            .O(N__19479),
            .I(\pid_alt.error_d_regZ0Z_13 ));
    InMux I__2120 (
            .O(N__19476),
            .I(N__19472));
    InMux I__2119 (
            .O(N__19475),
            .I(N__19469));
    LocalMux I__2118 (
            .O(N__19472),
            .I(\pid_alt.error_d_reg_prevZ0Z_13 ));
    LocalMux I__2117 (
            .O(N__19469),
            .I(\pid_alt.error_d_reg_prevZ0Z_13 ));
    InMux I__2116 (
            .O(N__19464),
            .I(N__19461));
    LocalMux I__2115 (
            .O(N__19461),
            .I(N__19458));
    Span4Mux_h I__2114 (
            .O(N__19458),
            .I(N__19455));
    Odrv4 I__2113 (
            .O(N__19455),
            .I(\pid_alt.O_0_15 ));
    InMux I__2112 (
            .O(N__19452),
            .I(N__19446));
    InMux I__2111 (
            .O(N__19451),
            .I(N__19446));
    LocalMux I__2110 (
            .O(N__19446),
            .I(N__19443));
    Span4Mux_h I__2109 (
            .O(N__19443),
            .I(N__19440));
    Span4Mux_v I__2108 (
            .O(N__19440),
            .I(N__19437));
    Odrv4 I__2107 (
            .O(N__19437),
            .I(\pid_alt.error_p_regZ0Z_18 ));
    CascadeMux I__2106 (
            .O(N__19434),
            .I(\pid_alt.error_d_reg_prev_esr_RNI53IM_0Z0Z_18_cascade_ ));
    InMux I__2105 (
            .O(N__19431),
            .I(N__19422));
    InMux I__2104 (
            .O(N__19430),
            .I(N__19422));
    InMux I__2103 (
            .O(N__19429),
            .I(N__19422));
    LocalMux I__2102 (
            .O(N__19422),
            .I(N__19419));
    Span4Mux_v I__2101 (
            .O(N__19419),
            .I(N__19416));
    Span4Mux_h I__2100 (
            .O(N__19416),
            .I(N__19413));
    Span4Mux_v I__2099 (
            .O(N__19413),
            .I(N__19410));
    Odrv4 I__2098 (
            .O(N__19410),
            .I(\pid_alt.error_d_regZ0Z_18 ));
    CascadeMux I__2097 (
            .O(N__19407),
            .I(N__19404));
    InMux I__2096 (
            .O(N__19404),
            .I(N__19398));
    InMux I__2095 (
            .O(N__19403),
            .I(N__19398));
    LocalMux I__2094 (
            .O(N__19398),
            .I(\pid_alt.error_d_reg_prevZ0Z_18 ));
    InMux I__2093 (
            .O(N__19395),
            .I(N__19392));
    LocalMux I__2092 (
            .O(N__19392),
            .I(\pid_alt.error_d_reg_prev_esr_RNI53IM_0Z0Z_18 ));
    InMux I__2091 (
            .O(N__19389),
            .I(N__19383));
    InMux I__2090 (
            .O(N__19388),
            .I(N__19383));
    LocalMux I__2089 (
            .O(N__19383),
            .I(N__19380));
    Span4Mux_h I__2088 (
            .O(N__19380),
            .I(N__19377));
    Span4Mux_v I__2087 (
            .O(N__19377),
            .I(N__19374));
    Odrv4 I__2086 (
            .O(N__19374),
            .I(\pid_alt.error_d_reg_prev_esr_RNI20IMZ0Z_17 ));
    InMux I__2085 (
            .O(N__19371),
            .I(N__19367));
    InMux I__2084 (
            .O(N__19370),
            .I(N__19364));
    LocalMux I__2083 (
            .O(N__19367),
            .I(N__19359));
    LocalMux I__2082 (
            .O(N__19364),
            .I(N__19359));
    Span4Mux_h I__2081 (
            .O(N__19359),
            .I(N__19356));
    Span4Mux_v I__2080 (
            .O(N__19356),
            .I(N__19353));
    Odrv4 I__2079 (
            .O(N__19353),
            .I(\pid_alt.error_p_regZ0Z_13 ));
    CascadeMux I__2078 (
            .O(N__19350),
            .I(\pid_alt.error_d_reg_prev_esr_RNIMJHM_0Z0Z_13_cascade_ ));
    InMux I__2077 (
            .O(N__19347),
            .I(N__19344));
    LocalMux I__2076 (
            .O(N__19344),
            .I(\pid_alt.error_d_reg_prev_esr_RNIJGHMZ0Z_12 ));
    InMux I__2075 (
            .O(N__19341),
            .I(N__19338));
    LocalMux I__2074 (
            .O(N__19338),
            .I(\pid_alt.error_d_reg_prev_esr_RNIMJHM_0Z0Z_13 ));
    CascadeMux I__2073 (
            .O(N__19335),
            .I(\pid_alt.error_d_reg_prev_esr_RNIJGHMZ0Z_12_cascade_ ));
    InMux I__2072 (
            .O(N__19332),
            .I(N__19329));
    LocalMux I__2071 (
            .O(N__19329),
            .I(\pid_alt.g0_4_0 ));
    InMux I__2070 (
            .O(N__19326),
            .I(N__19321));
    InMux I__2069 (
            .O(N__19325),
            .I(N__19318));
    CascadeMux I__2068 (
            .O(N__19324),
            .I(N__19314));
    LocalMux I__2067 (
            .O(N__19321),
            .I(N__19308));
    LocalMux I__2066 (
            .O(N__19318),
            .I(N__19308));
    InMux I__2065 (
            .O(N__19317),
            .I(N__19305));
    InMux I__2064 (
            .O(N__19314),
            .I(N__19300));
    InMux I__2063 (
            .O(N__19313),
            .I(N__19300));
    Odrv4 I__2062 (
            .O(N__19308),
            .I(\pid_alt.error_d_reg_prevZ0Z_2 ));
    LocalMux I__2061 (
            .O(N__19305),
            .I(\pid_alt.error_d_reg_prevZ0Z_2 ));
    LocalMux I__2060 (
            .O(N__19300),
            .I(\pid_alt.error_d_reg_prevZ0Z_2 ));
    InMux I__2059 (
            .O(N__19293),
            .I(N__19289));
    InMux I__2058 (
            .O(N__19292),
            .I(N__19286));
    LocalMux I__2057 (
            .O(N__19289),
            .I(N__19278));
    LocalMux I__2056 (
            .O(N__19286),
            .I(N__19278));
    InMux I__2055 (
            .O(N__19285),
            .I(N__19275));
    InMux I__2054 (
            .O(N__19284),
            .I(N__19270));
    InMux I__2053 (
            .O(N__19283),
            .I(N__19270));
    Span4Mux_h I__2052 (
            .O(N__19278),
            .I(N__19267));
    LocalMux I__2051 (
            .O(N__19275),
            .I(N__19262));
    LocalMux I__2050 (
            .O(N__19270),
            .I(N__19262));
    Odrv4 I__2049 (
            .O(N__19267),
            .I(\pid_alt.error_p_regZ0Z_2 ));
    Odrv12 I__2048 (
            .O(N__19262),
            .I(\pid_alt.error_p_regZ0Z_2 ));
    InMux I__2047 (
            .O(N__19257),
            .I(N__19253));
    InMux I__2046 (
            .O(N__19256),
            .I(N__19250));
    LocalMux I__2045 (
            .O(N__19253),
            .I(N__19242));
    LocalMux I__2044 (
            .O(N__19250),
            .I(N__19242));
    InMux I__2043 (
            .O(N__19249),
            .I(N__19238));
    InMux I__2042 (
            .O(N__19248),
            .I(N__19233));
    InMux I__2041 (
            .O(N__19247),
            .I(N__19233));
    Span4Mux_h I__2040 (
            .O(N__19242),
            .I(N__19230));
    InMux I__2039 (
            .O(N__19241),
            .I(N__19227));
    LocalMux I__2038 (
            .O(N__19238),
            .I(N__19222));
    LocalMux I__2037 (
            .O(N__19233),
            .I(N__19222));
    Odrv4 I__2036 (
            .O(N__19230),
            .I(\pid_alt.error_d_regZ0Z_2 ));
    LocalMux I__2035 (
            .O(N__19227),
            .I(\pid_alt.error_d_regZ0Z_2 ));
    Odrv4 I__2034 (
            .O(N__19222),
            .I(\pid_alt.error_d_regZ0Z_2 ));
    InMux I__2033 (
            .O(N__19215),
            .I(N__19212));
    LocalMux I__2032 (
            .O(N__19212),
            .I(\pid_alt.error_d_reg_prev_esr_RNI3M511_0Z0Z_3 ));
    CascadeMux I__2031 (
            .O(N__19209),
            .I(\pid_alt.error_d_reg_prev_esr_RNI0J511_0Z0Z_2_cascade_ ));
    InMux I__2030 (
            .O(N__19206),
            .I(N__19203));
    LocalMux I__2029 (
            .O(N__19203),
            .I(\pid_alt.error_d_reg_prev_esr_RNII5LS3Z0Z_2 ));
    InMux I__2028 (
            .O(N__19200),
            .I(N__19193));
    InMux I__2027 (
            .O(N__19199),
            .I(N__19193));
    InMux I__2026 (
            .O(N__19198),
            .I(N__19190));
    LocalMux I__2025 (
            .O(N__19193),
            .I(N__19187));
    LocalMux I__2024 (
            .O(N__19190),
            .I(N__19184));
    Span4Mux_h I__2023 (
            .O(N__19187),
            .I(N__19181));
    Odrv12 I__2022 (
            .O(N__19184),
            .I(\pid_alt.error_p_regZ0Z_3 ));
    Odrv4 I__2021 (
            .O(N__19181),
            .I(\pid_alt.error_p_regZ0Z_3 ));
    InMux I__2020 (
            .O(N__19176),
            .I(N__19169));
    InMux I__2019 (
            .O(N__19175),
            .I(N__19169));
    InMux I__2018 (
            .O(N__19174),
            .I(N__19166));
    LocalMux I__2017 (
            .O(N__19169),
            .I(N__19163));
    LocalMux I__2016 (
            .O(N__19166),
            .I(\pid_alt.error_d_reg_prevZ0Z_3 ));
    Odrv4 I__2015 (
            .O(N__19163),
            .I(\pid_alt.error_d_reg_prevZ0Z_3 ));
    InMux I__2014 (
            .O(N__19158),
            .I(N__19152));
    InMux I__2013 (
            .O(N__19157),
            .I(N__19149));
    InMux I__2012 (
            .O(N__19156),
            .I(N__19144));
    InMux I__2011 (
            .O(N__19155),
            .I(N__19144));
    LocalMux I__2010 (
            .O(N__19152),
            .I(N__19141));
    LocalMux I__2009 (
            .O(N__19149),
            .I(N__19138));
    LocalMux I__2008 (
            .O(N__19144),
            .I(N__19135));
    Span4Mux_v I__2007 (
            .O(N__19141),
            .I(N__19130));
    Span4Mux_h I__2006 (
            .O(N__19138),
            .I(N__19130));
    Span4Mux_h I__2005 (
            .O(N__19135),
            .I(N__19127));
    Odrv4 I__2004 (
            .O(N__19130),
            .I(\pid_alt.error_d_regZ0Z_3 ));
    Odrv4 I__2003 (
            .O(N__19127),
            .I(\pid_alt.error_d_regZ0Z_3 ));
    InMux I__2002 (
            .O(N__19122),
            .I(N__19119));
    LocalMux I__2001 (
            .O(N__19119),
            .I(\pid_alt.error_d_reg_prev_esr_RNI53IMZ0Z_18 ));
    InMux I__2000 (
            .O(N__19116),
            .I(N__19110));
    InMux I__1999 (
            .O(N__19115),
            .I(N__19110));
    LocalMux I__1998 (
            .O(N__19110),
            .I(N__19107));
    Odrv4 I__1997 (
            .O(N__19107),
            .I(\pid_alt.error_d_reg_prev_esr_RNI86IM_0Z0Z_19 ));
    CascadeMux I__1996 (
            .O(N__19104),
            .I(\pid_alt.error_d_reg_prev_esr_RNI53IMZ0Z_18_cascade_ ));
    InMux I__1995 (
            .O(N__19101),
            .I(N__19097));
    InMux I__1994 (
            .O(N__19100),
            .I(N__19094));
    LocalMux I__1993 (
            .O(N__19097),
            .I(\pid_alt.error_d_reg_prevZ0Z_20 ));
    LocalMux I__1992 (
            .O(N__19094),
            .I(\pid_alt.error_d_reg_prevZ0Z_20 ));
    InMux I__1991 (
            .O(N__19089),
            .I(N__19083));
    InMux I__1990 (
            .O(N__19088),
            .I(N__19083));
    LocalMux I__1989 (
            .O(N__19083),
            .I(N__19079));
    InMux I__1988 (
            .O(N__19082),
            .I(N__19076));
    Span4Mux_h I__1987 (
            .O(N__19079),
            .I(N__19073));
    LocalMux I__1986 (
            .O(N__19076),
            .I(N__19070));
    Sp12to4 I__1985 (
            .O(N__19073),
            .I(N__19065));
    Span12Mux_h I__1984 (
            .O(N__19070),
            .I(N__19065));
    Odrv12 I__1983 (
            .O(N__19065),
            .I(\pid_alt.error_d_regZ0Z_20 ));
    InMux I__1982 (
            .O(N__19062),
            .I(N__19059));
    LocalMux I__1981 (
            .O(N__19059),
            .I(N__19056));
    Span4Mux_h I__1980 (
            .O(N__19056),
            .I(N__19053));
    Span4Mux_v I__1979 (
            .O(N__19053),
            .I(N__19050));
    Odrv4 I__1978 (
            .O(N__19050),
            .I(\pid_alt.O_1_7 ));
    InMux I__1977 (
            .O(N__19047),
            .I(N__19044));
    LocalMux I__1976 (
            .O(N__19044),
            .I(N__19041));
    Span4Mux_v I__1975 (
            .O(N__19041),
            .I(N__19038));
    Span4Mux_h I__1974 (
            .O(N__19038),
            .I(N__19035));
    Odrv4 I__1973 (
            .O(N__19035),
            .I(alt_kp_0));
    InMux I__1972 (
            .O(N__19032),
            .I(N__19029));
    LocalMux I__1971 (
            .O(N__19029),
            .I(N__19026));
    Span4Mux_h I__1970 (
            .O(N__19026),
            .I(N__19023));
    Odrv4 I__1969 (
            .O(N__19023),
            .I(alt_kp_6));
    InMux I__1968 (
            .O(N__19020),
            .I(N__19017));
    LocalMux I__1967 (
            .O(N__19017),
            .I(N__19014));
    Span4Mux_s3_h I__1966 (
            .O(N__19014),
            .I(N__19011));
    Odrv4 I__1965 (
            .O(N__19011),
            .I(alt_kp_5));
    InMux I__1964 (
            .O(N__19008),
            .I(N__19005));
    LocalMux I__1963 (
            .O(N__19005),
            .I(N__19002));
    Span4Mux_h I__1962 (
            .O(N__19002),
            .I(N__18999));
    Odrv4 I__1961 (
            .O(N__18999),
            .I(\pid_alt.O_0_16 ));
    InMux I__1960 (
            .O(N__18996),
            .I(N__18993));
    LocalMux I__1959 (
            .O(N__18993),
            .I(N__18989));
    InMux I__1958 (
            .O(N__18992),
            .I(N__18986));
    Span4Mux_v I__1957 (
            .O(N__18989),
            .I(N__18983));
    LocalMux I__1956 (
            .O(N__18986),
            .I(N__18980));
    Span4Mux_h I__1955 (
            .O(N__18983),
            .I(N__18975));
    Span4Mux_h I__1954 (
            .O(N__18980),
            .I(N__18975));
    Odrv4 I__1953 (
            .O(N__18975),
            .I(alt_kd_4));
    CEMux I__1952 (
            .O(N__18972),
            .I(N__18969));
    LocalMux I__1951 (
            .O(N__18969),
            .I(N__18966));
    Span4Mux_h I__1950 (
            .O(N__18966),
            .I(N__18961));
    CEMux I__1949 (
            .O(N__18965),
            .I(N__18958));
    CEMux I__1948 (
            .O(N__18964),
            .I(N__18955));
    Odrv4 I__1947 (
            .O(N__18961),
            .I(\Commands_frame_decoder.source_alt_kd_1_sqmuxa ));
    LocalMux I__1946 (
            .O(N__18958),
            .I(\Commands_frame_decoder.source_alt_kd_1_sqmuxa ));
    LocalMux I__1945 (
            .O(N__18955),
            .I(\Commands_frame_decoder.source_alt_kd_1_sqmuxa ));
    InMux I__1944 (
            .O(N__18948),
            .I(N__18945));
    LocalMux I__1943 (
            .O(N__18945),
            .I(\pid_alt.error_d_reg_prev_esr_RNI0J511_3Z0Z_2 ));
    CascadeMux I__1942 (
            .O(N__18942),
            .I(\pid_alt.error_d_reg_esr_RNITF511_0Z0Z_1_cascade_ ));
    InMux I__1941 (
            .O(N__18939),
            .I(N__18936));
    LocalMux I__1940 (
            .O(N__18936),
            .I(\pid_alt.error_p_reg_esr_RNIL2AQ1Z0Z_0 ));
    InMux I__1939 (
            .O(N__18933),
            .I(N__18930));
    LocalMux I__1938 (
            .O(N__18930),
            .I(\pid_alt.N_1078_0 ));
    InMux I__1937 (
            .O(N__18927),
            .I(N__18924));
    LocalMux I__1936 (
            .O(N__18924),
            .I(N__18915));
    InMux I__1935 (
            .O(N__18923),
            .I(N__18910));
    InMux I__1934 (
            .O(N__18922),
            .I(N__18910));
    InMux I__1933 (
            .O(N__18921),
            .I(N__18907));
    InMux I__1932 (
            .O(N__18920),
            .I(N__18900));
    InMux I__1931 (
            .O(N__18919),
            .I(N__18900));
    InMux I__1930 (
            .O(N__18918),
            .I(N__18900));
    Span4Mux_h I__1929 (
            .O(N__18915),
            .I(N__18895));
    LocalMux I__1928 (
            .O(N__18910),
            .I(N__18895));
    LocalMux I__1927 (
            .O(N__18907),
            .I(N__18890));
    LocalMux I__1926 (
            .O(N__18900),
            .I(N__18890));
    Span4Mux_v I__1925 (
            .O(N__18895),
            .I(N__18887));
    Span4Mux_v I__1924 (
            .O(N__18890),
            .I(N__18884));
    Odrv4 I__1923 (
            .O(N__18887),
            .I(\pid_alt.error_p_regZ0Z_1 ));
    Odrv4 I__1922 (
            .O(N__18884),
            .I(\pid_alt.error_p_regZ0Z_1 ));
    CascadeMux I__1921 (
            .O(N__18879),
            .I(N__18875));
    InMux I__1920 (
            .O(N__18878),
            .I(N__18869));
    InMux I__1919 (
            .O(N__18875),
            .I(N__18864));
    InMux I__1918 (
            .O(N__18874),
            .I(N__18864));
    CascadeMux I__1917 (
            .O(N__18873),
            .I(N__18861));
    InMux I__1916 (
            .O(N__18872),
            .I(N__18856));
    LocalMux I__1915 (
            .O(N__18869),
            .I(N__18851));
    LocalMux I__1914 (
            .O(N__18864),
            .I(N__18851));
    InMux I__1913 (
            .O(N__18861),
            .I(N__18844));
    InMux I__1912 (
            .O(N__18860),
            .I(N__18844));
    InMux I__1911 (
            .O(N__18859),
            .I(N__18844));
    LocalMux I__1910 (
            .O(N__18856),
            .I(\pid_alt.error_d_reg_prevZ0Z_1 ));
    Odrv4 I__1909 (
            .O(N__18851),
            .I(\pid_alt.error_d_reg_prevZ0Z_1 ));
    LocalMux I__1908 (
            .O(N__18844),
            .I(\pid_alt.error_d_reg_prevZ0Z_1 ));
    InMux I__1907 (
            .O(N__18837),
            .I(N__18830));
    InMux I__1906 (
            .O(N__18836),
            .I(N__18830));
    InMux I__1905 (
            .O(N__18835),
            .I(N__18826));
    LocalMux I__1904 (
            .O(N__18830),
            .I(N__18823));
    InMux I__1903 (
            .O(N__18829),
            .I(N__18818));
    LocalMux I__1902 (
            .O(N__18826),
            .I(N__18813));
    Span4Mux_h I__1901 (
            .O(N__18823),
            .I(N__18813));
    InMux I__1900 (
            .O(N__18822),
            .I(N__18808));
    InMux I__1899 (
            .O(N__18821),
            .I(N__18808));
    LocalMux I__1898 (
            .O(N__18818),
            .I(\pid_alt.error_d_regZ0Z_1 ));
    Odrv4 I__1897 (
            .O(N__18813),
            .I(\pid_alt.error_d_regZ0Z_1 ));
    LocalMux I__1896 (
            .O(N__18808),
            .I(\pid_alt.error_d_regZ0Z_1 ));
    InMux I__1895 (
            .O(N__18801),
            .I(N__18798));
    LocalMux I__1894 (
            .O(N__18798),
            .I(\pid_alt.N_1074_1 ));
    CascadeMux I__1893 (
            .O(N__18795),
            .I(\pid_alt.N_3_1_cascade_ ));
    InMux I__1892 (
            .O(N__18792),
            .I(N__18789));
    LocalMux I__1891 (
            .O(N__18789),
            .I(\pid_alt.error_d_reg_prev_esr_RNI0J511_1Z0Z_2 ));
    InMux I__1890 (
            .O(N__18786),
            .I(N__18783));
    LocalMux I__1889 (
            .O(N__18783),
            .I(N__18780));
    Odrv4 I__1888 (
            .O(N__18780),
            .I(\pid_alt.g1_0 ));
    InMux I__1887 (
            .O(N__18777),
            .I(N__18774));
    LocalMux I__1886 (
            .O(N__18774),
            .I(N__18771));
    Span4Mux_s3_h I__1885 (
            .O(N__18771),
            .I(N__18768));
    Odrv4 I__1884 (
            .O(N__18768),
            .I(alt_kp_2));
    InMux I__1883 (
            .O(N__18765),
            .I(N__18762));
    LocalMux I__1882 (
            .O(N__18762),
            .I(N__18759));
    Span4Mux_h I__1881 (
            .O(N__18759),
            .I(N__18756));
    Odrv4 I__1880 (
            .O(N__18756),
            .I(\pid_alt.O_0_22 ));
    InMux I__1879 (
            .O(N__18753),
            .I(N__18749));
    InMux I__1878 (
            .O(N__18752),
            .I(N__18746));
    LocalMux I__1877 (
            .O(N__18749),
            .I(N__18743));
    LocalMux I__1876 (
            .O(N__18746),
            .I(N__18740));
    Span4Mux_v I__1875 (
            .O(N__18743),
            .I(N__18735));
    Span4Mux_v I__1874 (
            .O(N__18740),
            .I(N__18735));
    Odrv4 I__1873 (
            .O(N__18735),
            .I(alt_kd_6));
    InMux I__1872 (
            .O(N__18732),
            .I(N__18728));
    InMux I__1871 (
            .O(N__18731),
            .I(N__18725));
    LocalMux I__1870 (
            .O(N__18728),
            .I(N__18722));
    LocalMux I__1869 (
            .O(N__18725),
            .I(N__18719));
    Span4Mux_s3_h I__1868 (
            .O(N__18722),
            .I(N__18716));
    Span4Mux_s3_h I__1867 (
            .O(N__18719),
            .I(N__18713));
    Odrv4 I__1866 (
            .O(N__18716),
            .I(alt_kd_5));
    Odrv4 I__1865 (
            .O(N__18713),
            .I(alt_kd_5));
    InMux I__1864 (
            .O(N__18708),
            .I(N__18705));
    LocalMux I__1863 (
            .O(N__18705),
            .I(N__18702));
    Odrv4 I__1862 (
            .O(N__18702),
            .I(\pid_alt.O_4 ));
    InMux I__1861 (
            .O(N__18699),
            .I(N__18696));
    LocalMux I__1860 (
            .O(N__18696),
            .I(\pid_alt.N_1074_0 ));
    InMux I__1859 (
            .O(N__18693),
            .I(N__18690));
    LocalMux I__1858 (
            .O(N__18690),
            .I(\pid_alt.N_5_0 ));
    InMux I__1857 (
            .O(N__18687),
            .I(N__18684));
    LocalMux I__1856 (
            .O(N__18684),
            .I(\pid_alt.g1_1 ));
    CascadeMux I__1855 (
            .O(N__18681),
            .I(\pid_alt.N_1080_0_cascade_ ));
    InMux I__1854 (
            .O(N__18678),
            .I(N__18674));
    InMux I__1853 (
            .O(N__18677),
            .I(N__18671));
    LocalMux I__1852 (
            .O(N__18674),
            .I(N__18666));
    LocalMux I__1851 (
            .O(N__18671),
            .I(N__18666));
    Span4Mux_h I__1850 (
            .O(N__18666),
            .I(N__18663));
    Odrv4 I__1849 (
            .O(N__18663),
            .I(\pid_alt.error_d_reg_fastZ0Z_1 ));
    CascadeMux I__1848 (
            .O(N__18660),
            .I(N__18657));
    InMux I__1847 (
            .O(N__18657),
            .I(N__18654));
    LocalMux I__1846 (
            .O(N__18654),
            .I(\pid_alt.N_3_0 ));
    InMux I__1845 (
            .O(N__18651),
            .I(N__18646));
    InMux I__1844 (
            .O(N__18650),
            .I(N__18641));
    InMux I__1843 (
            .O(N__18649),
            .I(N__18641));
    LocalMux I__1842 (
            .O(N__18646),
            .I(N__18636));
    LocalMux I__1841 (
            .O(N__18641),
            .I(N__18636));
    Span4Mux_v I__1840 (
            .O(N__18636),
            .I(N__18633));
    Span4Mux_v I__1839 (
            .O(N__18633),
            .I(N__18630));
    Odrv4 I__1838 (
            .O(N__18630),
            .I(\pid_alt.error_d_regZ0Z_19 ));
    CascadeMux I__1837 (
            .O(N__18627),
            .I(N__18624));
    InMux I__1836 (
            .O(N__18624),
            .I(N__18618));
    InMux I__1835 (
            .O(N__18623),
            .I(N__18618));
    LocalMux I__1834 (
            .O(N__18618),
            .I(\pid_alt.error_d_reg_prevZ0Z_19 ));
    InMux I__1833 (
            .O(N__18615),
            .I(N__18609));
    InMux I__1832 (
            .O(N__18614),
            .I(N__18609));
    LocalMux I__1831 (
            .O(N__18609),
            .I(N__18606));
    Span4Mux_v I__1830 (
            .O(N__18606),
            .I(N__18603));
    Odrv4 I__1829 (
            .O(N__18603),
            .I(\pid_alt.error_p_regZ0Z_19 ));
    InMux I__1828 (
            .O(N__18600),
            .I(N__18597));
    LocalMux I__1827 (
            .O(N__18597),
            .I(N__18594));
    Span12Mux_v I__1826 (
            .O(N__18594),
            .I(N__18591));
    Odrv12 I__1825 (
            .O(N__18591),
            .I(\pid_alt.O_1_6 ));
    InMux I__1824 (
            .O(N__18588),
            .I(N__18585));
    LocalMux I__1823 (
            .O(N__18585),
            .I(N__18582));
    Span4Mux_h I__1822 (
            .O(N__18582),
            .I(N__18579));
    Span4Mux_v I__1821 (
            .O(N__18579),
            .I(N__18576));
    Odrv4 I__1820 (
            .O(N__18576),
            .I(\pid_alt.O_1_5 ));
    InMux I__1819 (
            .O(N__18573),
            .I(N__18570));
    LocalMux I__1818 (
            .O(N__18570),
            .I(N__18567));
    Span12Mux_v I__1817 (
            .O(N__18567),
            .I(N__18564));
    Odrv12 I__1816 (
            .O(N__18564),
            .I(\pid_alt.O_1_14 ));
    InMux I__1815 (
            .O(N__18561),
            .I(N__18558));
    LocalMux I__1814 (
            .O(N__18558),
            .I(N__18555));
    Span4Mux_s2_h I__1813 (
            .O(N__18555),
            .I(N__18552));
    Span4Mux_v I__1812 (
            .O(N__18552),
            .I(N__18549));
    Odrv4 I__1811 (
            .O(N__18549),
            .I(alt_kp_3));
    InMux I__1810 (
            .O(N__18546),
            .I(N__18543));
    LocalMux I__1809 (
            .O(N__18543),
            .I(N__18540));
    Span4Mux_s2_h I__1808 (
            .O(N__18540),
            .I(N__18537));
    Odrv4 I__1807 (
            .O(N__18537),
            .I(alt_kp_1));
    InMux I__1806 (
            .O(N__18534),
            .I(N__18531));
    LocalMux I__1805 (
            .O(N__18531),
            .I(N__18528));
    Span4Mux_s2_h I__1804 (
            .O(N__18528),
            .I(N__18525));
    Odrv4 I__1803 (
            .O(N__18525),
            .I(alt_kp_7));
    CascadeMux I__1802 (
            .O(N__18522),
            .I(\pid_alt.g0_0_0_cascade_ ));
    InMux I__1801 (
            .O(N__18519),
            .I(N__18516));
    LocalMux I__1800 (
            .O(N__18516),
            .I(N__18513));
    Odrv4 I__1799 (
            .O(N__18513),
            .I(\pid_alt.O_0_18 ));
    InMux I__1798 (
            .O(N__18510),
            .I(N__18507));
    LocalMux I__1797 (
            .O(N__18507),
            .I(\pid_alt.O_0_19 ));
    InMux I__1796 (
            .O(N__18504),
            .I(N__18501));
    LocalMux I__1795 (
            .O(N__18501),
            .I(N__18497));
    InMux I__1794 (
            .O(N__18500),
            .I(N__18494));
    Span4Mux_v I__1793 (
            .O(N__18497),
            .I(N__18491));
    LocalMux I__1792 (
            .O(N__18494),
            .I(N__18488));
    Span4Mux_v I__1791 (
            .O(N__18491),
            .I(N__18485));
    Span12Mux_s11_v I__1790 (
            .O(N__18488),
            .I(N__18482));
    Span4Mux_v I__1789 (
            .O(N__18485),
            .I(N__18479));
    Odrv12 I__1788 (
            .O(N__18482),
            .I(\pid_alt.error_p_regZ0Z_17 ));
    Odrv4 I__1787 (
            .O(N__18479),
            .I(\pid_alt.error_p_regZ0Z_17 ));
    InMux I__1786 (
            .O(N__18474),
            .I(N__18470));
    InMux I__1785 (
            .O(N__18473),
            .I(N__18467));
    LocalMux I__1784 (
            .O(N__18470),
            .I(\pid_alt.error_d_reg_prevZ0Z_17 ));
    LocalMux I__1783 (
            .O(N__18467),
            .I(\pid_alt.error_d_reg_prevZ0Z_17 ));
    InMux I__1782 (
            .O(N__18462),
            .I(N__18457));
    InMux I__1781 (
            .O(N__18461),
            .I(N__18454));
    InMux I__1780 (
            .O(N__18460),
            .I(N__18451));
    LocalMux I__1779 (
            .O(N__18457),
            .I(N__18444));
    LocalMux I__1778 (
            .O(N__18454),
            .I(N__18444));
    LocalMux I__1777 (
            .O(N__18451),
            .I(N__18444));
    Odrv4 I__1776 (
            .O(N__18444),
            .I(\pid_alt.error_d_regZ0Z_17 ));
    InMux I__1775 (
            .O(N__18441),
            .I(N__18437));
    InMux I__1774 (
            .O(N__18440),
            .I(N__18434));
    LocalMux I__1773 (
            .O(N__18437),
            .I(N__18431));
    LocalMux I__1772 (
            .O(N__18434),
            .I(N__18428));
    Span4Mux_s2_h I__1771 (
            .O(N__18431),
            .I(N__18425));
    Span4Mux_s2_h I__1770 (
            .O(N__18428),
            .I(N__18422));
    Odrv4 I__1769 (
            .O(N__18425),
            .I(alt_kd_2));
    Odrv4 I__1768 (
            .O(N__18422),
            .I(alt_kd_2));
    InMux I__1767 (
            .O(N__18417),
            .I(N__18413));
    InMux I__1766 (
            .O(N__18416),
            .I(N__18410));
    LocalMux I__1765 (
            .O(N__18413),
            .I(N__18407));
    LocalMux I__1764 (
            .O(N__18410),
            .I(N__18404));
    Span4Mux_s3_h I__1763 (
            .O(N__18407),
            .I(N__18401));
    Span4Mux_v I__1762 (
            .O(N__18404),
            .I(N__18398));
    Odrv4 I__1761 (
            .O(N__18401),
            .I(alt_kd_3));
    Odrv4 I__1760 (
            .O(N__18398),
            .I(alt_kd_3));
    InMux I__1759 (
            .O(N__18393),
            .I(N__18389));
    InMux I__1758 (
            .O(N__18392),
            .I(N__18386));
    LocalMux I__1757 (
            .O(N__18389),
            .I(N__18383));
    LocalMux I__1756 (
            .O(N__18386),
            .I(N__18380));
    Span4Mux_s2_h I__1755 (
            .O(N__18383),
            .I(N__18377));
    Span4Mux_v I__1754 (
            .O(N__18380),
            .I(N__18374));
    Odrv4 I__1753 (
            .O(N__18377),
            .I(alt_kd_7));
    Odrv4 I__1752 (
            .O(N__18374),
            .I(alt_kd_7));
    InMux I__1751 (
            .O(N__18369),
            .I(N__18365));
    InMux I__1750 (
            .O(N__18368),
            .I(N__18362));
    LocalMux I__1749 (
            .O(N__18365),
            .I(N__18359));
    LocalMux I__1748 (
            .O(N__18362),
            .I(N__18356));
    Span12Mux_s9_v I__1747 (
            .O(N__18359),
            .I(N__18353));
    Span4Mux_s2_h I__1746 (
            .O(N__18356),
            .I(N__18350));
    Odrv12 I__1745 (
            .O(N__18353),
            .I(alt_kd_1));
    Odrv4 I__1744 (
            .O(N__18350),
            .I(alt_kd_1));
    InMux I__1743 (
            .O(N__18345),
            .I(N__18342));
    LocalMux I__1742 (
            .O(N__18342),
            .I(N__18338));
    InMux I__1741 (
            .O(N__18341),
            .I(N__18335));
    Span4Mux_s1_h I__1740 (
            .O(N__18338),
            .I(N__18332));
    LocalMux I__1739 (
            .O(N__18335),
            .I(N__18329));
    Span4Mux_v I__1738 (
            .O(N__18332),
            .I(N__18326));
    Span4Mux_s2_h I__1737 (
            .O(N__18329),
            .I(N__18323));
    Odrv4 I__1736 (
            .O(N__18326),
            .I(alt_kd_0));
    Odrv4 I__1735 (
            .O(N__18323),
            .I(alt_kd_0));
    CascadeMux I__1734 (
            .O(N__18318),
            .I(N__18311));
    CascadeMux I__1733 (
            .O(N__18317),
            .I(N__18307));
    CascadeMux I__1732 (
            .O(N__18316),
            .I(N__18303));
    InMux I__1731 (
            .O(N__18315),
            .I(N__18288));
    InMux I__1730 (
            .O(N__18314),
            .I(N__18288));
    InMux I__1729 (
            .O(N__18311),
            .I(N__18288));
    InMux I__1728 (
            .O(N__18310),
            .I(N__18288));
    InMux I__1727 (
            .O(N__18307),
            .I(N__18288));
    InMux I__1726 (
            .O(N__18306),
            .I(N__18288));
    InMux I__1725 (
            .O(N__18303),
            .I(N__18288));
    LocalMux I__1724 (
            .O(N__18288),
            .I(\pid_alt.O_1_21 ));
    InMux I__1723 (
            .O(N__18285),
            .I(\pid_alt.error_filt_cry_21 ));
    InMux I__1722 (
            .O(N__18282),
            .I(N__18279));
    LocalMux I__1721 (
            .O(N__18279),
            .I(N__18276));
    Span4Mux_v I__1720 (
            .O(N__18276),
            .I(N__18273));
    Odrv4 I__1719 (
            .O(N__18273),
            .I(\pid_alt.O_1_11 ));
    InMux I__1718 (
            .O(N__18270),
            .I(N__18267));
    LocalMux I__1717 (
            .O(N__18267),
            .I(N__18264));
    Span4Mux_h I__1716 (
            .O(N__18264),
            .I(N__18261));
    Odrv4 I__1715 (
            .O(N__18261),
            .I(\pid_alt.O_1_12 ));
    InMux I__1714 (
            .O(N__18258),
            .I(N__18255));
    LocalMux I__1713 (
            .O(N__18255),
            .I(N__18252));
    Odrv4 I__1712 (
            .O(N__18252),
            .I(\pid_alt.O_1_10 ));
    InMux I__1711 (
            .O(N__18249),
            .I(N__18246));
    LocalMux I__1710 (
            .O(N__18246),
            .I(N__18243));
    Span4Mux_h I__1709 (
            .O(N__18243),
            .I(N__18240));
    Odrv4 I__1708 (
            .O(N__18240),
            .I(\pid_alt.O_0_17 ));
    InMux I__1707 (
            .O(N__18237),
            .I(N__18234));
    LocalMux I__1706 (
            .O(N__18234),
            .I(N__18231));
    Odrv4 I__1705 (
            .O(N__18231),
            .I(\pid_alt.O_0_20 ));
    InMux I__1704 (
            .O(N__18228),
            .I(N__18225));
    LocalMux I__1703 (
            .O(N__18225),
            .I(N__18222));
    Span4Mux_h I__1702 (
            .O(N__18222),
            .I(N__18219));
    Odrv4 I__1701 (
            .O(N__18219),
            .I(\pid_alt.O_0_23 ));
    InMux I__1700 (
            .O(N__18216),
            .I(N__18213));
    LocalMux I__1699 (
            .O(N__18213),
            .I(N__18210));
    Odrv4 I__1698 (
            .O(N__18210),
            .I(\pid_alt.O_1_13 ));
    InMux I__1697 (
            .O(N__18207),
            .I(N__18204));
    LocalMux I__1696 (
            .O(N__18204),
            .I(N__18201));
    Odrv4 I__1695 (
            .O(N__18201),
            .I(\pid_alt.O_0_21 ));
    InMux I__1694 (
            .O(N__18198),
            .I(N__18195));
    LocalMux I__1693 (
            .O(N__18195),
            .I(N__18192));
    Odrv4 I__1692 (
            .O(N__18192),
            .I(\pid_alt.O_0_24 ));
    InMux I__1691 (
            .O(N__18189),
            .I(N__18186));
    LocalMux I__1690 (
            .O(N__18186),
            .I(\pid_alt.O_1_19 ));
    InMux I__1689 (
            .O(N__18183),
            .I(\pid_alt.error_filt_cry_13 ));
    CascadeMux I__1688 (
            .O(N__18180),
            .I(N__18177));
    InMux I__1687 (
            .O(N__18177),
            .I(N__18174));
    LocalMux I__1686 (
            .O(N__18174),
            .I(\pid_alt.O_1_20 ));
    InMux I__1685 (
            .O(N__18171),
            .I(\pid_alt.error_filt_cry_14 ));
    InMux I__1684 (
            .O(N__18168),
            .I(bfn_1_18_0_));
    InMux I__1683 (
            .O(N__18165),
            .I(\pid_alt.error_filt_cry_16 ));
    InMux I__1682 (
            .O(N__18162),
            .I(\pid_alt.error_filt_cry_17 ));
    InMux I__1681 (
            .O(N__18159),
            .I(\pid_alt.error_filt_cry_18 ));
    InMux I__1680 (
            .O(N__18156),
            .I(\pid_alt.error_filt_cry_19 ));
    InMux I__1679 (
            .O(N__18153),
            .I(\pid_alt.error_filt_cry_20 ));
    InMux I__1678 (
            .O(N__18150),
            .I(\pid_alt.error_filt_cry_4 ));
    InMux I__1677 (
            .O(N__18147),
            .I(N__18144));
    LocalMux I__1676 (
            .O(N__18144),
            .I(N__18141));
    Span4Mux_s2_h I__1675 (
            .O(N__18141),
            .I(N__18138));
    Span4Mux_h I__1674 (
            .O(N__18138),
            .I(N__18135));
    Span4Mux_h I__1673 (
            .O(N__18135),
            .I(N__18132));
    Span4Mux_h I__1672 (
            .O(N__18132),
            .I(N__18129));
    Span4Mux_h I__1671 (
            .O(N__18129),
            .I(N__18126));
    Span4Mux_h I__1670 (
            .O(N__18126),
            .I(N__18123));
    Odrv4 I__1669 (
            .O(N__18123),
            .I(\pid_alt.O_3_11 ));
    CascadeMux I__1668 (
            .O(N__18120),
            .I(N__18117));
    InMux I__1667 (
            .O(N__18117),
            .I(N__18114));
    LocalMux I__1666 (
            .O(N__18114),
            .I(\pid_alt.O_2_11 ));
    InMux I__1665 (
            .O(N__18111),
            .I(\pid_alt.error_filt_cry_5 ));
    InMux I__1664 (
            .O(N__18108),
            .I(N__18105));
    LocalMux I__1663 (
            .O(N__18105),
            .I(\pid_alt.O_2_12 ));
    CascadeMux I__1662 (
            .O(N__18102),
            .I(N__18099));
    InMux I__1661 (
            .O(N__18099),
            .I(N__18096));
    LocalMux I__1660 (
            .O(N__18096),
            .I(N__18093));
    Span4Mux_h I__1659 (
            .O(N__18093),
            .I(N__18090));
    Sp12to4 I__1658 (
            .O(N__18090),
            .I(N__18087));
    Span12Mux_h I__1657 (
            .O(N__18087),
            .I(N__18084));
    Odrv12 I__1656 (
            .O(N__18084),
            .I(\pid_alt.O_3_12 ));
    InMux I__1655 (
            .O(N__18081),
            .I(\pid_alt.error_filt_cry_6 ));
    InMux I__1654 (
            .O(N__18078),
            .I(N__18075));
    LocalMux I__1653 (
            .O(N__18075),
            .I(N__18072));
    Span12Mux_v I__1652 (
            .O(N__18072),
            .I(N__18069));
    Span12Mux_h I__1651 (
            .O(N__18069),
            .I(N__18066));
    Span12Mux_h I__1650 (
            .O(N__18066),
            .I(N__18063));
    Odrv12 I__1649 (
            .O(N__18063),
            .I(\pid_alt.O_3_13 ));
    CascadeMux I__1648 (
            .O(N__18060),
            .I(N__18057));
    InMux I__1647 (
            .O(N__18057),
            .I(N__18054));
    LocalMux I__1646 (
            .O(N__18054),
            .I(\pid_alt.O_2_13 ));
    InMux I__1645 (
            .O(N__18051),
            .I(bfn_1_17_0_));
    InMux I__1644 (
            .O(N__18048),
            .I(N__18045));
    LocalMux I__1643 (
            .O(N__18045),
            .I(N__18042));
    Span4Mux_v I__1642 (
            .O(N__18042),
            .I(N__18039));
    Sp12to4 I__1641 (
            .O(N__18039),
            .I(N__18036));
    Span12Mux_h I__1640 (
            .O(N__18036),
            .I(N__18033));
    Odrv12 I__1639 (
            .O(N__18033),
            .I(\pid_alt.O_3_14 ));
    CascadeMux I__1638 (
            .O(N__18030),
            .I(N__18027));
    InMux I__1637 (
            .O(N__18027),
            .I(N__18024));
    LocalMux I__1636 (
            .O(N__18024),
            .I(\pid_alt.O_2_14 ));
    InMux I__1635 (
            .O(N__18021),
            .I(\pid_alt.error_filt_cry_8 ));
    CascadeMux I__1634 (
            .O(N__18018),
            .I(N__18015));
    InMux I__1633 (
            .O(N__18015),
            .I(N__18012));
    LocalMux I__1632 (
            .O(N__18012),
            .I(\pid_alt.O_1_15 ));
    InMux I__1631 (
            .O(N__18009),
            .I(\pid_alt.error_filt_cry_9 ));
    CascadeMux I__1630 (
            .O(N__18006),
            .I(N__18003));
    InMux I__1629 (
            .O(N__18003),
            .I(N__18000));
    LocalMux I__1628 (
            .O(N__18000),
            .I(\pid_alt.O_1_16 ));
    InMux I__1627 (
            .O(N__17997),
            .I(\pid_alt.error_filt_cry_10 ));
    CascadeMux I__1626 (
            .O(N__17994),
            .I(N__17991));
    InMux I__1625 (
            .O(N__17991),
            .I(N__17988));
    LocalMux I__1624 (
            .O(N__17988),
            .I(\pid_alt.O_1_17 ));
    InMux I__1623 (
            .O(N__17985),
            .I(\pid_alt.error_filt_cry_11 ));
    CascadeMux I__1622 (
            .O(N__17982),
            .I(N__17979));
    InMux I__1621 (
            .O(N__17979),
            .I(N__17976));
    LocalMux I__1620 (
            .O(N__17976),
            .I(\pid_alt.O_1_18 ));
    InMux I__1619 (
            .O(N__17973),
            .I(\pid_alt.error_filt_cry_12 ));
    InMux I__1618 (
            .O(N__17970),
            .I(N__17967));
    LocalMux I__1617 (
            .O(N__17967),
            .I(N__17964));
    Span12Mux_h I__1616 (
            .O(N__17964),
            .I(N__17961));
    Odrv12 I__1615 (
            .O(N__17961),
            .I(\pid_alt.O_1_4 ));
    InMux I__1614 (
            .O(N__17958),
            .I(N__17955));
    LocalMux I__1613 (
            .O(N__17955),
            .I(N__17952));
    Span4Mux_s3_h I__1612 (
            .O(N__17952),
            .I(N__17949));
    Span4Mux_h I__1611 (
            .O(N__17949),
            .I(N__17946));
    Span4Mux_h I__1610 (
            .O(N__17946),
            .I(N__17943));
    Span4Mux_h I__1609 (
            .O(N__17943),
            .I(N__17940));
    Span4Mux_h I__1608 (
            .O(N__17940),
            .I(N__17937));
    Span4Mux_h I__1607 (
            .O(N__17937),
            .I(N__17934));
    Odrv4 I__1606 (
            .O(N__17934),
            .I(\pid_alt.error_filt_prevZ0Z_0 ));
    InMux I__1605 (
            .O(N__17931),
            .I(N__17927));
    InMux I__1604 (
            .O(N__17930),
            .I(N__17924));
    LocalMux I__1603 (
            .O(N__17927),
            .I(N__17921));
    LocalMux I__1602 (
            .O(N__17924),
            .I(N__17918));
    Span12Mux_v I__1601 (
            .O(N__17921),
            .I(N__17915));
    Span12Mux_s4_h I__1600 (
            .O(N__17918),
            .I(N__17912));
    Span12Mux_h I__1599 (
            .O(N__17915),
            .I(N__17909));
    Span12Mux_h I__1598 (
            .O(N__17912),
            .I(N__17906));
    Span12Mux_h I__1597 (
            .O(N__17909),
            .I(N__17903));
    Odrv12 I__1596 (
            .O(N__17906),
            .I(\pid_alt.error_filt ));
    Odrv12 I__1595 (
            .O(N__17903),
            .I(\pid_alt.error_filt ));
    CascadeMux I__1594 (
            .O(N__17898),
            .I(N__17894));
    InMux I__1593 (
            .O(N__17897),
            .I(N__17891));
    InMux I__1592 (
            .O(N__17894),
            .I(N__17888));
    LocalMux I__1591 (
            .O(N__17891),
            .I(\pid_alt.O_2_5 ));
    LocalMux I__1590 (
            .O(N__17888),
            .I(\pid_alt.O_2_5 ));
    InMux I__1589 (
            .O(N__17883),
            .I(N__17880));
    LocalMux I__1588 (
            .O(N__17880),
            .I(N__17877));
    Span4Mux_s2_h I__1587 (
            .O(N__17877),
            .I(N__17874));
    Odrv4 I__1586 (
            .O(N__17874),
            .I(\pid_alt.error_filt_0 ));
    InMux I__1585 (
            .O(N__17871),
            .I(N__17868));
    LocalMux I__1584 (
            .O(N__17868),
            .I(N__17865));
    Span4Mux_v I__1583 (
            .O(N__17865),
            .I(N__17862));
    Sp12to4 I__1582 (
            .O(N__17862),
            .I(N__17859));
    Span12Mux_h I__1581 (
            .O(N__17859),
            .I(N__17856));
    Odrv12 I__1580 (
            .O(N__17856),
            .I(\pid_alt.O_3_6 ));
    CascadeMux I__1579 (
            .O(N__17853),
            .I(N__17850));
    InMux I__1578 (
            .O(N__17850),
            .I(N__17847));
    LocalMux I__1577 (
            .O(N__17847),
            .I(\pid_alt.O_2_6 ));
    InMux I__1576 (
            .O(N__17844),
            .I(\pid_alt.error_filt_cry_0 ));
    InMux I__1575 (
            .O(N__17841),
            .I(N__17838));
    LocalMux I__1574 (
            .O(N__17838),
            .I(N__17835));
    Span4Mux_v I__1573 (
            .O(N__17835),
            .I(N__17832));
    Sp12to4 I__1572 (
            .O(N__17832),
            .I(N__17829));
    Span12Mux_h I__1571 (
            .O(N__17829),
            .I(N__17826));
    Odrv12 I__1570 (
            .O(N__17826),
            .I(\pid_alt.O_3_7 ));
    CascadeMux I__1569 (
            .O(N__17823),
            .I(N__17820));
    InMux I__1568 (
            .O(N__17820),
            .I(N__17817));
    LocalMux I__1567 (
            .O(N__17817),
            .I(\pid_alt.O_2_7 ));
    InMux I__1566 (
            .O(N__17814),
            .I(\pid_alt.error_filt_cry_1 ));
    InMux I__1565 (
            .O(N__17811),
            .I(N__17808));
    LocalMux I__1564 (
            .O(N__17808),
            .I(N__17805));
    Span12Mux_s9_h I__1563 (
            .O(N__17805),
            .I(N__17802));
    Span12Mux_h I__1562 (
            .O(N__17802),
            .I(N__17799));
    Odrv12 I__1561 (
            .O(N__17799),
            .I(\pid_alt.O_3_8 ));
    CascadeMux I__1560 (
            .O(N__17796),
            .I(N__17793));
    InMux I__1559 (
            .O(N__17793),
            .I(N__17790));
    LocalMux I__1558 (
            .O(N__17790),
            .I(\pid_alt.O_2_8 ));
    InMux I__1557 (
            .O(N__17787),
            .I(\pid_alt.error_filt_cry_2 ));
    InMux I__1556 (
            .O(N__17784),
            .I(N__17781));
    LocalMux I__1555 (
            .O(N__17781),
            .I(N__17778));
    Span12Mux_v I__1554 (
            .O(N__17778),
            .I(N__17775));
    Span12Mux_h I__1553 (
            .O(N__17775),
            .I(N__17772));
    Span12Mux_h I__1552 (
            .O(N__17772),
            .I(N__17769));
    Odrv12 I__1551 (
            .O(N__17769),
            .I(\pid_alt.O_3_9 ));
    CascadeMux I__1550 (
            .O(N__17766),
            .I(N__17763));
    InMux I__1549 (
            .O(N__17763),
            .I(N__17760));
    LocalMux I__1548 (
            .O(N__17760),
            .I(\pid_alt.O_2_9 ));
    InMux I__1547 (
            .O(N__17757),
            .I(\pid_alt.error_filt_cry_3 ));
    InMux I__1546 (
            .O(N__17754),
            .I(N__17751));
    LocalMux I__1545 (
            .O(N__17751),
            .I(\pid_alt.O_2_10 ));
    CascadeMux I__1544 (
            .O(N__17748),
            .I(N__17745));
    InMux I__1543 (
            .O(N__17745),
            .I(N__17742));
    LocalMux I__1542 (
            .O(N__17742),
            .I(N__17739));
    Span12Mux_s7_h I__1541 (
            .O(N__17739),
            .I(N__17736));
    Span12Mux_h I__1540 (
            .O(N__17736),
            .I(N__17733));
    Odrv12 I__1539 (
            .O(N__17733),
            .I(\pid_alt.O_3_10 ));
    InMux I__1538 (
            .O(N__17730),
            .I(N__17727));
    LocalMux I__1537 (
            .O(N__17727),
            .I(\pid_alt.O_13 ));
    InMux I__1536 (
            .O(N__17724),
            .I(N__17721));
    LocalMux I__1535 (
            .O(N__17721),
            .I(\pid_alt.O_11 ));
    CascadeMux I__1534 (
            .O(N__17718),
            .I(N__17715));
    InMux I__1533 (
            .O(N__17715),
            .I(N__17709));
    InMux I__1532 (
            .O(N__17714),
            .I(N__17709));
    LocalMux I__1531 (
            .O(N__17709),
            .I(\pid_alt.O_5 ));
    InMux I__1530 (
            .O(N__17706),
            .I(N__17703));
    LocalMux I__1529 (
            .O(N__17703),
            .I(\pid_alt.O_14 ));
    InMux I__1528 (
            .O(N__17700),
            .I(N__17697));
    LocalMux I__1527 (
            .O(N__17697),
            .I(\pid_alt.O_6 ));
    InMux I__1526 (
            .O(N__17694),
            .I(N__17691));
    LocalMux I__1525 (
            .O(N__17691),
            .I(\pid_alt.O_12 ));
    InMux I__1524 (
            .O(N__17688),
            .I(N__17685));
    LocalMux I__1523 (
            .O(N__17685),
            .I(\pid_alt.O_9 ));
    InMux I__1522 (
            .O(N__17682),
            .I(N__17679));
    LocalMux I__1521 (
            .O(N__17679),
            .I(N__17676));
    Odrv4 I__1520 (
            .O(N__17676),
            .I(\pid_alt.O_7 ));
    InMux I__1519 (
            .O(N__17673),
            .I(\pid_alt.un1_error_d_reg_add_1_cry_10 ));
    CascadeMux I__1518 (
            .O(N__17670),
            .I(N__17667));
    InMux I__1517 (
            .O(N__17667),
            .I(N__17664));
    LocalMux I__1516 (
            .O(N__17664),
            .I(\pid_alt.un1_error_d_reg_2_12 ));
    InMux I__1515 (
            .O(N__17661),
            .I(\pid_alt.un1_error_d_reg_add_1_cry_11 ));
    CascadeMux I__1514 (
            .O(N__17658),
            .I(N__17655));
    InMux I__1513 (
            .O(N__17655),
            .I(N__17652));
    LocalMux I__1512 (
            .O(N__17652),
            .I(\pid_alt.un1_error_d_reg_2_13 ));
    InMux I__1511 (
            .O(N__17649),
            .I(\pid_alt.un1_error_d_reg_add_1_cry_12 ));
    CascadeMux I__1510 (
            .O(N__17646),
            .I(N__17643));
    InMux I__1509 (
            .O(N__17643),
            .I(N__17640));
    LocalMux I__1508 (
            .O(N__17640),
            .I(\pid_alt.un1_error_d_reg_2_14 ));
    InMux I__1507 (
            .O(N__17637),
            .I(\pid_alt.un1_error_d_reg_add_1_cry_13 ));
    CascadeMux I__1506 (
            .O(N__17634),
            .I(N__17631));
    InMux I__1505 (
            .O(N__17631),
            .I(N__17628));
    LocalMux I__1504 (
            .O(N__17628),
            .I(\pid_alt.un1_error_d_reg_2_15 ));
    InMux I__1503 (
            .O(N__17625),
            .I(\pid_alt.un1_error_d_reg_add_1_cry_14 ));
    InMux I__1502 (
            .O(N__17622),
            .I(N__17612));
    InMux I__1501 (
            .O(N__17621),
            .I(N__17605));
    InMux I__1500 (
            .O(N__17620),
            .I(N__17605));
    InMux I__1499 (
            .O(N__17619),
            .I(N__17605));
    InMux I__1498 (
            .O(N__17618),
            .I(N__17596));
    InMux I__1497 (
            .O(N__17617),
            .I(N__17596));
    InMux I__1496 (
            .O(N__17616),
            .I(N__17596));
    InMux I__1495 (
            .O(N__17615),
            .I(N__17596));
    LocalMux I__1494 (
            .O(N__17612),
            .I(N__17591));
    LocalMux I__1493 (
            .O(N__17605),
            .I(N__17591));
    LocalMux I__1492 (
            .O(N__17596),
            .I(N__17588));
    Span4Mux_v I__1491 (
            .O(N__17591),
            .I(N__17585));
    Span4Mux_v I__1490 (
            .O(N__17588),
            .I(N__17582));
    Odrv4 I__1489 (
            .O(N__17585),
            .I(\pid_alt.un1_error_d_reg_1_24 ));
    Odrv4 I__1488 (
            .O(N__17582),
            .I(\pid_alt.un1_error_d_reg_1_24 ));
    CascadeMux I__1487 (
            .O(N__17577),
            .I(N__17574));
    InMux I__1486 (
            .O(N__17574),
            .I(N__17571));
    LocalMux I__1485 (
            .O(N__17571),
            .I(\pid_alt.un1_error_d_reg_2_16 ));
    InMux I__1484 (
            .O(N__17568),
            .I(bfn_1_8_0_));
    InMux I__1483 (
            .O(N__17565),
            .I(N__17562));
    LocalMux I__1482 (
            .O(N__17562),
            .I(N__17559));
    Odrv4 I__1481 (
            .O(N__17559),
            .I(\pid_alt.O_10 ));
    InMux I__1480 (
            .O(N__17556),
            .I(N__17553));
    LocalMux I__1479 (
            .O(N__17553),
            .I(N__17550));
    Span4Mux_v I__1478 (
            .O(N__17550),
            .I(N__17546));
    InMux I__1477 (
            .O(N__17549),
            .I(N__17543));
    Odrv4 I__1476 (
            .O(N__17546),
            .I(\pid_alt.un1_error_d_reg_2_0 ));
    LocalMux I__1475 (
            .O(N__17543),
            .I(\pid_alt.un1_error_d_reg_2_0 ));
    CascadeMux I__1474 (
            .O(N__17538),
            .I(N__17535));
    InMux I__1473 (
            .O(N__17535),
            .I(N__17531));
    InMux I__1472 (
            .O(N__17534),
            .I(N__17528));
    LocalMux I__1471 (
            .O(N__17531),
            .I(N__17525));
    LocalMux I__1470 (
            .O(N__17528),
            .I(N__17520));
    Span4Mux_v I__1469 (
            .O(N__17525),
            .I(N__17520));
    Odrv4 I__1468 (
            .O(N__17520),
            .I(\pid_alt.un1_error_d_reg_1_15 ));
    InMux I__1467 (
            .O(N__17517),
            .I(\pid_alt.un1_error_d_reg_add_1_cry_2 ));
    InMux I__1466 (
            .O(N__17514),
            .I(N__17511));
    LocalMux I__1465 (
            .O(N__17511),
            .I(N__17508));
    Odrv4 I__1464 (
            .O(N__17508),
            .I(\pid_alt.un1_error_d_reg_2_4 ));
    CascadeMux I__1463 (
            .O(N__17505),
            .I(N__17502));
    InMux I__1462 (
            .O(N__17502),
            .I(N__17499));
    LocalMux I__1461 (
            .O(N__17499),
            .I(N__17496));
    Span4Mux_v I__1460 (
            .O(N__17496),
            .I(N__17493));
    Odrv4 I__1459 (
            .O(N__17493),
            .I(\pid_alt.un1_error_d_reg_1_19 ));
    InMux I__1458 (
            .O(N__17490),
            .I(\pid_alt.un1_error_d_reg_add_1_cry_3 ));
    InMux I__1457 (
            .O(N__17487),
            .I(N__17484));
    LocalMux I__1456 (
            .O(N__17484),
            .I(\pid_alt.un1_error_d_reg_2_5 ));
    CascadeMux I__1455 (
            .O(N__17481),
            .I(N__17478));
    InMux I__1454 (
            .O(N__17478),
            .I(N__17475));
    LocalMux I__1453 (
            .O(N__17475),
            .I(N__17472));
    Span4Mux_v I__1452 (
            .O(N__17472),
            .I(N__17469));
    Odrv4 I__1451 (
            .O(N__17469),
            .I(\pid_alt.un1_error_d_reg_1_20 ));
    InMux I__1450 (
            .O(N__17466),
            .I(\pid_alt.un1_error_d_reg_add_1_cry_4 ));
    InMux I__1449 (
            .O(N__17463),
            .I(N__17460));
    LocalMux I__1448 (
            .O(N__17460),
            .I(\pid_alt.un1_error_d_reg_2_6 ));
    CascadeMux I__1447 (
            .O(N__17457),
            .I(N__17454));
    InMux I__1446 (
            .O(N__17454),
            .I(N__17451));
    LocalMux I__1445 (
            .O(N__17451),
            .I(N__17448));
    Span4Mux_v I__1444 (
            .O(N__17448),
            .I(N__17445));
    Odrv4 I__1443 (
            .O(N__17445),
            .I(\pid_alt.un1_error_d_reg_1_21 ));
    InMux I__1442 (
            .O(N__17442),
            .I(\pid_alt.un1_error_d_reg_add_1_cry_5 ));
    InMux I__1441 (
            .O(N__17439),
            .I(N__17436));
    LocalMux I__1440 (
            .O(N__17436),
            .I(N__17433));
    Span4Mux_v I__1439 (
            .O(N__17433),
            .I(N__17430));
    Odrv4 I__1438 (
            .O(N__17430),
            .I(\pid_alt.un1_error_d_reg_1_22 ));
    CascadeMux I__1437 (
            .O(N__17427),
            .I(N__17424));
    InMux I__1436 (
            .O(N__17424),
            .I(N__17421));
    LocalMux I__1435 (
            .O(N__17421),
            .I(\pid_alt.un1_error_d_reg_2_7 ));
    InMux I__1434 (
            .O(N__17418),
            .I(\pid_alt.un1_error_d_reg_add_1_cry_6 ));
    InMux I__1433 (
            .O(N__17415),
            .I(N__17412));
    LocalMux I__1432 (
            .O(N__17412),
            .I(N__17409));
    Span4Mux_v I__1431 (
            .O(N__17409),
            .I(N__17406));
    Span4Mux_s1_h I__1430 (
            .O(N__17406),
            .I(N__17403));
    Odrv4 I__1429 (
            .O(N__17403),
            .I(\pid_alt.un1_error_d_reg_1_23 ));
    CascadeMux I__1428 (
            .O(N__17400),
            .I(N__17397));
    InMux I__1427 (
            .O(N__17397),
            .I(N__17394));
    LocalMux I__1426 (
            .O(N__17394),
            .I(\pid_alt.un1_error_d_reg_2_8 ));
    InMux I__1425 (
            .O(N__17391),
            .I(bfn_1_7_0_));
    CascadeMux I__1424 (
            .O(N__17388),
            .I(N__17385));
    InMux I__1423 (
            .O(N__17385),
            .I(N__17382));
    LocalMux I__1422 (
            .O(N__17382),
            .I(\pid_alt.un1_error_d_reg_2_9 ));
    InMux I__1421 (
            .O(N__17379),
            .I(\pid_alt.un1_error_d_reg_add_1_cry_8 ));
    CascadeMux I__1420 (
            .O(N__17376),
            .I(N__17373));
    InMux I__1419 (
            .O(N__17373),
            .I(N__17370));
    LocalMux I__1418 (
            .O(N__17370),
            .I(\pid_alt.un1_error_d_reg_2_10 ));
    InMux I__1417 (
            .O(N__17367),
            .I(\pid_alt.un1_error_d_reg_add_1_cry_9 ));
    CascadeMux I__1416 (
            .O(N__17364),
            .I(N__17361));
    InMux I__1415 (
            .O(N__17361),
            .I(N__17358));
    LocalMux I__1414 (
            .O(N__17358),
            .I(\pid_alt.un1_error_d_reg_2_11 ));
    InMux I__1413 (
            .O(N__17355),
            .I(N__17352));
    LocalMux I__1412 (
            .O(N__17352),
            .I(\pid_alt.un1_error_d_reg_2_1 ));
    CascadeMux I__1411 (
            .O(N__17349),
            .I(N__17346));
    InMux I__1410 (
            .O(N__17346),
            .I(N__17343));
    LocalMux I__1409 (
            .O(N__17343),
            .I(N__17340));
    Span4Mux_v I__1408 (
            .O(N__17340),
            .I(N__17337));
    Odrv4 I__1407 (
            .O(N__17337),
            .I(\pid_alt.un1_error_d_reg_1_16 ));
    InMux I__1406 (
            .O(N__17334),
            .I(\pid_alt.un1_error_d_reg_add_1_cry_0 ));
    InMux I__1405 (
            .O(N__17331),
            .I(N__17328));
    LocalMux I__1404 (
            .O(N__17328),
            .I(\pid_alt.un1_error_d_reg_2_2 ));
    CascadeMux I__1403 (
            .O(N__17325),
            .I(N__17322));
    InMux I__1402 (
            .O(N__17322),
            .I(N__17319));
    LocalMux I__1401 (
            .O(N__17319),
            .I(N__17316));
    Span4Mux_v I__1400 (
            .O(N__17316),
            .I(N__17313));
    Odrv4 I__1399 (
            .O(N__17313),
            .I(\pid_alt.un1_error_d_reg_1_17 ));
    InMux I__1398 (
            .O(N__17310),
            .I(\pid_alt.un1_error_d_reg_add_1_cry_1 ));
    InMux I__1397 (
            .O(N__17307),
            .I(N__17304));
    LocalMux I__1396 (
            .O(N__17304),
            .I(N__17301));
    Odrv4 I__1395 (
            .O(N__17301),
            .I(\pid_alt.un1_error_d_reg_2_3 ));
    CascadeMux I__1394 (
            .O(N__17298),
            .I(N__17295));
    InMux I__1393 (
            .O(N__17295),
            .I(N__17292));
    LocalMux I__1392 (
            .O(N__17292),
            .I(N__17289));
    Span4Mux_v I__1391 (
            .O(N__17289),
            .I(N__17286));
    Odrv4 I__1390 (
            .O(N__17286),
            .I(\pid_alt.un1_error_d_reg_1_18 ));
    defparam IN_MUX_bfv_7_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_13_0_));
    defparam IN_MUX_bfv_7_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_14_0_ (
            .carryinitin(\pid_alt.un1_pid_prereg_0_cry_6 ),
            .carryinitout(bfn_7_14_0_));
    defparam IN_MUX_bfv_7_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_15_0_ (
            .carryinitin(\pid_alt.un1_pid_prereg_0_cry_14 ),
            .carryinitout(bfn_7_15_0_));
    defparam IN_MUX_bfv_7_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_16_0_ (
            .carryinitin(\pid_alt.un1_pid_prereg_0_cry_22 ),
            .carryinitout(bfn_7_16_0_));
    defparam IN_MUX_bfv_11_16_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_16_0_));
    defparam IN_MUX_bfv_11_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_17_0_ (
            .carryinitin(\scaler_4.un3_source_data_0_cry_7 ),
            .carryinitout(bfn_11_17_0_));
    defparam IN_MUX_bfv_12_16_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_16_0_));
    defparam IN_MUX_bfv_12_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_17_0_ (
            .carryinitin(\scaler_4.un2_source_data_0_cry_8 ),
            .carryinitout(bfn_12_17_0_));
    defparam IN_MUX_bfv_11_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_13_0_));
    defparam IN_MUX_bfv_11_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_14_0_ (
            .carryinitin(\scaler_3.un3_source_data_0_cry_7 ),
            .carryinitout(bfn_11_14_0_));
    defparam IN_MUX_bfv_12_14_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_14_0_));
    defparam IN_MUX_bfv_12_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_15_0_ (
            .carryinitin(\scaler_3.un2_source_data_0_cry_8 ),
            .carryinitout(bfn_12_15_0_));
    defparam IN_MUX_bfv_12_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_11_0_));
    defparam IN_MUX_bfv_12_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_12_0_ (
            .carryinitin(\scaler_2.un3_source_data_0_cry_7 ),
            .carryinitout(bfn_12_12_0_));
    defparam IN_MUX_bfv_14_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_13_0_));
    defparam IN_MUX_bfv_14_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_14_0_ (
            .carryinitin(\scaler_2.un2_source_data_0_cry_8 ),
            .carryinitout(bfn_14_14_0_));
    defparam IN_MUX_bfv_16_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_7_0_));
    defparam IN_MUX_bfv_16_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_8_0_ (
            .carryinitin(\reset_module_System.count_1_cry_8 ),
            .carryinitout(bfn_16_8_0_));
    defparam IN_MUX_bfv_16_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_9_0_ (
            .carryinitin(\reset_module_System.count_1_cry_16 ),
            .carryinitout(bfn_16_9_0_));
    defparam IN_MUX_bfv_13_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_13_0_));
    defparam IN_MUX_bfv_13_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_14_0_ (
            .carryinitin(\ppm_encoder_1.un1_throttle_cry_7 ),
            .carryinitout(bfn_13_14_0_));
    defparam IN_MUX_bfv_13_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_17_0_));
    defparam IN_MUX_bfv_13_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_18_0_ (
            .carryinitin(\ppm_encoder_1.un1_rudder_cry_13 ),
            .carryinitout(bfn_13_18_0_));
    defparam IN_MUX_bfv_13_19_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_19_0_));
    defparam IN_MUX_bfv_13_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_20_0_ (
            .carryinitin(\ppm_encoder_1.un1_elevator_cry_13 ),
            .carryinitout(bfn_13_20_0_));
    defparam IN_MUX_bfv_16_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_15_0_));
    defparam IN_MUX_bfv_16_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_16_0_ (
            .carryinitin(\ppm_encoder_1.un1_aileron_cry_13 ),
            .carryinitout(bfn_16_16_0_));
    defparam IN_MUX_bfv_17_14_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_14_0_));
    defparam IN_MUX_bfv_17_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_15_0_ (
            .carryinitin(\ppm_encoder_1.un1_init_pulses_0_cry_7 ),
            .carryinitout(bfn_17_15_0_));
    defparam IN_MUX_bfv_17_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_16_0_ (
            .carryinitin(\ppm_encoder_1.un1_init_pulses_0_cry_15 ),
            .carryinitout(bfn_17_16_0_));
    defparam IN_MUX_bfv_18_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_11_0_));
    defparam IN_MUX_bfv_18_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_12_0_ (
            .carryinitin(\ppm_encoder_1.un1_init_pulses_3_cry_7 ),
            .carryinitout(bfn_18_12_0_));
    defparam IN_MUX_bfv_18_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_13_0_ (
            .carryinitin(\ppm_encoder_1.un1_init_pulses_3_cry_15 ),
            .carryinitout(bfn_18_13_0_));
    defparam IN_MUX_bfv_18_20_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_20_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_20_0_));
    defparam IN_MUX_bfv_18_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_21_0_ (
            .carryinitin(\ppm_encoder_1.counter24_0_data_tmp_7 ),
            .carryinitout(bfn_18_21_0_));
    defparam IN_MUX_bfv_8_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_11_0_));
    defparam IN_MUX_bfv_8_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_12_0_ (
            .carryinitin(\pid_alt.un9lto29_i_a2_6 ),
            .carryinitout(bfn_8_12_0_));
    defparam IN_MUX_bfv_1_6_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_6_0_));
    defparam IN_MUX_bfv_1_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_7_0_ (
            .carryinitin(\pid_alt.un1_error_d_reg_add_1_cry_7 ),
            .carryinitout(bfn_1_7_0_));
    defparam IN_MUX_bfv_1_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_8_0_ (
            .carryinitin(\pid_alt.un1_error_d_reg_add_1_cry_15 ),
            .carryinitout(bfn_1_8_0_));
    defparam IN_MUX_bfv_7_19_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_19_0_));
    defparam IN_MUX_bfv_7_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_20_0_ (
            .carryinitin(\pid_alt.error_cry_7 ),
            .carryinitout(bfn_7_20_0_));
    defparam IN_MUX_bfv_11_6_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_6_0_));
    defparam IN_MUX_bfv_15_6_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_6_0_));
    defparam IN_MUX_bfv_16_19_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_19_0_));
    defparam IN_MUX_bfv_16_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_20_0_ (
            .carryinitin(\ppm_encoder_1.un1_counter_13_cry_7 ),
            .carryinitout(bfn_16_20_0_));
    defparam IN_MUX_bfv_16_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_21_0_ (
            .carryinitin(\ppm_encoder_1.un1_counter_13_cry_15 ),
            .carryinitout(bfn_16_21_0_));
    defparam IN_MUX_bfv_17_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_17_0_));
    defparam IN_MUX_bfv_17_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_18_0_ (
            .carryinitin(\pid_alt.un9_error_filt_add_1_cry_7 ),
            .carryinitout(bfn_17_18_0_));
    defparam IN_MUX_bfv_13_21_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_21_0_));
    defparam IN_MUX_bfv_13_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_22_0_ (
            .carryinitin(\pid_alt.un1_error_i_acumm_prereg_cry_7 ),
            .carryinitout(bfn_13_22_0_));
    defparam IN_MUX_bfv_13_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_23_0_ (
            .carryinitin(\pid_alt.un1_error_i_acumm_prereg_cry_15 ),
            .carryinitout(bfn_13_23_0_));
    defparam IN_MUX_bfv_1_16_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_16_0_));
    defparam IN_MUX_bfv_1_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_17_0_ (
            .carryinitin(\pid_alt.error_filt_cry_7 ),
            .carryinitout(bfn_1_17_0_));
    defparam IN_MUX_bfv_1_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_18_0_ (
            .carryinitin(\pid_alt.error_filt_cry_15 ),
            .carryinitout(bfn_1_18_0_));
    defparam IN_MUX_bfv_7_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_7_0_));
    defparam IN_MUX_bfv_7_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_8_0_ (
            .carryinitin(\dron_frame_decoder_1.un1_WDT_cry_7 ),
            .carryinitout(bfn_7_8_0_));
    defparam IN_MUX_bfv_9_5_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_5_0_));
    defparam IN_MUX_bfv_9_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_6_0_ (
            .carryinitin(\Commands_frame_decoder.un1_WDT_cry_7 ),
            .carryinitout(bfn_9_6_0_));
    ICE_GB \reset_module_System.reset_RNITC69_0  (
            .USERSIGNALTOGLOBALBUFFER(N__43371),
            .GLOBALBUFFEROUTPUT(N_411_g));
    ICE_GB \reset_module_System.reset_RNITC69  (
            .USERSIGNALTOGLOBALBUFFER(N__32938),
            .GLOBALBUFFEROUTPUT(reset_system_g));
    ICE_GB \pid_alt.state_RNICP2N1_0_0  (
            .USERSIGNALTOGLOBALBUFFER(N__22293),
            .GLOBALBUFFEROUTPUT(\pid_alt.N_410_0_g ));
    ICE_GB debug_CH3_20A_c_0_g_gb (
            .USERSIGNALTOGLOBALBUFFER(N__30507),
            .GLOBALBUFFEROUTPUT(debug_CH3_20A_c_0_g));
    ICE_GB \pid_alt.state_RNIH1EN_0_0  (
            .USERSIGNALTOGLOBALBUFFER(N__24912),
            .GLOBALBUFFEROUTPUT(\pid_alt.state_0_g_0 ));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    ICE_GB \ppm_encoder_1.counter24_0_I_57_c_RNIGCO83_0  (
            .USERSIGNALTOGLOBALBUFFER(N__32886),
            .GLOBALBUFFEROUTPUT(\ppm_encoder_1.N_322_g ));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \pid_alt.un1_error_d_reg_add_1_cry_0_c_LC_1_6_0 .C_ON=1'b1;
    defparam \pid_alt.un1_error_d_reg_add_1_cry_0_c_LC_1_6_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un1_error_d_reg_add_1_cry_0_c_LC_1_6_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_alt.un1_error_d_reg_add_1_cry_0_c_LC_1_6_0  (
            .in0(_gnd_net_),
            .in1(N__17549),
            .in2(N__17538),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_6_0_),
            .carryout(\pid_alt.un1_error_d_reg_add_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_esr_12_LC_1_6_1 .C_ON=1'b1;
    defparam \pid_alt.error_d_reg_esr_12_LC_1_6_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_12_LC_1_6_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_d_reg_esr_12_LC_1_6_1  (
            .in0(_gnd_net_),
            .in1(N__17355),
            .in2(N__17349),
            .in3(N__17334),
            .lcout(\pid_alt.error_d_regZ0Z_12 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_d_reg_add_1_cry_0 ),
            .carryout(\pid_alt.un1_error_d_reg_add_1_cry_1 ),
            .clk(N__47478),
            .ce(N__46815),
            .sr(N__46628));
    defparam \pid_alt.error_d_reg_esr_13_LC_1_6_2 .C_ON=1'b1;
    defparam \pid_alt.error_d_reg_esr_13_LC_1_6_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_13_LC_1_6_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_d_reg_esr_13_LC_1_6_2  (
            .in0(_gnd_net_),
            .in1(N__17331),
            .in2(N__17325),
            .in3(N__17310),
            .lcout(\pid_alt.error_d_regZ0Z_13 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_d_reg_add_1_cry_1 ),
            .carryout(\pid_alt.un1_error_d_reg_add_1_cry_2 ),
            .clk(N__47478),
            .ce(N__46815),
            .sr(N__46628));
    defparam \pid_alt.error_d_reg_esr_14_LC_1_6_3 .C_ON=1'b1;
    defparam \pid_alt.error_d_reg_esr_14_LC_1_6_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_14_LC_1_6_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_d_reg_esr_14_LC_1_6_3  (
            .in0(_gnd_net_),
            .in1(N__17307),
            .in2(N__17298),
            .in3(N__17517),
            .lcout(\pid_alt.error_d_regZ0Z_14 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_d_reg_add_1_cry_2 ),
            .carryout(\pid_alt.un1_error_d_reg_add_1_cry_3 ),
            .clk(N__47478),
            .ce(N__46815),
            .sr(N__46628));
    defparam \pid_alt.error_d_reg_esr_15_LC_1_6_4 .C_ON=1'b1;
    defparam \pid_alt.error_d_reg_esr_15_LC_1_6_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_15_LC_1_6_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_d_reg_esr_15_LC_1_6_4  (
            .in0(_gnd_net_),
            .in1(N__17514),
            .in2(N__17505),
            .in3(N__17490),
            .lcout(\pid_alt.error_d_regZ0Z_15 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_d_reg_add_1_cry_3 ),
            .carryout(\pid_alt.un1_error_d_reg_add_1_cry_4 ),
            .clk(N__47478),
            .ce(N__46815),
            .sr(N__46628));
    defparam \pid_alt.error_d_reg_esr_16_LC_1_6_5 .C_ON=1'b1;
    defparam \pid_alt.error_d_reg_esr_16_LC_1_6_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_16_LC_1_6_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_d_reg_esr_16_LC_1_6_5  (
            .in0(_gnd_net_),
            .in1(N__17487),
            .in2(N__17481),
            .in3(N__17466),
            .lcout(\pid_alt.error_d_regZ0Z_16 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_d_reg_add_1_cry_4 ),
            .carryout(\pid_alt.un1_error_d_reg_add_1_cry_5 ),
            .clk(N__47478),
            .ce(N__46815),
            .sr(N__46628));
    defparam \pid_alt.error_d_reg_esr_17_LC_1_6_6 .C_ON=1'b1;
    defparam \pid_alt.error_d_reg_esr_17_LC_1_6_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_17_LC_1_6_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_d_reg_esr_17_LC_1_6_6  (
            .in0(_gnd_net_),
            .in1(N__17463),
            .in2(N__17457),
            .in3(N__17442),
            .lcout(\pid_alt.error_d_regZ0Z_17 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_d_reg_add_1_cry_5 ),
            .carryout(\pid_alt.un1_error_d_reg_add_1_cry_6 ),
            .clk(N__47478),
            .ce(N__46815),
            .sr(N__46628));
    defparam \pid_alt.error_d_reg_esr_18_LC_1_6_7 .C_ON=1'b1;
    defparam \pid_alt.error_d_reg_esr_18_LC_1_6_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_18_LC_1_6_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_d_reg_esr_18_LC_1_6_7  (
            .in0(_gnd_net_),
            .in1(N__17439),
            .in2(N__17427),
            .in3(N__17418),
            .lcout(\pid_alt.error_d_regZ0Z_18 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_d_reg_add_1_cry_6 ),
            .carryout(\pid_alt.un1_error_d_reg_add_1_cry_7 ),
            .clk(N__47478),
            .ce(N__46815),
            .sr(N__46628));
    defparam \pid_alt.error_d_reg_esr_19_LC_1_7_0 .C_ON=1'b1;
    defparam \pid_alt.error_d_reg_esr_19_LC_1_7_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_19_LC_1_7_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_d_reg_esr_19_LC_1_7_0  (
            .in0(_gnd_net_),
            .in1(N__17415),
            .in2(N__17400),
            .in3(N__17391),
            .lcout(\pid_alt.error_d_regZ0Z_19 ),
            .ltout(),
            .carryin(bfn_1_7_0_),
            .carryout(\pid_alt.un1_error_d_reg_add_1_cry_8 ),
            .clk(N__47477),
            .ce(N__46814),
            .sr(N__46627));
    defparam \pid_alt.error_d_reg_esr_20_LC_1_7_1 .C_ON=1'b1;
    defparam \pid_alt.error_d_reg_esr_20_LC_1_7_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_20_LC_1_7_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_d_reg_esr_20_LC_1_7_1  (
            .in0(_gnd_net_),
            .in1(N__17615),
            .in2(N__17388),
            .in3(N__17379),
            .lcout(\pid_alt.error_d_regZ0Z_20 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_d_reg_add_1_cry_8 ),
            .carryout(\pid_alt.un1_error_d_reg_add_1_cry_9 ),
            .clk(N__47477),
            .ce(N__46814),
            .sr(N__46627));
    defparam \pid_alt.error_d_reg_esr_21_LC_1_7_2 .C_ON=1'b1;
    defparam \pid_alt.error_d_reg_esr_21_LC_1_7_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_21_LC_1_7_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_d_reg_esr_21_LC_1_7_2  (
            .in0(_gnd_net_),
            .in1(N__17619),
            .in2(N__17376),
            .in3(N__17367),
            .lcout(\pid_alt.error_d_regZ0Z_21 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_d_reg_add_1_cry_9 ),
            .carryout(\pid_alt.un1_error_d_reg_add_1_cry_10 ),
            .clk(N__47477),
            .ce(N__46814),
            .sr(N__46627));
    defparam \pid_alt.error_d_reg_esr_22_LC_1_7_3 .C_ON=1'b1;
    defparam \pid_alt.error_d_reg_esr_22_LC_1_7_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_22_LC_1_7_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_d_reg_esr_22_LC_1_7_3  (
            .in0(_gnd_net_),
            .in1(N__17616),
            .in2(N__17364),
            .in3(N__17673),
            .lcout(\pid_alt.error_d_regZ0Z_22 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_d_reg_add_1_cry_10 ),
            .carryout(\pid_alt.un1_error_d_reg_add_1_cry_11 ),
            .clk(N__47477),
            .ce(N__46814),
            .sr(N__46627));
    defparam \pid_alt.error_d_reg_esr_23_LC_1_7_4 .C_ON=1'b1;
    defparam \pid_alt.error_d_reg_esr_23_LC_1_7_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_23_LC_1_7_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_d_reg_esr_23_LC_1_7_4  (
            .in0(_gnd_net_),
            .in1(N__17620),
            .in2(N__17670),
            .in3(N__17661),
            .lcout(\pid_alt.error_d_regZ0Z_23 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_d_reg_add_1_cry_11 ),
            .carryout(\pid_alt.un1_error_d_reg_add_1_cry_12 ),
            .clk(N__47477),
            .ce(N__46814),
            .sr(N__46627));
    defparam \pid_alt.error_d_reg_esr_24_LC_1_7_5 .C_ON=1'b1;
    defparam \pid_alt.error_d_reg_esr_24_LC_1_7_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_24_LC_1_7_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_d_reg_esr_24_LC_1_7_5  (
            .in0(_gnd_net_),
            .in1(N__17617),
            .in2(N__17658),
            .in3(N__17649),
            .lcout(\pid_alt.error_d_regZ0Z_24 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_d_reg_add_1_cry_12 ),
            .carryout(\pid_alt.un1_error_d_reg_add_1_cry_13 ),
            .clk(N__47477),
            .ce(N__46814),
            .sr(N__46627));
    defparam \pid_alt.error_d_reg_esr_25_LC_1_7_6 .C_ON=1'b1;
    defparam \pid_alt.error_d_reg_esr_25_LC_1_7_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_25_LC_1_7_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_d_reg_esr_25_LC_1_7_6  (
            .in0(_gnd_net_),
            .in1(N__17621),
            .in2(N__17646),
            .in3(N__17637),
            .lcout(\pid_alt.error_d_regZ0Z_25 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_d_reg_add_1_cry_13 ),
            .carryout(\pid_alt.un1_error_d_reg_add_1_cry_14 ),
            .clk(N__47477),
            .ce(N__46814),
            .sr(N__46627));
    defparam \pid_alt.error_d_reg_esr_26_LC_1_7_7 .C_ON=1'b1;
    defparam \pid_alt.error_d_reg_esr_26_LC_1_7_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_26_LC_1_7_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_d_reg_esr_26_LC_1_7_7  (
            .in0(_gnd_net_),
            .in1(N__17618),
            .in2(N__17634),
            .in3(N__17625),
            .lcout(\pid_alt.error_d_regZ0Z_26 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_d_reg_add_1_cry_14 ),
            .carryout(\pid_alt.un1_error_d_reg_add_1_cry_15 ),
            .clk(N__47477),
            .ce(N__46814),
            .sr(N__46627));
    defparam \pid_alt.error_d_reg_esr_27_LC_1_8_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_27_LC_1_8_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_27_LC_1_8_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_d_reg_esr_27_LC_1_8_0  (
            .in0(_gnd_net_),
            .in1(N__17622),
            .in2(N__17577),
            .in3(N__17568),
            .lcout(\pid_alt.error_d_regZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47476),
            .ce(N__46812),
            .sr(N__46626));
    defparam \pid_alt.error_d_reg_esr_6_LC_1_8_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_6_LC_1_8_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_6_LC_1_8_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_6_LC_1_8_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17565),
            .lcout(\pid_alt.error_d_regZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47476),
            .ce(N__46812),
            .sr(N__46626));
    defparam \pid_alt.error_d_reg_11_LC_1_9_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_11_LC_1_9_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_11_LC_1_9_0 .LUT_INIT=16'b0111001011011000;
    LogicCell40 \pid_alt.error_d_reg_11_LC_1_9_0  (
            .in0(N__24128),
            .in1(N__17556),
            .in2(N__19664),
            .in3(N__17534),
            .lcout(\pid_alt.error_d_regZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47472),
            .ce(),
            .sr(N__46625));
    defparam \pid_alt.error_d_reg_prev_esr_RNI20IM_17_LC_1_9_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI20IM_17_LC_1_9_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI20IM_17_LC_1_9_7 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI20IM_17_LC_1_9_7  (
            .in0(N__18500),
            .in1(N__18474),
            .in2(_gnd_net_),
            .in3(N__18461),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI20IMZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_esr_9_LC_1_10_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_9_LC_1_10_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_9_LC_1_10_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_9_LC_1_10_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17730),
            .lcout(\pid_alt.error_d_regZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47470),
            .ce(N__46809),
            .sr(N__46624));
    defparam \pid_alt.error_d_reg_esr_7_LC_1_10_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_7_LC_1_10_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_7_LC_1_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_7_LC_1_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17724),
            .lcout(\pid_alt.error_d_regZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47470),
            .ce(N__46809),
            .sr(N__46624));
    defparam \pid_alt.error_d_reg_esr_1_LC_1_11_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_1_LC_1_11_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_1_LC_1_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_1_LC_1_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17714),
            .lcout(\pid_alt.error_d_regZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47464),
            .ce(N__46805),
            .sr(N__46623));
    defparam \pid_alt.error_d_reg_fast_esr_1_LC_1_11_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_fast_esr_1_LC_1_11_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_fast_esr_1_LC_1_11_2 .LUT_INIT=16'b1111000011110000;
    LogicCell40 \pid_alt.error_d_reg_fast_esr_1_LC_1_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17718),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_d_reg_fastZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47464),
            .ce(N__46805),
            .sr(N__46623));
    defparam \pid_alt.error_d_reg_esr_10_LC_1_11_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_10_LC_1_11_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_10_LC_1_11_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_10_LC_1_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17706),
            .lcout(\pid_alt.error_d_regZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47464),
            .ce(N__46805),
            .sr(N__46623));
    defparam \pid_alt.error_d_reg_esr_2_LC_1_11_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_2_LC_1_11_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_2_LC_1_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_2_LC_1_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17700),
            .lcout(\pid_alt.error_d_regZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47464),
            .ce(N__46805),
            .sr(N__46623));
    defparam \pid_alt.error_d_reg_esr_8_LC_1_11_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_8_LC_1_11_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_8_LC_1_11_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_8_LC_1_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17694),
            .lcout(\pid_alt.error_d_regZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47464),
            .ce(N__46805),
            .sr(N__46623));
    defparam \pid_alt.error_d_reg_esr_5_LC_1_11_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_5_LC_1_11_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_5_LC_1_11_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_5_LC_1_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17688),
            .lcout(\pid_alt.error_d_regZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47464),
            .ce(N__46805),
            .sr(N__46623));
    defparam \pid_alt.error_d_reg_esr_3_LC_1_12_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_3_LC_1_12_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_3_LC_1_12_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_3_LC_1_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17682),
            .lcout(\pid_alt.error_d_regZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47459),
            .ce(N__46801),
            .sr(N__46621));
    defparam \pid_alt.error_d_reg_prev_esr_2_LC_1_13_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_2_LC_1_13_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_2_LC_1_13_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_2_LC_1_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19249),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47452),
            .ce(N__33622),
            .sr(N__43831));
    defparam \pid_alt.error_p_reg_esr_0_LC_1_15_3 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_0_LC_1_15_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_0_LC_1_15_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_0_LC_1_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17970),
            .lcout(\pid_alt.error_p_regZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47438),
            .ce(N__46800),
            .sr(N__46620));
    defparam \pid_alt.error_filt_prev_esr_0_LC_1_15_7 .C_ON=1'b0;
    defparam \pid_alt.error_filt_prev_esr_0_LC_1_15_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_filt_prev_esr_0_LC_1_15_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_alt.error_filt_prev_esr_0_LC_1_15_7  (
            .in0(_gnd_net_),
            .in1(N__17930),
            .in2(_gnd_net_),
            .in3(N__17897),
            .lcout(\pid_alt.error_filt_prevZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47438),
            .ce(N__46800),
            .sr(N__46620));
    defparam \pid_alt.error_filt_error_filt_axb_0_LC_1_16_0 .C_ON=1'b1;
    defparam \pid_alt.error_filt_error_filt_axb_0_LC_1_16_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_filt_error_filt_axb_0_LC_1_16_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \pid_alt.error_filt_error_filt_axb_0_LC_1_16_0  (
            .in0(_gnd_net_),
            .in1(N__17931),
            .in2(N__17898),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_filt_0 ),
            .ltout(),
            .carryin(bfn_1_16_0_),
            .carryout(\pid_alt.error_filt_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_filt_error_filt_cry_0_c_RNIBLFT_LC_1_16_1 .C_ON=1'b1;
    defparam \pid_alt.error_filt_error_filt_cry_0_c_RNIBLFT_LC_1_16_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_filt_error_filt_cry_0_c_RNIBLFT_LC_1_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_filt_error_filt_cry_0_c_RNIBLFT_LC_1_16_1  (
            .in0(_gnd_net_),
            .in1(N__17871),
            .in2(N__17853),
            .in3(N__17844),
            .lcout(\pid_alt.error_filt_1 ),
            .ltout(),
            .carryin(\pid_alt.error_filt_cry_0 ),
            .carryout(\pid_alt.error_filt_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_filt_error_filt_cry_1_c_RNICNGT_LC_1_16_2 .C_ON=1'b1;
    defparam \pid_alt.error_filt_error_filt_cry_1_c_RNICNGT_LC_1_16_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_filt_error_filt_cry_1_c_RNICNGT_LC_1_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_filt_error_filt_cry_1_c_RNICNGT_LC_1_16_2  (
            .in0(_gnd_net_),
            .in1(N__17841),
            .in2(N__17823),
            .in3(N__17814),
            .lcout(\pid_alt.error_filt_2 ),
            .ltout(),
            .carryin(\pid_alt.error_filt_cry_1 ),
            .carryout(\pid_alt.error_filt_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_filt_error_filt_cry_2_c_RNIDPHT_LC_1_16_3 .C_ON=1'b1;
    defparam \pid_alt.error_filt_error_filt_cry_2_c_RNIDPHT_LC_1_16_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_filt_error_filt_cry_2_c_RNIDPHT_LC_1_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_filt_error_filt_cry_2_c_RNIDPHT_LC_1_16_3  (
            .in0(_gnd_net_),
            .in1(N__17811),
            .in2(N__17796),
            .in3(N__17787),
            .lcout(\pid_alt.error_filt_3 ),
            .ltout(),
            .carryin(\pid_alt.error_filt_cry_2 ),
            .carryout(\pid_alt.error_filt_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_filt_error_filt_cry_3_c_RNIERIT_LC_1_16_4 .C_ON=1'b1;
    defparam \pid_alt.error_filt_error_filt_cry_3_c_RNIERIT_LC_1_16_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_filt_error_filt_cry_3_c_RNIERIT_LC_1_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_filt_error_filt_cry_3_c_RNIERIT_LC_1_16_4  (
            .in0(_gnd_net_),
            .in1(N__17784),
            .in2(N__17766),
            .in3(N__17757),
            .lcout(\pid_alt.error_filt_4 ),
            .ltout(),
            .carryin(\pid_alt.error_filt_cry_3 ),
            .carryout(\pid_alt.error_filt_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_filt_error_filt_cry_4_c_RNIFTJT_LC_1_16_5 .C_ON=1'b1;
    defparam \pid_alt.error_filt_error_filt_cry_4_c_RNIFTJT_LC_1_16_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_filt_error_filt_cry_4_c_RNIFTJT_LC_1_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_filt_error_filt_cry_4_c_RNIFTJT_LC_1_16_5  (
            .in0(_gnd_net_),
            .in1(N__17754),
            .in2(N__17748),
            .in3(N__18150),
            .lcout(\pid_alt.error_filt_5 ),
            .ltout(),
            .carryin(\pid_alt.error_filt_cry_4 ),
            .carryout(\pid_alt.error_filt_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_filt_error_filt_cry_5_c_RNIGVKT_LC_1_16_6 .C_ON=1'b1;
    defparam \pid_alt.error_filt_error_filt_cry_5_c_RNIGVKT_LC_1_16_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_filt_error_filt_cry_5_c_RNIGVKT_LC_1_16_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_filt_error_filt_cry_5_c_RNIGVKT_LC_1_16_6  (
            .in0(_gnd_net_),
            .in1(N__18147),
            .in2(N__18120),
            .in3(N__18111),
            .lcout(\pid_alt.error_filt_6 ),
            .ltout(),
            .carryin(\pid_alt.error_filt_cry_5 ),
            .carryout(\pid_alt.error_filt_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_filt_error_filt_cry_6_c_RNIH1MT_LC_1_16_7 .C_ON=1'b1;
    defparam \pid_alt.error_filt_error_filt_cry_6_c_RNIH1MT_LC_1_16_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_filt_error_filt_cry_6_c_RNIH1MT_LC_1_16_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_filt_error_filt_cry_6_c_RNIH1MT_LC_1_16_7  (
            .in0(_gnd_net_),
            .in1(N__18108),
            .in2(N__18102),
            .in3(N__18081),
            .lcout(\pid_alt.error_filt_7 ),
            .ltout(),
            .carryin(\pid_alt.error_filt_cry_6 ),
            .carryout(\pid_alt.error_filt_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_filt_error_filt_cry_7_c_RNII3NT_LC_1_17_0 .C_ON=1'b1;
    defparam \pid_alt.error_filt_error_filt_cry_7_c_RNII3NT_LC_1_17_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_filt_error_filt_cry_7_c_RNII3NT_LC_1_17_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_filt_error_filt_cry_7_c_RNII3NT_LC_1_17_0  (
            .in0(_gnd_net_),
            .in1(N__18078),
            .in2(N__18060),
            .in3(N__18051),
            .lcout(\pid_alt.error_filt_8 ),
            .ltout(),
            .carryin(bfn_1_17_0_),
            .carryout(\pid_alt.error_filt_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_filt_error_filt_cry_8_c_RNIJ5OT_LC_1_17_1 .C_ON=1'b1;
    defparam \pid_alt.error_filt_error_filt_cry_8_c_RNIJ5OT_LC_1_17_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_filt_error_filt_cry_8_c_RNIJ5OT_LC_1_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_filt_error_filt_cry_8_c_RNIJ5OT_LC_1_17_1  (
            .in0(_gnd_net_),
            .in1(N__18048),
            .in2(N__18030),
            .in3(N__18021),
            .lcout(\pid_alt.error_filt_9 ),
            .ltout(),
            .carryin(\pid_alt.error_filt_cry_8 ),
            .carryout(\pid_alt.error_filt_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un9_error_filt_add_1_axb_0_RNIRHEM_LC_1_17_2 .C_ON=1'b1;
    defparam \pid_alt.un9_error_filt_add_1_axb_0_RNIRHEM_LC_1_17_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un9_error_filt_add_1_axb_0_RNIRHEM_LC_1_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.un9_error_filt_add_1_axb_0_RNIRHEM_LC_1_17_2  (
            .in0(_gnd_net_),
            .in1(N__38310),
            .in2(N__18018),
            .in3(N__18009),
            .lcout(\pid_alt.error_filt_10 ),
            .ltout(),
            .carryin(\pid_alt.error_filt_cry_9 ),
            .carryout(\pid_alt.error_filt_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un9_error_filt_add_1_cry_1_s_RNI9PB01_LC_1_17_3 .C_ON=1'b1;
    defparam \pid_alt.un9_error_filt_add_1_cry_1_s_RNI9PB01_LC_1_17_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un9_error_filt_add_1_cry_1_s_RNI9PB01_LC_1_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.un9_error_filt_add_1_cry_1_s_RNI9PB01_LC_1_17_3  (
            .in0(_gnd_net_),
            .in1(N__38250),
            .in2(N__18006),
            .in3(N__17997),
            .lcout(\pid_alt.error_filt_11 ),
            .ltout(),
            .carryin(\pid_alt.error_filt_cry_10 ),
            .carryout(\pid_alt.error_filt_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un9_error_filt_add_1_cry_2_s_RNIBTD01_LC_1_17_4 .C_ON=1'b1;
    defparam \pid_alt.un9_error_filt_add_1_cry_2_s_RNIBTD01_LC_1_17_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un9_error_filt_add_1_cry_2_s_RNIBTD01_LC_1_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.un9_error_filt_add_1_cry_2_s_RNIBTD01_LC_1_17_4  (
            .in0(_gnd_net_),
            .in1(N__38739),
            .in2(N__17994),
            .in3(N__17985),
            .lcout(\pid_alt.error_filt_12 ),
            .ltout(),
            .carryin(\pid_alt.error_filt_cry_11 ),
            .carryout(\pid_alt.error_filt_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un9_error_filt_add_1_cry_3_s_RNID1G01_LC_1_17_5 .C_ON=1'b1;
    defparam \pid_alt.un9_error_filt_add_1_cry_3_s_RNID1G01_LC_1_17_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un9_error_filt_add_1_cry_3_s_RNID1G01_LC_1_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.un9_error_filt_add_1_cry_3_s_RNID1G01_LC_1_17_5  (
            .in0(_gnd_net_),
            .in1(N__38679),
            .in2(N__17982),
            .in3(N__17973),
            .lcout(\pid_alt.error_filt_13 ),
            .ltout(),
            .carryin(\pid_alt.error_filt_cry_12 ),
            .carryout(\pid_alt.error_filt_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un9_error_filt_add_1_cry_4_s_RNIF5I01_LC_1_17_6 .C_ON=1'b1;
    defparam \pid_alt.un9_error_filt_add_1_cry_4_s_RNIF5I01_LC_1_17_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un9_error_filt_add_1_cry_4_s_RNIF5I01_LC_1_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.un9_error_filt_add_1_cry_4_s_RNIF5I01_LC_1_17_6  (
            .in0(_gnd_net_),
            .in1(N__18189),
            .in2(N__38640),
            .in3(N__18183),
            .lcout(\pid_alt.error_filt_14 ),
            .ltout(),
            .carryin(\pid_alt.error_filt_cry_13 ),
            .carryout(\pid_alt.error_filt_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un9_error_filt_add_1_cry_5_s_RNIH9K01_LC_1_17_7 .C_ON=1'b1;
    defparam \pid_alt.un9_error_filt_add_1_cry_5_s_RNIH9K01_LC_1_17_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un9_error_filt_add_1_cry_5_s_RNIH9K01_LC_1_17_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.un9_error_filt_add_1_cry_5_s_RNIH9K01_LC_1_17_7  (
            .in0(_gnd_net_),
            .in1(N__38604),
            .in2(N__18180),
            .in3(N__18171),
            .lcout(\pid_alt.error_filt_15 ),
            .ltout(),
            .carryin(\pid_alt.error_filt_cry_14 ),
            .carryout(\pid_alt.error_filt_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un9_error_filt_add_1_cry_6_s_RNIJDM01_LC_1_18_0 .C_ON=1'b1;
    defparam \pid_alt.un9_error_filt_add_1_cry_6_s_RNIJDM01_LC_1_18_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un9_error_filt_add_1_cry_6_s_RNIJDM01_LC_1_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.un9_error_filt_add_1_cry_6_s_RNIJDM01_LC_1_18_0  (
            .in0(_gnd_net_),
            .in1(N__38568),
            .in2(N__18316),
            .in3(N__18168),
            .lcout(\pid_alt.error_filt_16 ),
            .ltout(),
            .carryin(bfn_1_18_0_),
            .carryout(\pid_alt.error_filt_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un9_error_filt_add_1_cry_7_s_RNILHO01_LC_1_18_1 .C_ON=1'b1;
    defparam \pid_alt.un9_error_filt_add_1_cry_7_s_RNILHO01_LC_1_18_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un9_error_filt_add_1_cry_7_s_RNILHO01_LC_1_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.un9_error_filt_add_1_cry_7_s_RNILHO01_LC_1_18_1  (
            .in0(_gnd_net_),
            .in1(N__18306),
            .in2(N__38526),
            .in3(N__18165),
            .lcout(\pid_alt.error_filt_17 ),
            .ltout(),
            .carryin(\pid_alt.error_filt_cry_16 ),
            .carryout(\pid_alt.error_filt_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un9_error_filt_add_1_cry_8_s_RNINLQ01_LC_1_18_2 .C_ON=1'b1;
    defparam \pid_alt.un9_error_filt_add_1_cry_8_s_RNINLQ01_LC_1_18_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un9_error_filt_add_1_cry_8_s_RNINLQ01_LC_1_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.un9_error_filt_add_1_cry_8_s_RNINLQ01_LC_1_18_2  (
            .in0(_gnd_net_),
            .in1(N__38475),
            .in2(N__18317),
            .in3(N__18162),
            .lcout(\pid_alt.error_filt_18 ),
            .ltout(),
            .carryin(\pid_alt.error_filt_cry_17 ),
            .carryout(\pid_alt.error_filt_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un9_error_filt_add_1_cry_9_s_RNIPPS01_LC_1_18_3 .C_ON=1'b1;
    defparam \pid_alt.un9_error_filt_add_1_cry_9_s_RNIPPS01_LC_1_18_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un9_error_filt_add_1_cry_9_s_RNIPPS01_LC_1_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.un9_error_filt_add_1_cry_9_s_RNIPPS01_LC_1_18_3  (
            .in0(_gnd_net_),
            .in1(N__18310),
            .in2(N__39195),
            .in3(N__18159),
            .lcout(\pid_alt.error_filt_19 ),
            .ltout(),
            .carryin(\pid_alt.error_filt_cry_18 ),
            .carryout(\pid_alt.error_filt_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un9_error_filt_add_1_cry_10_s_RNI20BR_LC_1_18_4 .C_ON=1'b1;
    defparam \pid_alt.un9_error_filt_add_1_cry_10_s_RNI20BR_LC_1_18_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un9_error_filt_add_1_cry_10_s_RNI20BR_LC_1_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.un9_error_filt_add_1_cry_10_s_RNI20BR_LC_1_18_4  (
            .in0(_gnd_net_),
            .in1(N__39156),
            .in2(N__18318),
            .in3(N__18156),
            .lcout(\pid_alt.error_filt_20 ),
            .ltout(),
            .carryin(\pid_alt.error_filt_cry_19 ),
            .carryout(\pid_alt.error_filt_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_filt_error_filt_cry_20_c_RNIEB1O_LC_1_18_5 .C_ON=1'b1;
    defparam \pid_alt.error_filt_error_filt_cry_20_c_RNIEB1O_LC_1_18_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_filt_error_filt_cry_20_c_RNIEB1O_LC_1_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_filt_error_filt_cry_20_c_RNIEB1O_LC_1_18_5  (
            .in0(_gnd_net_),
            .in1(N__18314),
            .in2(N__39060),
            .in3(N__18153),
            .lcout(\pid_alt.error_filt_21 ),
            .ltout(),
            .carryin(\pid_alt.error_filt_cry_20 ),
            .carryout(\pid_alt.error_filt_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_filt_error_filt_cry_21_c_RNIFD2O_LC_1_18_6 .C_ON=1'b0;
    defparam \pid_alt.error_filt_error_filt_cry_21_c_RNIFD2O_LC_1_18_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_filt_error_filt_cry_21_c_RNIFD2O_LC_1_18_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_filt_error_filt_cry_21_c_RNIFD2O_LC_1_18_6  (
            .in0(N__18315),
            .in1(N__39059),
            .in2(_gnd_net_),
            .in3(N__18285),
            .lcout(\pid_alt.error_filt_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_p_reg_esr_7_LC_1_19_2 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_7_LC_1_19_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_7_LC_1_19_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_7_LC_1_19_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18282),
            .lcout(\pid_alt.error_p_regZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47393),
            .ce(N__46793),
            .sr(N__46616));
    defparam \pid_alt.error_p_reg_esr_8_LC_1_20_4 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_8_LC_1_20_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_8_LC_1_20_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_8_LC_1_20_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18270),
            .lcout(\pid_alt.error_p_regZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47378),
            .ce(N__46791),
            .sr(N__46614));
    defparam \pid_alt.error_p_reg_esr_6_LC_1_21_2 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_6_LC_1_21_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_6_LC_1_21_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_6_LC_1_21_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18258),
            .lcout(\pid_alt.error_p_regZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47366),
            .ce(N__46790),
            .sr(N__46613));
    defparam \pid_alt.error_p_reg_esr_13_LC_1_21_4 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_13_LC_1_21_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_13_LC_1_21_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_13_LC_1_21_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18249),
            .lcout(\pid_alt.error_p_regZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47366),
            .ce(N__46790),
            .sr(N__46613));
    defparam \pid_alt.error_p_reg_esr_16_LC_1_22_3 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_16_LC_1_22_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_16_LC_1_22_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_16_LC_1_22_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18237),
            .lcout(\pid_alt.error_p_regZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47352),
            .ce(N__46789),
            .sr(N__46612));
    defparam \pid_alt.error_p_reg_esr_19_LC_1_22_4 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_19_LC_1_22_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_19_LC_1_22_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_19_LC_1_22_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18228),
            .lcout(\pid_alt.error_p_regZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47352),
            .ce(N__46789),
            .sr(N__46612));
    defparam \pid_alt.error_p_reg_esr_9_LC_1_22_6 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_9_LC_1_22_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_9_LC_1_22_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_9_LC_1_22_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18216),
            .lcout(\pid_alt.error_p_regZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47352),
            .ce(N__46789),
            .sr(N__46612));
    defparam \pid_alt.error_p_reg_esr_17_LC_1_23_1 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_17_LC_1_23_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_17_LC_1_23_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_17_LC_1_23_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18207),
            .lcout(\pid_alt.error_p_regZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47336),
            .ce(N__46788),
            .sr(N__46610));
    defparam \pid_alt.error_p_reg_esr_20_LC_1_23_4 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_20_LC_1_23_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_20_LC_1_23_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_20_LC_1_23_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18198),
            .lcout(\pid_alt.error_p_regZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47336),
            .ce(N__46788),
            .sr(N__46610));
    defparam \pid_alt.error_p_reg_esr_14_LC_1_23_6 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_14_LC_1_23_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_14_LC_1_23_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_14_LC_1_23_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18519),
            .lcout(\pid_alt.error_p_regZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47336),
            .ce(N__46788),
            .sr(N__46610));
    defparam \pid_alt.error_p_reg_esr_15_LC_1_24_3 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_15_LC_1_24_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_15_LC_1_24_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_15_LC_1_24_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18510),
            .lcout(\pid_alt.error_p_regZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47323),
            .ce(N__46785),
            .sr(N__46606));
    defparam \pid_alt.error_d_reg_prev_esr_17_LC_2_8_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_17_LC_2_8_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_17_LC_2_8_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_17_LC_2_8_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18462),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47474),
            .ce(N__33599),
            .sr(N__43803));
    defparam \pid_alt.error_d_reg_prev_esr_RNI20IM_0_17_LC_2_9_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI20IM_0_17_LC_2_9_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI20IM_0_17_LC_2_9_6 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI20IM_0_17_LC_2_9_6  (
            .in0(N__18504),
            .in1(N__18473),
            .in2(_gnd_net_),
            .in3(N__18460),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI20IM_0Z0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kd_2_LC_2_10_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kd_2_LC_2_10_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kd_2_LC_2_10_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Commands_frame_decoder.source_alt_kd_2_LC_2_10_2  (
            .in0(N__36871),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(alt_kd_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47467),
            .ce(N__18972),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kd_3_LC_2_10_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kd_3_LC_2_10_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kd_3_LC_2_10_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_alt_kd_3_LC_2_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43353),
            .lcout(alt_kd_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47467),
            .ce(N__18972),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kd_7_LC_2_10_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kd_7_LC_2_10_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kd_7_LC_2_10_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Commands_frame_decoder.source_alt_kd_7_LC_2_10_5  (
            .in0(N__45012),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(alt_kd_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47467),
            .ce(N__18972),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kd_1_LC_2_10_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kd_1_LC_2_10_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kd_1_LC_2_10_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_alt_kd_1_LC_2_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45200),
            .lcout(alt_kd_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47467),
            .ce(N__18972),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kd_0_LC_2_10_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kd_0_LC_2_10_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kd_0_LC_2_10_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_alt_kd_0_LC_2_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27677),
            .lcout(alt_kd_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47467),
            .ce(N__18972),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_1_LC_2_11_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_1_LC_2_11_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_1_LC_2_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_1_LC_2_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18829),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47461),
            .ce(N__33610),
            .sr(N__43814));
    defparam \pid_alt.error_d_reg_esr_RNITF511_1_LC_2_12_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_RNITF511_1_LC_2_12_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_esr_RNITF511_1_LC_2_12_1 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_alt.error_d_reg_esr_RNITF511_1_LC_2_12_1  (
            .in0(N__18918),
            .in1(N__18859),
            .in2(_gnd_net_),
            .in3(N__18821),
            .lcout(\pid_alt.N_1074_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_p_reg_esr_RNIOI4P_0_0_LC_2_12_3 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_RNIOI4P_0_0_LC_2_12_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_p_reg_esr_RNIOI4P_0_0_LC_2_12_3 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \pid_alt.error_p_reg_esr_RNIOI4P_0_0_LC_2_12_3  (
            .in0(N__20723),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20777),
            .lcout(\pid_alt.g1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_esr_RNITF511_2_1_LC_2_12_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_RNITF511_2_1_LC_2_12_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_esr_RNITF511_2_1_LC_2_12_4 .LUT_INIT=16'b0101101010100101;
    LogicCell40 \pid_alt.error_d_reg_esr_RNITF511_2_1_LC_2_12_4  (
            .in0(N__18822),
            .in1(_gnd_net_),
            .in2(N__18873),
            .in3(N__18920),
            .lcout(\pid_alt.error_d_reg_esr_RNITF511_2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_fast_esr_RNIA7JS_1_LC_2_12_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_fast_esr_RNIA7JS_1_LC_2_12_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_fast_esr_RNIA7JS_1_LC_2_12_6 .LUT_INIT=16'b1101110101000100;
    LogicCell40 \pid_alt.error_d_reg_fast_esr_RNIA7JS_1_LC_2_12_6  (
            .in0(N__18860),
            .in1(N__18678),
            .in2(_gnd_net_),
            .in3(N__18919),
            .lcout(\pid_alt.N_1074_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI0J511_2_2_LC_2_12_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI0J511_2_2_LC_2_12_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI0J511_2_2_LC_2_12_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI0J511_2_2_LC_2_12_7  (
            .in0(N__19285),
            .in1(N__19317),
            .in2(_gnd_net_),
            .in3(N__19241),
            .lcout(\pid_alt.N_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI0J511_3_2_LC_2_13_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI0J511_3_2_LC_2_13_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI0J511_3_2_LC_2_13_1 .LUT_INIT=16'b0101101010100101;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI0J511_3_2_LC_2_13_1  (
            .in0(N__19248),
            .in1(_gnd_net_),
            .in2(N__19324),
            .in3(N__19284),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI0J511_3Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI0J511_1_2_LC_2_13_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI0J511_1_2_LC_2_13_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI0J511_1_2_LC_2_13_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI0J511_1_2_LC_2_13_2  (
            .in0(N__19283),
            .in1(N__19247),
            .in2(_gnd_net_),
            .in3(N__19313),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI0J511_1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_esr_RNIA37K_1_LC_2_13_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_RNIA37K_1_LC_2_13_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_esr_RNIA37K_1_LC_2_13_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \pid_alt.error_d_reg_esr_RNIA37K_1_LC_2_13_3  (
            .in0(N__18878),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18835),
            .lcout(),
            .ltout(\pid_alt.g0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_p_reg_esr_RNIL2AQ1_0_LC_2_13_4 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_RNIL2AQ1_0_LC_2_13_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_p_reg_esr_RNIL2AQ1_0_LC_2_13_4 .LUT_INIT=16'b1110000000001110;
    LogicCell40 \pid_alt.error_p_reg_esr_RNIL2AQ1_0_LC_2_13_4  (
            .in0(N__20724),
            .in1(N__20778),
            .in2(N__18522),
            .in3(N__18921),
            .lcout(\pid_alt.error_p_reg_esr_RNIL2AQ1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_19_LC_2_14_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_19_LC_2_14_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_19_LC_2_14_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_19_LC_2_14_0  (
            .in0(N__18651),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47440),
            .ce(N__33623),
            .sr(N__43832));
    defparam \pid_alt.error_d_reg_prev_esr_RNI86IM_0_19_LC_2_15_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI86IM_0_19_LC_2_15_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI86IM_0_19_LC_2_15_4 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI86IM_0_19_LC_2_15_4  (
            .in0(N__18614),
            .in1(N__18623),
            .in2(_gnd_net_),
            .in3(N__18649),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI86IM_0Z0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI86IM_19_LC_2_15_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI86IM_19_LC_2_15_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI86IM_19_LC_2_15_7 .LUT_INIT=16'b1010111100001010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI86IM_19_LC_2_15_7  (
            .in0(N__18650),
            .in1(_gnd_net_),
            .in2(N__18627),
            .in3(N__18615),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI86IMZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_p_reg_esr_2_LC_2_16_7 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_2_LC_2_16_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_2_LC_2_16_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_2_LC_2_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18600),
            .lcout(\pid_alt.error_p_regZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47418),
            .ce(N__46799),
            .sr(N__46619));
    defparam \pid_alt.error_p_reg_esr_1_LC_2_17_7 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_1_LC_2_17_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_1_LC_2_17_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_1_LC_2_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18588),
            .lcout(\pid_alt.error_p_regZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47408),
            .ce(N__46796),
            .sr(N__46618));
    defparam \pid_alt.error_p_reg_esr_10_LC_2_19_2 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_10_LC_2_19_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_10_LC_2_19_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_10_LC_2_19_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18573),
            .lcout(\pid_alt.error_p_regZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47380),
            .ce(N__46792),
            .sr(N__46615));
    defparam \Commands_frame_decoder.source_alt_kp_e_0_3_LC_2_20_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_3_LC_2_20_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_3_LC_2_20_3 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_kp_e_0_3_LC_2_20_3  (
            .in0(_gnd_net_),
            .in1(N__43365),
            .in2(_gnd_net_),
            .in3(N__46689),
            .lcout(alt_kp_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47368),
            .ce(N__22472),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kp_e_0_1_LC_2_21_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_1_LC_2_21_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_1_LC_2_21_7 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_kp_e_0_1_LC_2_21_7  (
            .in0(_gnd_net_),
            .in1(N__45225),
            .in2(_gnd_net_),
            .in3(N__46688),
            .lcout(alt_kp_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47355),
            .ce(N__22474),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kp_e_0_6_LC_2_22_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_6_LC_2_22_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_6_LC_2_22_5 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_kp_e_0_6_LC_2_22_5  (
            .in0(_gnd_net_),
            .in1(N__45015),
            .in2(_gnd_net_),
            .in3(N__46687),
            .lcout(alt_kp_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47341),
            .ce(N__22482),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kp_e_0_2_LC_2_22_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_2_LC_2_22_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_2_LC_2_22_7 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_kp_e_0_2_LC_2_22_7  (
            .in0(_gnd_net_),
            .in1(N__36880),
            .in2(_gnd_net_),
            .in3(N__46686),
            .lcout(alt_kp_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47341),
            .ce(N__22482),
            .sr(_gnd_net_));
    defparam \pid_alt.error_p_reg_esr_18_LC_2_23_4 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_18_LC_2_23_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_18_LC_2_23_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_18_LC_2_23_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18765),
            .lcout(\pid_alt.error_p_regZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47326),
            .ce(N__46786),
            .sr(N__46608));
    defparam \Commands_frame_decoder.source_alt_kd_6_LC_3_9_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kd_6_LC_3_9_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kd_6_LC_3_9_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_alt_kd_6_LC_3_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33439),
            .lcout(alt_kd_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47468),
            .ce(N__18964),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kd_5_LC_3_9_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kd_5_LC_3_9_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kd_5_LC_3_9_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_alt_kd_5_LC_3_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44240),
            .lcout(alt_kd_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47468),
            .ce(N__18964),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_esr_0_LC_3_10_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_0_LC_3_10_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_0_LC_3_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_0_LC_3_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18708),
            .lcout(\pid_alt.error_d_regZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47462),
            .ce(N__46804),
            .sr(N__46622));
    defparam \pid_alt.error_d_reg_fast_esr_RNICKGJ3_1_LC_3_12_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_fast_esr_RNICKGJ3_1_LC_3_12_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_fast_esr_RNICKGJ3_1_LC_3_12_0 .LUT_INIT=16'b0010101100100010;
    LogicCell40 \pid_alt.error_d_reg_fast_esr_RNICKGJ3_1_LC_3_12_0  (
            .in0(N__18699),
            .in1(N__18693),
            .in2(N__18660),
            .in3(N__18687),
            .lcout(),
            .ltout(\pid_alt.N_1080_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_p_reg_esr_RNIFTRL5_3_LC_3_12_1 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_RNIFTRL5_3_LC_3_12_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_p_reg_esr_RNIFTRL5_3_LC_3_12_1 .LUT_INIT=16'b1110100011010100;
    LogicCell40 \pid_alt.error_p_reg_esr_RNIFTRL5_3_LC_3_12_1  (
            .in0(N__19332),
            .in1(N__18933),
            .in2(N__18681),
            .in3(N__19198),
            .lcout(\pid_alt.error_p_reg_esr_RNIFTRL5Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_fast_esr_RNIA7JS_0_1_LC_3_12_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_fast_esr_RNIA7JS_0_1_LC_3_12_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_fast_esr_RNIA7JS_0_1_LC_3_12_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_d_reg_fast_esr_RNIA7JS_0_1_LC_3_12_7  (
            .in0(N__18677),
            .in1(N__18927),
            .in2(_gnd_net_),
            .in3(N__18872),
            .lcout(\pid_alt.N_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_esr_RNITF511_0_1_LC_3_13_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_RNITF511_0_1_LC_3_13_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_esr_RNITF511_0_1_LC_3_13_1 .LUT_INIT=16'b1010111100001010;
    LogicCell40 \pid_alt.error_d_reg_esr_RNITF511_0_1_LC_3_13_1  (
            .in0(N__18837),
            .in1(_gnd_net_),
            .in2(N__18879),
            .in3(N__18923),
            .lcout(),
            .ltout(\pid_alt.error_d_reg_esr_RNITF511_0Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIF0465_2_LC_3_13_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIF0465_2_LC_3_13_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIF0465_2_LC_3_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIF0465_2_LC_3_13_2  (
            .in0(N__30039),
            .in1(N__18948),
            .in2(N__18942),
            .in3(N__18939),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIF0465Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI0J511_2_LC_3_13_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI0J511_2_LC_3_13_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI0J511_2_LC_3_13_4 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI0J511_2_LC_3_13_4  (
            .in0(N__19292),
            .in1(N__19325),
            .in2(_gnd_net_),
            .in3(N__19256),
            .lcout(\pid_alt.N_1078_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_esr_RNITF511_1_1_LC_3_13_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_RNITF511_1_1_LC_3_13_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_esr_RNITF511_1_1_LC_3_13_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_d_reg_esr_RNITF511_1_1_LC_3_13_6  (
            .in0(N__18922),
            .in1(N__18874),
            .in2(_gnd_net_),
            .in3(N__18836),
            .lcout(),
            .ltout(\pid_alt.N_3_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNII5LS3_2_LC_3_13_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNII5LS3_2_LC_3_13_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNII5LS3_2_LC_3_13_7 .LUT_INIT=16'b0000100011001110;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNII5LS3_2_LC_3_13_7  (
            .in0(N__18786),
            .in1(N__18801),
            .in2(N__18795),
            .in3(N__18792),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNII5LS3Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_p_reg_esr_RNIOI4P_0_LC_3_14_2 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_RNIOI4P_0_LC_3_14_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_p_reg_esr_RNIOI4P_0_LC_3_14_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \pid_alt.error_p_reg_esr_RNIOI4P_0_LC_3_14_2  (
            .in0(_gnd_net_),
            .in1(N__20782),
            .in2(_gnd_net_),
            .in3(N__20722),
            .lcout(\pid_alt.g1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIK3024_19_LC_3_15_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIK3024_19_LC_3_15_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIK3024_19_LC_3_15_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIK3024_19_LC_3_15_0  (
            .in0(N__23195),
            .in1(N__23174),
            .in2(N__21227),
            .in3(N__30771),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIK3024Z0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_20_LC_3_15_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_20_LC_3_15_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_20_LC_3_15_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_20_LC_3_15_5  (
            .in0(N__19089),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47419),
            .ce(N__33624),
            .sr(N__43833));
    defparam \pid_alt.error_d_reg_prev_esr_RNIGGKM_20_LC_3_15_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIGGKM_20_LC_3_15_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIGGKM_20_LC_3_15_6 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIGGKM_20_LC_3_15_6  (
            .in0(N__24634),
            .in1(N__19101),
            .in2(_gnd_net_),
            .in3(N__19088),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIGGKMZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIMJHM_13_LC_3_16_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIMJHM_13_LC_3_16_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIMJHM_13_LC_3_16_1 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIMJHM_13_LC_3_16_1  (
            .in0(N__19371),
            .in1(N__19476),
            .in2(_gnd_net_),
            .in3(N__19500),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIMJHMZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIGGKM_0_20_LC_3_16_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIGGKM_0_20_LC_3_16_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIGGKM_0_20_LC_3_16_5 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIGGKM_0_20_LC_3_16_5  (
            .in0(N__19100),
            .in1(N__24608),
            .in2(_gnd_net_),
            .in3(N__19082),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIGGKM_0Z0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_p_reg_esr_3_LC_3_17_0 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_3_LC_3_17_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_3_LC_3_17_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_3_LC_3_17_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19062),
            .lcout(\pid_alt.error_p_regZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47394),
            .ce(N__46794),
            .sr(N__46617));
    defparam \Commands_frame_decoder.source_alt_kp_e_0_0_LC_3_21_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_0_LC_3_21_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_0_LC_3_21_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_kp_e_0_0_LC_3_21_0  (
            .in0(_gnd_net_),
            .in1(N__27681),
            .in2(_gnd_net_),
            .in3(N__46684),
            .lcout(alt_kp_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47342),
            .ce(N__22473),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kp_e_0_5_LC_3_21_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_5_LC_3_21_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_5_LC_3_21_5 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Commands_frame_decoder.source_alt_kp_e_0_5_LC_3_21_5  (
            .in0(N__46685),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33435),
            .lcout(alt_kp_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47342),
            .ce(N__22473),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kp_0_e_0_4_LC_3_22_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kp_0_e_0_4_LC_3_22_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kp_0_e_0_4_LC_3_22_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_kp_0_e_0_4_LC_3_22_6  (
            .in0(_gnd_net_),
            .in1(N__44291),
            .in2(_gnd_net_),
            .in3(N__46683),
            .lcout(alt_kp_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47327),
            .ce(N__22481),
            .sr(_gnd_net_));
    defparam \pid_alt.error_p_reg_esr_12_LC_3_23_1 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_12_LC_3_23_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_12_LC_3_23_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_12_LC_3_23_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19008),
            .lcout(\pid_alt.error_p_regZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47313),
            .ce(N__46783),
            .sr(N__46605));
    defparam \Commands_frame_decoder.state_RNIRSI31_11_LC_4_9_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIRSI31_11_LC_4_9_3 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIRSI31_11_LC_4_9_3 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \Commands_frame_decoder.state_RNIRSI31_11_LC_4_9_3  (
            .in0(N__23709),
            .in1(N__27040),
            .in2(_gnd_net_),
            .in3(N__44092),
            .lcout(\Commands_frame_decoder.source_alt_kd_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kd_4_LC_4_10_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kd_4_LC_4_10_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kd_4_LC_4_10_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_alt_kd_4_LC_4_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45350),
            .lcout(alt_kd_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47455),
            .ce(N__18965),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_3_LC_4_11_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_3_LC_4_11_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_3_LC_4_11_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_3_LC_4_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19158),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47447),
            .ce(N__33602),
            .sr(N__43808));
    defparam \pid_alt.error_d_reg_prev_esr_RNIE77K_3_LC_4_12_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIE77K_3_LC_4_12_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIE77K_3_LC_4_12_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIE77K_3_LC_4_12_6  (
            .in0(N__19174),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19157),
            .lcout(\pid_alt.g0_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI3M511_0_3_LC_4_13_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI3M511_0_3_LC_4_13_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI3M511_0_3_LC_4_13_0 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI3M511_0_3_LC_4_13_0  (
            .in0(N__19199),
            .in1(N__19175),
            .in2(_gnd_net_),
            .in3(N__19156),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI3M511_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI0J511_0_2_LC_4_13_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI0J511_0_2_LC_4_13_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI0J511_0_2_LC_4_13_1 .LUT_INIT=16'b1101110101000100;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI0J511_0_2_LC_4_13_1  (
            .in0(N__19326),
            .in1(N__19293),
            .in2(_gnd_net_),
            .in3(N__19257),
            .lcout(),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNI0J511_0Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNILDG87_2_LC_4_13_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNILDG87_2_LC_4_13_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNILDG87_2_LC_4_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNILDG87_2_LC_4_13_2  (
            .in0(N__29997),
            .in1(N__19215),
            .in2(N__19209),
            .in3(N__19206),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNILDG87Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI3M511_3_LC_4_13_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI3M511_3_LC_4_13_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI3M511_3_LC_4_13_4 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI3M511_3_LC_4_13_4  (
            .in0(N__19200),
            .in1(N__19176),
            .in2(_gnd_net_),
            .in3(N__19155),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI3M511Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_p_reg_esr_RNI3SMI1_0_LC_4_14_7 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_RNI3SMI1_0_LC_4_14_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_p_reg_esr_RNI3SMI1_0_LC_4_14_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \pid_alt.error_p_reg_esr_RNI3SMI1_0_LC_4_14_7  (
            .in0(N__30138),
            .in1(N__20783),
            .in2(_gnd_net_),
            .in3(N__20734),
            .lcout(\pid_alt.error_p_reg_esr_RNI3SMI1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI8IQ14_18_LC_4_15_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI8IQ14_18_LC_4_15_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI8IQ14_18_LC_4_15_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI8IQ14_18_LC_4_15_0  (
            .in0(N__19115),
            .in1(N__19122),
            .in2(N__20888),
            .in3(N__30809),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI8IQ14Z0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI53IM_18_LC_4_15_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI53IM_18_LC_4_15_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI53IM_18_LC_4_15_1 .LUT_INIT=16'b1010111100001010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI53IM_18_LC_4_15_1  (
            .in0(N__19430),
            .in1(_gnd_net_),
            .in2(N__19407),
            .in3(N__19452),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI53IMZ0Z_18 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNI53IMZ0Z_18_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIOTT02_18_LC_4_15_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIOTT02_18_LC_4_15_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIOTT02_18_LC_4_15_2 .LUT_INIT=16'b1111101010100000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIOTT02_18_LC_4_15_2  (
            .in0(N__19116),
            .in1(_gnd_net_),
            .in2(N__19104),
            .in3(N__30810),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIOTT02Z0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI53IM_0_18_LC_4_15_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI53IM_0_18_LC_4_15_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI53IM_0_18_LC_4_15_4 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI53IM_0_18_LC_4_15_4  (
            .in0(N__19451),
            .in1(N__19403),
            .in2(_gnd_net_),
            .in3(N__19429),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI53IM_0Z0Z_18 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNI53IM_0Z0Z_18_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIGKS02_17_LC_4_15_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIGKS02_17_LC_4_15_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIGKS02_17_LC_4_15_5 .LUT_INIT=16'b1111110011000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIGKS02_17_LC_4_15_5  (
            .in0(_gnd_net_),
            .in1(N__19389),
            .in2(N__19434),
            .in3(N__30846),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIGKS02Z0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_18_LC_4_15_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_18_LC_4_15_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_18_LC_4_15_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_18_LC_4_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19431),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47409),
            .ce(N__33620),
            .sr(N__43824));
    defparam \pid_alt.error_d_reg_prev_esr_RNIOVN14_17_LC_4_15_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIOVN14_17_LC_4_15_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIOVN14_17_LC_4_15_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIOVN14_17_LC_4_15_7  (
            .in0(N__19395),
            .in1(N__19388),
            .in2(N__20930),
            .in3(N__30845),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIOVN14Z0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_12_LC_4_16_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_12_LC_4_16_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_12_LC_4_16_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_12_LC_4_16_0  (
            .in0(N__19524),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47395),
            .ce(N__33625),
            .sr(N__43834));
    defparam \pid_alt.error_d_reg_prev_esr_RNIMJHM_0_13_LC_4_16_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIMJHM_0_13_LC_4_16_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIMJHM_0_13_LC_4_16_1 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIMJHM_0_13_LC_4_16_1  (
            .in0(N__19370),
            .in1(N__19475),
            .in2(_gnd_net_),
            .in3(N__19498),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIMJHM_0Z0Z_13 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNIMJHM_0Z0Z_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNISAO32_12_LC_4_16_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNISAO32_12_LC_4_16_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNISAO32_12_LC_4_16_2 .LUT_INIT=16'b1111110011000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNISAO32_12_LC_4_16_2  (
            .in0(_gnd_net_),
            .in1(N__19347),
            .in2(N__19350),
            .in3(N__30215),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNISAO32Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIJGHM_12_LC_4_16_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIJGHM_12_LC_4_16_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIJGHM_12_LC_4_16_3 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIJGHM_12_LC_4_16_3  (
            .in0(N__19548),
            .in1(N__19533),
            .in2(_gnd_net_),
            .in3(N__19523),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIJGHMZ0Z_12 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNIJGHMZ0Z_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIT4AF4_12_LC_4_16_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIT4AF4_12_LC_4_16_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIT4AF4_12_LC_4_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIT4AF4_12_LC_4_16_4  (
            .in0(N__21119),
            .in1(N__19341),
            .in2(N__19335),
            .in3(N__30214),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIT4AF4Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIJGHM_0_12_LC_4_16_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIJGHM_0_12_LC_4_16_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIJGHM_0_12_LC_4_16_5 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIJGHM_0_12_LC_4_16_5  (
            .in0(N__19547),
            .in1(N__19532),
            .in2(_gnd_net_),
            .in3(N__19522),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIJGHM_0Z0Z_12 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNIJGHM_0Z0Z_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI1QHB2_11_LC_4_16_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI1QHB2_11_LC_4_16_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI1QHB2_11_LC_4_16_6 .LUT_INIT=16'b1111101010100000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI1QHB2_11_LC_4_16_6  (
            .in0(N__19617),
            .in1(_gnd_net_),
            .in2(N__19503),
            .in3(N__30255),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI1QHB2Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_13_LC_4_16_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_13_LC_4_16_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_13_LC_4_16_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_13_LC_4_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19499),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47395),
            .ce(N__33625),
            .sr(N__43834));
    defparam \pid_alt.error_d_reg_prev_esr_0_LC_4_17_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_0_LC_4_17_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_0_LC_4_17_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_0_LC_4_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20739),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47381),
            .ce(N__33628),
            .sr(N__43840));
    defparam \pid_alt.error_d_reg_prev_esr_RNIKKKM_0_22_LC_4_18_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIKKKM_0_22_LC_4_18_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIKKKM_0_22_LC_4_18_7 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIKKKM_0_22_LC_4_18_7  (
            .in0(N__20015),
            .in1(N__19997),
            .in2(_gnd_net_),
            .in3(N__24622),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIKKKM_0Z0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIMMKM_23_LC_4_19_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIMMKM_23_LC_4_19_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIMMKM_23_LC_4_19_1 .LUT_INIT=16'b1101110101000100;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIMMKM_23_LC_4_19_1  (
            .in0(N__20187),
            .in1(N__24614),
            .in2(_gnd_net_),
            .in3(N__20211),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIMMKMZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_CH4data_esr_5_LC_4_20_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH4data_esr_5_LC_4_20_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH4data_esr_5_LC_4_20_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH4data_esr_5_LC_4_20_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44292),
            .lcout(frame_decoder_CH4data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47343),
            .ce(N__26400),
            .sr(N__43863));
    defparam \pid_alt.error_p_reg_esr_11_LC_4_21_6 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_11_LC_4_21_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_11_LC_4_21_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_11_LC_4_21_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19464),
            .lcout(\pid_alt.error_p_regZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47328),
            .ce(N__46787),
            .sr(N__46609));
    defparam \dron_frame_decoder_1.WDT_RNIA9RK1_11_LC_5_8_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.WDT_RNIA9RK1_11_LC_5_8_1 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.WDT_RNIA9RK1_11_LC_5_8_1 .LUT_INIT=16'b0000001100010011;
    LogicCell40 \dron_frame_decoder_1.WDT_RNIA9RK1_11_LC_5_8_1  (
            .in0(N__20243),
            .in1(N__20495),
            .in2(N__20531),
            .in3(N__20264),
            .lcout(\dron_frame_decoder_1.WDT10_0_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.WDT_RNIM3K1_4_LC_5_8_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.WDT_RNIM3K1_4_LC_5_8_2 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.WDT_RNIM3K1_4_LC_5_8_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \dron_frame_decoder_1.WDT_RNIM3K1_4_LC_5_8_2  (
            .in0(N__20322),
            .in1(N__20385),
            .in2(N__20304),
            .in3(N__20406),
            .lcout(),
            .ltout(\dron_frame_decoder_1.WDT10lto9_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.WDT_RNI9TKF_6_LC_5_8_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.WDT_RNI9TKF_6_LC_5_8_3 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.WDT_RNI9TKF_6_LC_5_8_3 .LUT_INIT=16'b1010101010001010;
    LogicCell40 \dron_frame_decoder_1.WDT_RNI9TKF_6_LC_5_8_3  (
            .in0(N__20283),
            .in1(N__20343),
            .in2(N__19578),
            .in3(N__20364),
            .lcout(\dron_frame_decoder_1.WDT10lt12_0 ),
            .ltout(\dron_frame_decoder_1.WDT10lt12_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.WDT_RNIBUTU2_15_LC_5_8_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.WDT_RNIBUTU2_15_LC_5_8_4 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.WDT_RNIBUTU2_15_LC_5_8_4 .LUT_INIT=16'b0111111101010101;
    LogicCell40 \dron_frame_decoder_1.WDT_RNIBUTU2_15_LC_5_8_4  (
            .in0(N__20465),
            .in1(N__20527),
            .in2(N__19575),
            .in3(N__19572),
            .lcout(\dron_frame_decoder_1.WDT10_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.WDT_RNINA9N1_11_LC_5_8_6 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.WDT_RNINA9N1_11_LC_5_8_6 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.WDT_RNINA9N1_11_LC_5_8_6 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \dron_frame_decoder_1.WDT_RNINA9N1_11_LC_5_8_6  (
            .in0(N__20265),
            .in1(N__20244),
            .in2(N__20535),
            .in3(N__19566),
            .lcout(\dron_frame_decoder_1.WDT10lt14_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.WDT_RNIPI9R2_15_LC_5_9_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.WDT_RNIPI9R2_15_LC_5_9_3 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.WDT_RNIPI9R2_15_LC_5_9_3 .LUT_INIT=16'b0000010100010101;
    LogicCell40 \dron_frame_decoder_1.WDT_RNIPI9R2_15_LC_5_9_3  (
            .in0(N__29672),
            .in1(N__20499),
            .in2(N__20469),
            .in3(N__19560),
            .lcout(\dron_frame_decoder_1.WDT_RNIPI9R2Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.source_data_valid_esr_RNO_LC_5_11_3 .C_ON=1'b0;
    defparam \pid_alt.source_data_valid_esr_RNO_LC_5_11_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.source_data_valid_esr_RNO_LC_5_11_3 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \pid_alt.source_data_valid_esr_RNO_LC_5_11_3  (
            .in0(_gnd_net_),
            .in1(N__24961),
            .in2(_gnd_net_),
            .in3(N__44100),
            .lcout(\pid_alt.state_1_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.source_data_valid_esr_LC_5_12_0 .C_ON=1'b0;
    defparam \pid_alt.source_data_valid_esr_LC_5_12_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_data_valid_esr_LC_5_12_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.source_data_valid_esr_LC_5_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33229),
            .lcout(pid_altitude_dv),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47430),
            .ce(N__19554),
            .sr(N__43809));
    defparam \pid_alt.source_pid_1_4_LC_5_13_6 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_4_LC_5_13_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_4_LC_5_13_6 .LUT_INIT=16'b1111101011011000;
    LogicCell40 \pid_alt.source_pid_1_4_LC_5_13_6  (
            .in0(N__33204),
            .in1(N__25914),
            .in2(N__29396),
            .in3(N__24165),
            .lcout(throttle_command_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47420),
            .ce(),
            .sr(N__27875));
    defparam \pid_alt.error_d_reg_prev_esr_RNIKQBI4_10_LC_5_14_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIKQBI4_10_LC_5_14_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIKQBI4_10_LC_5_14_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIKQBI4_10_LC_5_14_0  (
            .in0(N__19637),
            .in1(N__19644),
            .in2(N__23082),
            .in3(N__30299),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIKQBI4Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIDAHM_10_LC_5_14_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIDAHM_10_LC_5_14_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIDAHM_10_LC_5_14_1 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIDAHM_10_LC_5_14_1  (
            .in0(N__22974),
            .in1(N__22946),
            .in2(_gnd_net_),
            .in3(N__22930),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIDAHMZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI7E8R_11_LC_5_14_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI7E8R_11_LC_5_14_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI7E8R_11_LC_5_14_2 .LUT_INIT=16'b1010111100001010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI7E8R_11_LC_5_14_2  (
            .in0(N__19673),
            .in1(_gnd_net_),
            .in2(N__19686),
            .in3(N__19704),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI7E8RZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_11_LC_5_14_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_11_LC_5_14_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_11_LC_5_14_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_11_LC_5_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19674),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47410),
            .ce(N__33611),
            .sr(N__43815));
    defparam \pid_alt.error_d_reg_prev_esr_10_LC_5_14_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_10_LC_5_14_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_10_LC_5_14_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_10_LC_5_14_4  (
            .in0(N__22931),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47410),
            .ce(N__33611),
            .sr(N__43815));
    defparam \pid_alt.error_d_reg_prev_esr_RNI7E8R_0_11_LC_5_14_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI7E8R_0_11_LC_5_14_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI7E8R_0_11_LC_5_14_5 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI7E8R_0_11_LC_5_14_5  (
            .in0(N__19703),
            .in1(N__19682),
            .in2(_gnd_net_),
            .in3(N__19672),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI7E8R_0Z0Z_11 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNI7E8R_0Z0Z_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIOFGB2_10_LC_5_14_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIOFGB2_10_LC_5_14_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIOFGB2_10_LC_5_14_6 .LUT_INIT=16'b1111101010100000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIOFGB2_10_LC_5_14_6  (
            .in0(N__19638),
            .in1(_gnd_net_),
            .in2(N__19629),
            .in3(N__30300),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIOFGB2Z0Z_10 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNIOFGB2Z0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIP92N4_11_LC_5_14_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIP92N4_11_LC_5_14_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIP92N4_11_LC_5_14_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIP92N4_11_LC_5_14_7  (
            .in0(N__19626),
            .in1(N__19613),
            .in2(N__19602),
            .in3(N__30250),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIP92N4Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI8BR02_16_LC_5_15_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI8BR02_16_LC_5_15_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI8BR02_16_LC_5_15_0 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI8BR02_16_LC_5_15_0  (
            .in0(N__19599),
            .in1(N__19593),
            .in2(_gnd_net_),
            .in3(N__30882),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI8BR02Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIVSHM_16_LC_5_15_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIVSHM_16_LC_5_15_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIVSHM_16_LC_5_15_1 .LUT_INIT=16'b1010111100001010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIVSHM_16_LC_5_15_1  (
            .in0(N__19754),
            .in1(_gnd_net_),
            .in2(N__19767),
            .in3(N__19785),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIVSHMZ0Z_16 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNIVSHMZ0Z_16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI8DL14_16_LC_5_15_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI8DL14_16_LC_5_15_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI8DL14_16_LC_5_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI8DL14_16_LC_5_15_2  (
            .in0(N__20966),
            .in1(N__19592),
            .in2(N__19788),
            .in3(N__30881),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI8DL14Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_16_LC_5_15_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_16_LC_5_15_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_16_LC_5_15_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_16_LC_5_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19755),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47396),
            .ce(N__33615),
            .sr(N__43819));
    defparam \pid_alt.error_d_reg_prev_esr_RNI02Q02_15_LC_5_15_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI02Q02_15_LC_5_15_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI02Q02_15_LC_5_15_5 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI02Q02_15_LC_5_15_5  (
            .in0(N__19731),
            .in1(N__19869),
            .in2(_gnd_net_),
            .in3(N__30915),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI02Q02Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIVSHM_0_16_LC_5_15_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIVSHM_0_16_LC_5_15_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIVSHM_0_16_LC_5_15_6 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIVSHM_0_16_LC_5_15_6  (
            .in0(N__19784),
            .in1(N__19763),
            .in2(_gnd_net_),
            .in3(N__19753),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIVSHM_0Z0Z_16 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNIVSHM_0Z0Z_16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIOQI14_15_LC_5_15_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIOQI14_15_LC_5_15_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIOQI14_15_LC_5_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIOQI14_15_LC_5_15_7  (
            .in0(N__21011),
            .in1(N__19868),
            .in2(N__19725),
            .in3(N__30914),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIOQI14Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_7_LC_5_16_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_7_LC_5_16_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_7_LC_5_16_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_7_LC_5_16_0  (
            .in0(N__19950),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47382),
            .ce(N__33621),
            .sr(N__43825));
    defparam \pid_alt.error_d_reg_prev_esr_RNII5611_0_8_LC_5_16_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNII5611_0_8_LC_5_16_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNII5611_0_8_LC_5_16_1 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNII5611_0_8_LC_5_16_1  (
            .in0(N__19928),
            .in1(N__19880),
            .in2(_gnd_net_),
            .in3(N__19903),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNII5611_0Z0Z_8 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNII5611_0Z0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI7T3T2_7_LC_5_16_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI7T3T2_7_LC_5_16_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI7T3T2_7_LC_5_16_2 .LUT_INIT=16'b1111110011000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI7T3T2_7_LC_5_16_2  (
            .in0(_gnd_net_),
            .in1(N__19719),
            .in2(N__19722),
            .in3(N__30432),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI7T3T2Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIF2611_7_LC_5_16_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIF2611_7_LC_5_16_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIF2611_7_LC_5_16_3 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIF2611_7_LC_5_16_3  (
            .in0(N__19974),
            .in1(N__19959),
            .in2(_gnd_net_),
            .in3(N__19949),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIF2611Z0Z_7 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNIF2611Z0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI5G6Q5_7_LC_5_16_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI5G6Q5_7_LC_5_16_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI5G6Q5_7_LC_5_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI5G6Q5_7_LC_5_16_4  (
            .in0(N__26316),
            .in1(N__19713),
            .in2(N__19707),
            .in3(N__30431),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI5G6Q5Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIF2611_0_7_LC_5_16_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIF2611_0_7_LC_5_16_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIF2611_0_7_LC_5_16_5 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIF2611_0_7_LC_5_16_5  (
            .in0(N__19973),
            .in1(N__19958),
            .in2(_gnd_net_),
            .in3(N__19948),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIF2611_0Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNII5611_8_LC_5_17_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNII5611_8_LC_5_17_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNII5611_8_LC_5_17_0 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNII5611_8_LC_5_17_0  (
            .in0(N__19929),
            .in1(N__19881),
            .in2(_gnd_net_),
            .in3(N__19904),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNII5611Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_8_LC_5_17_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_8_LC_5_17_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_8_LC_5_17_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_8_LC_5_17_1  (
            .in0(N__19905),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47369),
            .ce(N__33626),
            .sr(N__43835));
    defparam \pid_alt.error_d_reg_prev_esr_RNISPHM_15_LC_5_17_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNISPHM_15_LC_5_17_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNISPHM_15_LC_5_17_3 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNISPHM_15_LC_5_17_3  (
            .in0(N__19839),
            .in1(N__19851),
            .in2(_gnd_net_),
            .in3(N__19817),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNISPHMZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_15_LC_5_17_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_15_LC_5_17_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_15_LC_5_17_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_15_LC_5_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19818),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47369),
            .ce(N__33626),
            .sr(N__43835));
    defparam \pid_alt.error_d_reg_prev_esr_RNI2Q08_0_LC_5_17_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI2Q08_0_LC_5_17_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI2Q08_0_LC_5_17_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI2Q08_0_LC_5_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19857),
            .lcout(\pid_alt.error_d_reg_prev_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI88G14_14_LC_5_18_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI88G14_14_LC_5_18_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI88G14_14_LC_5_18_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI88G14_14_LC_5_18_0  (
            .in0(N__19794),
            .in1(N__20102),
            .in2(N__21047),
            .in3(N__30950),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI88G14Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNISPHM_0_15_LC_5_18_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNISPHM_0_15_LC_5_18_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNISPHM_0_15_LC_5_18_1 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNISPHM_0_15_LC_5_18_1  (
            .in0(N__19850),
            .in1(N__19838),
            .in2(_gnd_net_),
            .in3(N__19816),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNISPHM_0Z0Z_15 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNISPHM_0Z0Z_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIOOO02_14_LC_5_18_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIOOO02_14_LC_5_18_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIOOO02_14_LC_5_18_2 .LUT_INIT=16'b1111110011000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIOOO02_14_LC_5_18_2  (
            .in0(_gnd_net_),
            .in1(N__20103),
            .in2(N__20106),
            .in3(N__30951),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIOOO02Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIPMHM_14_LC_5_18_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIPMHM_14_LC_5_18_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIPMHM_14_LC_5_18_3 .LUT_INIT=16'b1010111100001010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIPMHM_14_LC_5_18_3  (
            .in0(N__20072),
            .in1(_gnd_net_),
            .in2(N__20052),
            .in3(N__20094),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIPMHMZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIPMHM_0_14_LC_5_18_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIPMHM_0_14_LC_5_18_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIPMHM_0_14_LC_5_18_4 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIPMHM_0_14_LC_5_18_4  (
            .in0(N__20093),
            .in1(N__20048),
            .in2(_gnd_net_),
            .in3(N__20071),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIPMHM_0Z0Z_14 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNIPMHM_0Z0Z_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNICQF44_13_LC_5_18_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNICQF44_13_LC_5_18_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNICQF44_13_LC_5_18_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNICQF44_13_LC_5_18_5  (
            .in0(N__20039),
            .in1(N__21086),
            .in2(N__20076),
            .in3(N__30185),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNICQF44Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_14_LC_5_18_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_14_LC_5_18_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_14_LC_5_18_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_14_LC_5_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20073),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47356),
            .ce(N__33629),
            .sr(N__43841));
    defparam \pid_alt.error_d_reg_prev_esr_RNIGFN02_13_LC_5_18_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIGFN02_13_LC_5_18_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIGFN02_13_LC_5_18_7 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIGFN02_13_LC_5_18_7  (
            .in0(N__20040),
            .in1(N__20025),
            .in2(_gnd_net_),
            .in3(N__30186),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIGFN02Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_22_LC_5_19_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_22_LC_5_19_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_22_LC_5_19_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_22_LC_5_19_0  (
            .in0(N__20004),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47344),
            .ce(N__33630),
            .sr(N__43849));
    defparam \pid_alt.error_d_reg_prev_esr_RNIMMKM_0_23_LC_5_19_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIMMKM_0_23_LC_5_19_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIMMKM_0_23_LC_5_19_1 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIMMKM_0_23_LC_5_19_1  (
            .in0(N__20186),
            .in1(N__20206),
            .in2(_gnd_net_),
            .in3(N__24612),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIMMKM_0Z0Z_23 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNIMMKM_0Z0Z_23_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI6BU12_22_LC_5_19_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI6BU12_22_LC_5_19_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI6BU12_22_LC_5_19_2 .LUT_INIT=16'b1111110011000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI6BU12_22_LC_5_19_2  (
            .in0(_gnd_net_),
            .in1(N__20226),
            .in2(N__20019),
            .in3(N__30703),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI6BU12Z0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIKKKM_22_LC_5_19_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIKKKM_22_LC_5_19_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIKKKM_22_LC_5_19_3 .LUT_INIT=16'b1101110101000100;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIKKKM_22_LC_5_19_3  (
            .in0(N__20016),
            .in1(N__20003),
            .in2(_gnd_net_),
            .in3(N__24613),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIKKKMZ0Z_22 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNIKKKMZ0Z_22_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI8IS34_22_LC_5_19_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI8IS34_22_LC_5_19_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI8IS34_22_LC_5_19_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI8IS34_22_LC_5_19_4  (
            .in0(N__20220),
            .in1(N__23052),
            .in2(N__20214),
            .in3(N__30704),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI8IS34Z0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_23_LC_5_19_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_23_LC_5_19_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_23_LC_5_19_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_23_LC_5_19_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20207),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47344),
            .ce(N__33630),
            .sr(N__43849));
    defparam \pid_alt.error_p_reg_esr_4_LC_5_23_4 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_4_LC_5_23_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_4_LC_5_23_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_4_LC_5_23_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20175),
            .lcout(\pid_alt.error_p_regZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47293),
            .ce(N__46782),
            .sr(N__46602));
    defparam \uart_drone_sync.Q_0__0_LC_7_6_3 .C_ON=1'b0;
    defparam \uart_drone_sync.Q_0__0_LC_7_6_3 .SEQ_MODE=4'b1000;
    defparam \uart_drone_sync.Q_0__0_LC_7_6_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone_sync.Q_0__0_LC_7_6_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22329),
            .lcout(debug_CH0_16A_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47463),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.WDT_0_LC_7_7_0 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_0_LC_7_7_0 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_0_LC_7_7_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_0_LC_7_7_0  (
            .in0(_gnd_net_),
            .in1(N__20139),
            .in2(N__20160),
            .in3(N__20159),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_0 ),
            .ltout(),
            .carryin(bfn_7_7_0_),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_0 ),
            .clk(N__47456),
            .ce(),
            .sr(N__22323));
    defparam \dron_frame_decoder_1.WDT_1_LC_7_7_1 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_1_LC_7_7_1 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_1_LC_7_7_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_1_LC_7_7_1  (
            .in0(_gnd_net_),
            .in1(N__20133),
            .in2(_gnd_net_),
            .in3(N__20127),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_1 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_0 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_1 ),
            .clk(N__47456),
            .ce(),
            .sr(N__22323));
    defparam \dron_frame_decoder_1.WDT_2_LC_7_7_2 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_2_LC_7_7_2 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_2_LC_7_7_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_2_LC_7_7_2  (
            .in0(_gnd_net_),
            .in1(N__20124),
            .in2(_gnd_net_),
            .in3(N__20118),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_2 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_1 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_2 ),
            .clk(N__47456),
            .ce(),
            .sr(N__22323));
    defparam \dron_frame_decoder_1.WDT_3_LC_7_7_3 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_3_LC_7_7_3 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_3_LC_7_7_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_3_LC_7_7_3  (
            .in0(_gnd_net_),
            .in1(N__20115),
            .in2(_gnd_net_),
            .in3(N__20109),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_3 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_2 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_3 ),
            .clk(N__47456),
            .ce(),
            .sr(N__22323));
    defparam \dron_frame_decoder_1.WDT_4_LC_7_7_4 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_4_LC_7_7_4 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_4_LC_7_7_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_4_LC_7_7_4  (
            .in0(_gnd_net_),
            .in1(N__20402),
            .in2(_gnd_net_),
            .in3(N__20388),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_4 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_3 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_4 ),
            .clk(N__47456),
            .ce(),
            .sr(N__22323));
    defparam \dron_frame_decoder_1.WDT_5_LC_7_7_5 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_5_LC_7_7_5 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_5_LC_7_7_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_5_LC_7_7_5  (
            .in0(_gnd_net_),
            .in1(N__20381),
            .in2(_gnd_net_),
            .in3(N__20367),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_5 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_4 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_5 ),
            .clk(N__47456),
            .ce(),
            .sr(N__22323));
    defparam \dron_frame_decoder_1.WDT_6_LC_7_7_6 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_6_LC_7_7_6 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_6_LC_7_7_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_6_LC_7_7_6  (
            .in0(_gnd_net_),
            .in1(N__20360),
            .in2(_gnd_net_),
            .in3(N__20346),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_6 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_5 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_6 ),
            .clk(N__47456),
            .ce(),
            .sr(N__22323));
    defparam \dron_frame_decoder_1.WDT_7_LC_7_7_7 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_7_LC_7_7_7 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_7_LC_7_7_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_7_LC_7_7_7  (
            .in0(_gnd_net_),
            .in1(N__20339),
            .in2(_gnd_net_),
            .in3(N__20325),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_7 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_6 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_7 ),
            .clk(N__47456),
            .ce(),
            .sr(N__22323));
    defparam \dron_frame_decoder_1.WDT_8_LC_7_8_0 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_8_LC_7_8_0 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_8_LC_7_8_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_8_LC_7_8_0  (
            .in0(_gnd_net_),
            .in1(N__20321),
            .in2(_gnd_net_),
            .in3(N__20307),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_8 ),
            .ltout(),
            .carryin(bfn_7_8_0_),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_8 ),
            .clk(N__47448),
            .ce(),
            .sr(N__22322));
    defparam \dron_frame_decoder_1.WDT_9_LC_7_8_1 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_9_LC_7_8_1 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_9_LC_7_8_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_9_LC_7_8_1  (
            .in0(_gnd_net_),
            .in1(N__20300),
            .in2(_gnd_net_),
            .in3(N__20286),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_9 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_8 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_9 ),
            .clk(N__47448),
            .ce(),
            .sr(N__22322));
    defparam \dron_frame_decoder_1.WDT_10_LC_7_8_2 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_10_LC_7_8_2 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_10_LC_7_8_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_10_LC_7_8_2  (
            .in0(_gnd_net_),
            .in1(N__20282),
            .in2(_gnd_net_),
            .in3(N__20268),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_10 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_9 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_10 ),
            .clk(N__47448),
            .ce(),
            .sr(N__22322));
    defparam \dron_frame_decoder_1.WDT_11_LC_7_8_3 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_11_LC_7_8_3 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_11_LC_7_8_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_11_LC_7_8_3  (
            .in0(_gnd_net_),
            .in1(N__20263),
            .in2(_gnd_net_),
            .in3(N__20247),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_11 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_10 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_11 ),
            .clk(N__47448),
            .ce(),
            .sr(N__22322));
    defparam \dron_frame_decoder_1.WDT_12_LC_7_8_4 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_12_LC_7_8_4 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_12_LC_7_8_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_12_LC_7_8_4  (
            .in0(_gnd_net_),
            .in1(N__20242),
            .in2(_gnd_net_),
            .in3(N__20538),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_12 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_11 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_12 ),
            .clk(N__47448),
            .ce(),
            .sr(N__22322));
    defparam \dron_frame_decoder_1.WDT_13_LC_7_8_5 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_13_LC_7_8_5 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_13_LC_7_8_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_13_LC_7_8_5  (
            .in0(_gnd_net_),
            .in1(N__20523),
            .in2(_gnd_net_),
            .in3(N__20502),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_13 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_12 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_13 ),
            .clk(N__47448),
            .ce(),
            .sr(N__22322));
    defparam \dron_frame_decoder_1.WDT_14_LC_7_8_6 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_14_LC_7_8_6 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_14_LC_7_8_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_14_LC_7_8_6  (
            .in0(_gnd_net_),
            .in1(N__20494),
            .in2(_gnd_net_),
            .in3(N__20475),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_14 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_13 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_14 ),
            .clk(N__47448),
            .ce(),
            .sr(N__22322));
    defparam \dron_frame_decoder_1.WDT_15_LC_7_8_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.WDT_15_LC_7_8_7 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_15_LC_7_8_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \dron_frame_decoder_1.WDT_15_LC_7_8_7  (
            .in0(_gnd_net_),
            .in1(N__20458),
            .in2(_gnd_net_),
            .in3(N__20472),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47448),
            .ce(),
            .sr(N__22322));
    defparam \dron_frame_decoder_1.state_3_LC_7_9_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_3_LC_7_9_3 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.state_3_LC_7_9_3 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \dron_frame_decoder_1.state_3_LC_7_9_3  (
            .in0(N__22515),
            .in1(N__20412),
            .in2(N__20559),
            .in3(N__20438),
            .lcout(\dron_frame_decoder_1.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47441),
            .ce(),
            .sr(N__43800));
    defparam \dron_frame_decoder_1.state_5_LC_7_9_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_5_LC_7_9_5 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.state_5_LC_7_9_5 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \dron_frame_decoder_1.state_5_LC_7_9_5  (
            .in0(N__22516),
            .in1(N__22392),
            .in2(N__20427),
            .in3(N__29662),
            .lcout(\dron_frame_decoder_1.stateZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47441),
            .ce(),
            .sr(N__43800));
    defparam \dron_frame_decoder_1.state_2_LC_7_9_6 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_2_LC_7_9_6 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.state_2_LC_7_9_6 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \dron_frame_decoder_1.state_2_LC_7_9_6  (
            .in0(N__29661),
            .in1(N__20423),
            .in2(N__20439),
            .in3(N__22514),
            .lcout(\dron_frame_decoder_1.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47441),
            .ce(),
            .sr(N__43800));
    defparam \dron_frame_decoder_1.state_ns_0_i_a2_0_4_3_LC_7_10_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_ns_0_i_a2_0_4_3_LC_7_10_3 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_ns_0_i_a2_0_4_3_LC_7_10_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \dron_frame_decoder_1.state_ns_0_i_a2_0_4_3_LC_7_10_3  (
            .in0(N__26190),
            .in1(N__25209),
            .in2(N__25137),
            .in3(N__25002),
            .lcout(\dron_frame_decoder_1.N_188_4 ),
            .ltout(\dron_frame_decoder_1.N_188_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_RNO_0_3_LC_7_10_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNO_0_3_LC_7_10_4 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNO_0_3_LC_7_10_4 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \dron_frame_decoder_1.state_RNO_0_3_LC_7_10_4  (
            .in0(N__20677),
            .in1(_gnd_net_),
            .in2(N__20415),
            .in3(_gnd_net_),
            .lcout(\dron_frame_decoder_1.state_ns_0_i_a2_0_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNIFJ1J_3_LC_7_10_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIFJ1J_3_LC_7_10_5 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIFJ1J_3_LC_7_10_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Commands_frame_decoder.state_RNIFJ1J_3_LC_7_10_5  (
            .in0(_gnd_net_),
            .in1(N__23757),
            .in2(_gnd_net_),
            .in3(N__27039),
            .lcout(\Commands_frame_decoder.source_CH2data_1_sqmuxa ),
            .ltout(\Commands_frame_decoder.source_CH2data_1_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNIC08S_3_LC_7_10_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIC08S_3_LC_7_10_6 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIC08S_3_LC_7_10_6 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \Commands_frame_decoder.state_RNIC08S_3_LC_7_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20586),
            .in3(N__44088),
            .lcout(\Commands_frame_decoder.source_CH2data_1_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_ns_0_i_a2_1_0_3_LC_7_11_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_ns_0_i_a2_1_0_3_LC_7_11_0 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_ns_0_i_a2_1_0_3_LC_7_11_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \dron_frame_decoder_1.state_ns_0_i_a2_1_0_3_LC_7_11_0  (
            .in0(_gnd_net_),
            .in1(N__25090),
            .in2(_gnd_net_),
            .in3(N__25174),
            .lcout(),
            .ltout(\dron_frame_decoder_1.state_ns_0_i_a2_1_0Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_ns_0_i_a2_1_3_LC_7_11_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_ns_0_i_a2_1_3_LC_7_11_1 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_ns_0_i_a2_1_3_LC_7_11_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \dron_frame_decoder_1.state_ns_0_i_a2_1_3_LC_7_11_1  (
            .in0(N__24732),
            .in1(N__25042),
            .in2(N__20583),
            .in3(N__29657),
            .lcout(\dron_frame_decoder_1.state_ns_0_i_a2_1Z0Z_3 ),
            .ltout(\dron_frame_decoder_1.state_ns_0_i_a2_1Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_RNO_0_0_LC_7_11_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNO_0_0_LC_7_11_2 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNO_0_0_LC_7_11_2 .LUT_INIT=16'b1111000010000000;
    LogicCell40 \dron_frame_decoder_1.state_RNO_0_0_LC_7_11_2  (
            .in0(N__22629),
            .in1(N__20580),
            .in2(N__20574),
            .in3(N__20565),
            .lcout(),
            .ltout(\dron_frame_decoder_1.state_RNO_0Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_0_LC_7_11_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_0_LC_7_11_3 .SEQ_MODE=4'b1001;
    defparam \dron_frame_decoder_1.state_0_LC_7_11_3 .LUT_INIT=16'b0000001100000001;
    LogicCell40 \dron_frame_decoder_1.state_0_LC_7_11_3  (
            .in0(N__22530),
            .in1(N__20658),
            .in2(N__20571),
            .in3(N__22648),
            .lcout(\dron_frame_decoder_1.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47421),
            .ce(),
            .sr(N__43804));
    defparam \dron_frame_decoder_1.state_ns_0_i_a2_0_0_1_1_LC_7_11_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_ns_0_i_a2_0_0_1_1_LC_7_11_4 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_ns_0_i_a2_0_0_1_1_LC_7_11_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \dron_frame_decoder_1.state_ns_0_i_a2_0_0_1_1_LC_7_11_4  (
            .in0(_gnd_net_),
            .in1(N__25216),
            .in2(_gnd_net_),
            .in3(N__25009),
            .lcout(),
            .ltout(\dron_frame_decoder_1.state_ns_0_i_a2_0_0_1Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_RNIN9KQ1_0_LC_7_11_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNIN9KQ1_0_LC_7_11_5 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNIN9KQ1_0_LC_7_11_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \dron_frame_decoder_1.state_RNIN9KQ1_0_LC_7_11_5  (
            .in0(N__25138),
            .in1(N__22647),
            .in2(N__20568),
            .in3(N__26200),
            .lcout(\dron_frame_decoder_1.state_ns_0_i_a2_0_1 ),
            .ltout(\dron_frame_decoder_1.state_ns_0_i_a2_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_1_LC_7_11_6 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_1_LC_7_11_6 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.state_1_LC_7_11_6 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \dron_frame_decoder_1.state_1_LC_7_11_6  (
            .in0(N__20682),
            .in1(N__20555),
            .in2(N__20541),
            .in3(N__22529),
            .lcout(\dron_frame_decoder_1.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47421),
            .ce(),
            .sr(N__43804));
    defparam \pid_alt.un9lto29_i_a2_7_c_RNO_LC_7_12_1 .C_ON=1'b0;
    defparam \pid_alt.un9lto29_i_a2_7_c_RNO_LC_7_12_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un9lto29_i_a2_7_c_RNO_LC_7_12_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \pid_alt.un9lto29_i_a2_7_c_RNO_LC_7_12_1  (
            .in0(_gnd_net_),
            .in1(N__22739),
            .in2(_gnd_net_),
            .in3(N__22566),
            .lcout(\pid_alt.N_232_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_p_reg_esr_RNIFPN33_0_LC_7_12_3 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_RNIFPN33_0_LC_7_12_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_p_reg_esr_RNIFPN33_0_LC_7_12_3 .LUT_INIT=16'b0101010101100110;
    LogicCell40 \pid_alt.error_p_reg_esr_RNIFPN33_0_LC_7_12_3  (
            .in0(N__20796),
            .in1(N__20787),
            .in2(N__30102),
            .in3(N__20738),
            .lcout(\pid_alt.error_p_reg_esr_RNIFPN33Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNO_0_12_LC_7_12_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNO_0_12_LC_7_12_4 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNO_0_12_LC_7_12_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Commands_frame_decoder.state_RNO_0_12_LC_7_12_4  (
            .in0(_gnd_net_),
            .in1(N__23708),
            .in2(_gnd_net_),
            .in3(N__27045),
            .lcout(\Commands_frame_decoder.N_354 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNIM4TM_16_LC_7_12_5 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNIM4TM_16_LC_7_12_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNIM4TM_16_LC_7_12_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_alt.pid_prereg_esr_RNIM4TM_16_LC_7_12_5  (
            .in0(N__20910),
            .in1(N__20952),
            .in2(N__20868),
            .in3(N__20991),
            .lcout(\pid_alt.un9lto29_i_a2_3_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_RNO_1_0_LC_7_12_6 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNO_1_0_LC_7_12_6 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNO_1_0_LC_7_12_6 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \dron_frame_decoder_1.state_RNO_1_0_LC_7_12_6  (
            .in0(N__22650),
            .in1(N__29713),
            .in2(N__20681),
            .in3(N__29667),
            .lcout(\dron_frame_decoder_1.state_RNO_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un1_pid_prereg_un1_pid_prereg_0_cry_0_c_THRU_CRY_0_LC_7_13_0 .C_ON=1'b1;
    defparam \pid_alt.un1_pid_prereg_un1_pid_prereg_0_cry_0_c_THRU_CRY_0_LC_7_13_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un1_pid_prereg_un1_pid_prereg_0_cry_0_c_THRU_CRY_0_LC_7_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_alt.un1_pid_prereg_un1_pid_prereg_0_cry_0_c_THRU_CRY_0_LC_7_13_0  (
            .in0(_gnd_net_),
            .in1(N__20642),
            .in2(N__20649),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_13_0_),
            .carryout(\pid_alt.un1_pid_prereg_un1_pid_prereg_0_cry_0_c_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_0_LC_7_13_1 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_0_LC_7_13_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_0_LC_7_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_0_LC_7_13_1  (
            .in0(_gnd_net_),
            .in1(N__20622),
            .in2(N__30137),
            .in3(N__20610),
            .lcout(\pid_alt.pid_preregZ0Z_0 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_un1_pid_prereg_0_cry_0_c_THRU_CO ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_0 ),
            .clk(N__47397),
            .ce(N__33600),
            .sr(N__43810));
    defparam \pid_alt.pid_prereg_esr_1_LC_7_13_2 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_1_LC_7_13_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_1_LC_7_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_1_LC_7_13_2  (
            .in0(_gnd_net_),
            .in1(N__20607),
            .in2(N__30101),
            .in3(N__20601),
            .lcout(\pid_alt.pid_preregZ0Z_1 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_0 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_1 ),
            .clk(N__47397),
            .ce(N__33600),
            .sr(N__43810));
    defparam \pid_alt.pid_prereg_esr_2_LC_7_13_3 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_2_LC_7_13_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_2_LC_7_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_2_LC_7_13_3  (
            .in0(_gnd_net_),
            .in1(N__20598),
            .in2(N__30035),
            .in3(N__20589),
            .lcout(\pid_alt.pid_preregZ0Z_2 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_1 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_2 ),
            .clk(N__47397),
            .ce(N__33600),
            .sr(N__43810));
    defparam \pid_alt.pid_prereg_esr_3_LC_7_13_4 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_3_LC_7_13_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_3_LC_7_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_3_LC_7_13_4  (
            .in0(_gnd_net_),
            .in1(N__20853),
            .in2(N__29996),
            .in3(N__20844),
            .lcout(\pid_alt.pid_preregZ0Z_3 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_2 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_3 ),
            .clk(N__47397),
            .ce(N__33600),
            .sr(N__43810));
    defparam \pid_alt.pid_prereg_esr_4_LC_7_13_5 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_4_LC_7_13_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_4_LC_7_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_4_LC_7_13_5  (
            .in0(_gnd_net_),
            .in1(N__26114),
            .in2(N__26091),
            .in3(N__20841),
            .lcout(\pid_alt.pid_preregZ0Z_4 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_3 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_4 ),
            .clk(N__47397),
            .ce(N__33600),
            .sr(N__43810));
    defparam \pid_alt.pid_prereg_esr_5_LC_7_13_6 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_5_LC_7_13_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_5_LC_7_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_5_LC_7_13_6  (
            .in0(_gnd_net_),
            .in1(N__22668),
            .in2(N__26049),
            .in3(N__20838),
            .lcout(\pid_alt.pid_preregZ0Z_5 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_4 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_5 ),
            .clk(N__47397),
            .ce(N__33600),
            .sr(N__43810));
    defparam \pid_alt.pid_prereg_esr_6_LC_7_13_7 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_6_LC_7_13_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_6_LC_7_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_6_LC_7_13_7  (
            .in0(_gnd_net_),
            .in1(N__22698),
            .in2(N__22692),
            .in3(N__20835),
            .lcout(\pid_alt.pid_preregZ0Z_6 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_5 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_6 ),
            .clk(N__47397),
            .ce(N__33600),
            .sr(N__43810));
    defparam \pid_alt.pid_prereg_esr_7_LC_7_14_0 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_7_LC_7_14_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_7_LC_7_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_7_LC_7_14_0  (
            .in0(_gnd_net_),
            .in1(N__22752),
            .in2(N__22772),
            .in3(N__20832),
            .lcout(\pid_alt.pid_preregZ0Z_7 ),
            .ltout(),
            .carryin(bfn_7_14_0_),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_7 ),
            .clk(N__47383),
            .ce(N__33603),
            .sr(N__43816));
    defparam \pid_alt.pid_prereg_esr_8_LC_7_14_1 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_8_LC_7_14_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_8_LC_7_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_8_LC_7_14_1  (
            .in0(_gnd_net_),
            .in1(N__20829),
            .in2(N__26315),
            .in3(N__20817),
            .lcout(\pid_alt.pid_preregZ0Z_8 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_7 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_8 ),
            .clk(N__47383),
            .ce(N__33603),
            .sr(N__43816));
    defparam \pid_alt.pid_prereg_esr_9_LC_7_14_2 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_9_LC_7_14_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_9_LC_7_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_9_LC_7_14_2  (
            .in0(_gnd_net_),
            .in1(N__22779),
            .in2(N__22808),
            .in3(N__20814),
            .lcout(\pid_alt.pid_preregZ0Z_9 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_8 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_9 ),
            .clk(N__47383),
            .ce(N__33603),
            .sr(N__43816));
    defparam \pid_alt.pid_prereg_esr_10_LC_7_14_3 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_10_LC_7_14_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_10_LC_7_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_10_LC_7_14_3  (
            .in0(_gnd_net_),
            .in1(N__22980),
            .in2(N__22902),
            .in3(N__20811),
            .lcout(\pid_alt.pid_preregZ0Z_10 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_9 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_10 ),
            .clk(N__47383),
            .ce(N__33603),
            .sr(N__43816));
    defparam \pid_alt.pid_prereg_esr_11_LC_7_14_4 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_11_LC_7_14_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_11_LC_7_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_11_LC_7_14_4  (
            .in0(_gnd_net_),
            .in1(N__20808),
            .in2(N__23081),
            .in3(N__20799),
            .lcout(\pid_alt.pid_preregZ0Z_11 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_10 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_11 ),
            .clk(N__47383),
            .ce(N__33603),
            .sr(N__43816));
    defparam \pid_alt.pid_prereg_esr_12_LC_7_14_5 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_12_LC_7_14_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_12_LC_7_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_12_LC_7_14_5  (
            .in0(_gnd_net_),
            .in1(N__21165),
            .in2(N__21156),
            .in3(N__21144),
            .lcout(\pid_alt.pid_preregZ0Z_12 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_11 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_12 ),
            .clk(N__47383),
            .ce(N__33603),
            .sr(N__43816));
    defparam \pid_alt.pid_prereg_esr_13_LC_7_14_6 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_13_LC_7_14_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_13_LC_7_14_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_13_LC_7_14_6  (
            .in0(_gnd_net_),
            .in1(N__21141),
            .in2(N__21126),
            .in3(N__21105),
            .lcout(\pid_alt.pid_preregZ0Z_13 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_12 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_13 ),
            .clk(N__47383),
            .ce(N__33603),
            .sr(N__43816));
    defparam \pid_alt.pid_prereg_esr_14_LC_7_14_7 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_14_LC_7_14_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_14_LC_7_14_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_14_LC_7_14_7  (
            .in0(_gnd_net_),
            .in1(N__21102),
            .in2(N__21090),
            .in3(N__21066),
            .lcout(\pid_alt.pid_preregZ0Z_14 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_13 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_14 ),
            .clk(N__47383),
            .ce(N__33603),
            .sr(N__43816));
    defparam \pid_alt.pid_prereg_esr_15_LC_7_15_0 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_15_LC_7_15_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_15_LC_7_15_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_15_LC_7_15_0  (
            .in0(_gnd_net_),
            .in1(N__21063),
            .in2(N__21051),
            .in3(N__21027),
            .lcout(\pid_alt.pid_preregZ0Z_15 ),
            .ltout(),
            .carryin(bfn_7_15_0_),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_15 ),
            .clk(N__47370),
            .ce(N__33607),
            .sr(N__43820));
    defparam \pid_alt.pid_prereg_esr_16_LC_7_15_1 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_16_LC_7_15_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_16_LC_7_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_16_LC_7_15_1  (
            .in0(_gnd_net_),
            .in1(N__21024),
            .in2(N__21015),
            .in3(N__20982),
            .lcout(\pid_alt.pid_preregZ0Z_16 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_15 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_16 ),
            .clk(N__47370),
            .ce(N__33607),
            .sr(N__43820));
    defparam \pid_alt.pid_prereg_esr_17_LC_7_15_2 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_17_LC_7_15_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_17_LC_7_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_17_LC_7_15_2  (
            .in0(_gnd_net_),
            .in1(N__20979),
            .in2(N__20970),
            .in3(N__20943),
            .lcout(\pid_alt.pid_preregZ0Z_17 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_16 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_17 ),
            .clk(N__47370),
            .ce(N__33607),
            .sr(N__43820));
    defparam \pid_alt.pid_prereg_esr_18_LC_7_15_3 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_18_LC_7_15_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_18_LC_7_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_18_LC_7_15_3  (
            .in0(_gnd_net_),
            .in1(N__20940),
            .in2(N__20931),
            .in3(N__20901),
            .lcout(\pid_alt.pid_preregZ0Z_18 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_17 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_18 ),
            .clk(N__47370),
            .ce(N__33607),
            .sr(N__43820));
    defparam \pid_alt.pid_prereg_esr_19_LC_7_15_4 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_19_LC_7_15_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_19_LC_7_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_19_LC_7_15_4  (
            .in0(_gnd_net_),
            .in1(N__20898),
            .in2(N__20889),
            .in3(N__20856),
            .lcout(\pid_alt.pid_preregZ0Z_19 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_18 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_19 ),
            .clk(N__47370),
            .ce(N__33607),
            .sr(N__43820));
    defparam \pid_alt.pid_prereg_esr_20_LC_7_15_5 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_20_LC_7_15_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_20_LC_7_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_20_LC_7_15_5  (
            .in0(_gnd_net_),
            .in1(N__21237),
            .in2(N__21228),
            .in3(N__21207),
            .lcout(\pid_alt.pid_preregZ0Z_20 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_19 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_20 ),
            .clk(N__47370),
            .ce(N__33607),
            .sr(N__43820));
    defparam \pid_alt.pid_prereg_esr_21_LC_7_15_6 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_21_LC_7_15_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_21_LC_7_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_21_LC_7_15_6  (
            .in0(_gnd_net_),
            .in1(N__23256),
            .in2(N__23292),
            .in3(N__21204),
            .lcout(\pid_alt.pid_preregZ0Z_21 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_20 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_21 ),
            .clk(N__47370),
            .ce(N__33607),
            .sr(N__43820));
    defparam \pid_alt.pid_prereg_esr_22_LC_7_15_7 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_22_LC_7_15_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_22_LC_7_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_22_LC_7_15_7  (
            .in0(_gnd_net_),
            .in1(N__22998),
            .in2(N__23010),
            .in3(N__21201),
            .lcout(\pid_alt.pid_preregZ0Z_22 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_21 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_22 ),
            .clk(N__47370),
            .ce(N__33607),
            .sr(N__43820));
    defparam \pid_alt.pid_prereg_esr_23_LC_7_16_0 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_23_LC_7_16_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_23_LC_7_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_23_LC_7_16_0  (
            .in0(_gnd_net_),
            .in1(N__23045),
            .in2(N__21198),
            .in3(N__21183),
            .lcout(\pid_alt.pid_preregZ0Z_23 ),
            .ltout(),
            .carryin(bfn_7_16_0_),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_23 ),
            .clk(N__47357),
            .ce(N__33612),
            .sr(N__43826));
    defparam \pid_alt.pid_prereg_esr_24_LC_7_16_1 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_24_LC_7_16_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_24_LC_7_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_24_LC_7_16_1  (
            .in0(_gnd_net_),
            .in1(N__26243),
            .in2(N__26220),
            .in3(N__21180),
            .lcout(\pid_alt.pid_preregZ0Z_24 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_23 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_24 ),
            .clk(N__47357),
            .ce(N__33612),
            .sr(N__43826));
    defparam \pid_alt.pid_prereg_esr_25_LC_7_16_2 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_25_LC_7_16_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_25_LC_7_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_25_LC_7_16_2  (
            .in0(_gnd_net_),
            .in1(N__24239),
            .in2(N__24324),
            .in3(N__21177),
            .lcout(\pid_alt.pid_preregZ0Z_25 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_24 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_25 ),
            .clk(N__47357),
            .ce(N__33612),
            .sr(N__43826));
    defparam \pid_alt.pid_prereg_esr_26_LC_7_16_3 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_26_LC_7_16_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_26_LC_7_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_26_LC_7_16_3  (
            .in0(_gnd_net_),
            .in1(N__24260),
            .in2(N__24384),
            .in3(N__21174),
            .lcout(\pid_alt.pid_preregZ0Z_26 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_25 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_26 ),
            .clk(N__47357),
            .ce(N__33612),
            .sr(N__43826));
    defparam \pid_alt.pid_prereg_esr_27_LC_7_16_4 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_27_LC_7_16_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_27_LC_7_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_27_LC_7_16_4  (
            .in0(_gnd_net_),
            .in1(N__21279),
            .in2(N__24347),
            .in3(N__21171),
            .lcout(\pid_alt.pid_preregZ0Z_27 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_26 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_27 ),
            .clk(N__47357),
            .ce(N__33612),
            .sr(N__43826));
    defparam \pid_alt.pid_prereg_esr_28_LC_7_16_5 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_28_LC_7_16_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_28_LC_7_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_28_LC_7_16_5  (
            .in0(_gnd_net_),
            .in1(N__21270),
            .in2(N__21246),
            .in3(N__21168),
            .lcout(\pid_alt.pid_preregZ0Z_28 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_27 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_28 ),
            .clk(N__47357),
            .ce(N__33612),
            .sr(N__43826));
    defparam \pid_alt.pid_prereg_esr_29_LC_7_16_6 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_29_LC_7_16_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_29_LC_7_16_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_29_LC_7_16_6  (
            .in0(_gnd_net_),
            .in1(N__21990),
            .in2(N__22068),
            .in3(N__21285),
            .lcout(\pid_alt.pid_preregZ0Z_29 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_28 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_29 ),
            .clk(N__47357),
            .ce(N__33612),
            .sr(N__43826));
    defparam \pid_alt.pid_prereg_esr_30_LC_7_16_7 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_30_LC_7_16_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_30_LC_7_16_7 .LUT_INIT=16'b1000000101111110;
    LogicCell40 \pid_alt.pid_prereg_esr_30_LC_7_16_7  (
            .in0(N__22015),
            .in1(N__30720),
            .in2(N__22053),
            .in3(N__21282),
            .lcout(\pid_alt.pid_preregZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47357),
            .ce(N__33612),
            .sr(N__43826));
    defparam \pid_alt.error_d_reg_prev_esr_RNI8JT34_26_LC_7_17_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI8JT34_26_LC_7_17_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI8JT34_26_LC_7_17_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI8JT34_26_LC_7_17_0  (
            .in0(N__22008),
            .in1(N__21260),
            .in2(N__24351),
            .in3(N__30718),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI8JT34Z0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNISSKM_26_LC_7_17_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNISSKM_26_LC_7_17_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNISSKM_26_LC_7_17_1 .LUT_INIT=16'b1101110101000100;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNISSKM_26_LC_7_17_1  (
            .in0(N__23153),
            .in1(N__23138),
            .in2(_gnd_net_),
            .in3(N__24635),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNISSKMZ0Z_26 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNISSKMZ0Z_26_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIMRU12_26_LC_7_17_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIMRU12_26_LC_7_17_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIMRU12_26_LC_7_17_2 .LUT_INIT=16'b1111101010100000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIMRU12_26_LC_7_17_2  (
            .in0(N__22009),
            .in1(_gnd_net_),
            .in2(N__21273),
            .in3(N__30717),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIMRU12Z0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_26_LC_7_17_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_26_LC_7_17_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_26_LC_7_17_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_26_LC_7_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23139),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47345),
            .ce(N__33616),
            .sr(N__43836));
    defparam \pid_alt.error_d_reg_prev_esr_RNIUUKM_0_27_LC_7_17_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIUUKM_0_27_LC_7_17_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIUUKM_0_27_LC_7_17_4 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIUUKM_0_27_LC_7_17_4  (
            .in0(N__24636),
            .in1(N__21494),
            .in2(_gnd_net_),
            .in3(N__21523),
            .lcout(\pid_alt.un1_pid_prereg_296_1 ),
            .ltout(\pid_alt.un1_pid_prereg_296_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIKQJO2_26_LC_7_17_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIKQJO2_26_LC_7_17_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIKQJO2_26_LC_7_17_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIKQJO2_26_LC_7_17_5  (
            .in0(N__30719),
            .in1(N__21261),
            .in2(N__21249),
            .in3(N__22047),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIKQJO2Z0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_27_LC_7_17_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_27_LC_7_17_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_27_LC_7_17_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_27_LC_7_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21525),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47345),
            .ce(N__33616),
            .sr(N__43836));
    defparam \pid_alt.error_d_reg_prev_esr_RNIUUKM_27_LC_7_17_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIUUKM_27_LC_7_17_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIUUKM_27_LC_7_17_7 .LUT_INIT=16'b1010111100001010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIUUKM_27_LC_7_17_7  (
            .in0(N__21524),
            .in1(_gnd_net_),
            .in2(N__21498),
            .in3(N__24637),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIUUKMZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_CH1data_1_LC_7_18_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH1data_1_LC_7_18_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH1data_1_LC_7_18_2 .LUT_INIT=16'b0100111101000000;
    LogicCell40 \Commands_frame_decoder.source_CH1data_1_LC_7_18_2  (
            .in0(N__24099),
            .in1(N__45186),
            .in2(N__31849),
            .in3(N__21977),
            .lcout(alt_command_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47329),
            .ce(),
            .sr(N__43842));
    defparam \Commands_frame_decoder.source_CH1data_2_LC_7_18_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH1data_2_LC_7_18_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH1data_2_LC_7_18_3 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \Commands_frame_decoder.source_CH1data_2_LC_7_18_3  (
            .in0(N__36888),
            .in1(N__24100),
            .in2(N__21909),
            .in3(N__31842),
            .lcout(alt_command_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47329),
            .ce(),
            .sr(N__43842));
    defparam \Commands_frame_decoder.source_CH1data_3_LC_7_18_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH1data_3_LC_7_18_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH1data_3_LC_7_18_4 .LUT_INIT=16'b0100111101000000;
    LogicCell40 \Commands_frame_decoder.source_CH1data_3_LC_7_18_4  (
            .in0(N__24101),
            .in1(N__43354),
            .in2(N__31850),
            .in3(N__21849),
            .lcout(alt_command_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47329),
            .ce(),
            .sr(N__43842));
    defparam \pid_alt.error_cry_0_c_LC_7_19_0 .C_ON=1'b1;
    defparam \pid_alt.error_cry_0_c_LC_7_19_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_0_c_LC_7_19_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_alt.error_cry_0_c_LC_7_19_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23244),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_19_0_),
            .carryout(\pid_alt.error_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_0_c_RNI1N2F_LC_7_19_1 .C_ON=1'b1;
    defparam \pid_alt.error_cry_0_c_RNI1N2F_LC_7_19_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_0_c_RNI1N2F_LC_7_19_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pid_alt.error_cry_0_c_RNI1N2F_LC_7_19_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23436),
            .in3(N__21438),
            .lcout(\pid_alt.error_1 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_0 ),
            .carryout(\pid_alt.error_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_1_c_RNI3Q3F_LC_7_19_2 .C_ON=1'b1;
    defparam \pid_alt.error_cry_1_c_RNI3Q3F_LC_7_19_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_1_c_RNI3Q3F_LC_7_19_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pid_alt.error_cry_1_c_RNI3Q3F_LC_7_19_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23400),
            .in3(N__21393),
            .lcout(\pid_alt.error_2 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_1 ),
            .carryout(\pid_alt.error_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_2_c_RNI5T4F_LC_7_19_3 .C_ON=1'b1;
    defparam \pid_alt.error_cry_2_c_RNI5T4F_LC_7_19_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_2_c_RNI5T4F_LC_7_19_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pid_alt.error_cry_2_c_RNI5T4F_LC_7_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23229),
            .in3(N__21342),
            .lcout(\pid_alt.error_3 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_2 ),
            .carryout(\pid_alt.error_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_3_c_RNIKE1T_LC_7_19_4 .C_ON=1'b1;
    defparam \pid_alt.error_cry_3_c_RNIKE1T_LC_7_19_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_3_c_RNIKE1T_LC_7_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_cry_3_c_RNIKE1T_LC_7_19_4  (
            .in0(_gnd_net_),
            .in1(N__23364),
            .in2(N__24810),
            .in3(N__21288),
            .lcout(\pid_alt.error_4 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_3 ),
            .carryout(\pid_alt.error_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_4_c_RNINI2T_LC_7_19_5 .C_ON=1'b1;
    defparam \pid_alt.error_cry_4_c_RNINI2T_LC_7_19_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_4_c_RNINI2T_LC_7_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_cry_4_c_RNINI2T_LC_7_19_5  (
            .in0(_gnd_net_),
            .in1(N__21978),
            .in2(N__24792),
            .in3(N__21912),
            .lcout(\pid_alt.error_5 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_4 ),
            .carryout(\pid_alt.error_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_5_c_RNIQM3T_LC_7_19_6 .C_ON=1'b1;
    defparam \pid_alt.error_cry_5_c_RNIQM3T_LC_7_19_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_5_c_RNIQM3T_LC_7_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_cry_5_c_RNIQM3T_LC_7_19_6  (
            .in0(_gnd_net_),
            .in1(N__24774),
            .in2(N__21908),
            .in3(N__21852),
            .lcout(\pid_alt.error_6 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_5 ),
            .carryout(\pid_alt.error_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_6_c_RNITQ4T_LC_7_19_7 .C_ON=1'b1;
    defparam \pid_alt.error_cry_6_c_RNITQ4T_LC_7_19_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_6_c_RNITQ4T_LC_7_19_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_cry_6_c_RNITQ4T_LC_7_19_7  (
            .in0(_gnd_net_),
            .in1(N__21848),
            .in2(N__24759),
            .in3(N__21783),
            .lcout(\pid_alt.error_7 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_6 ),
            .carryout(\pid_alt.error_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_7_c_RNI9LEM_LC_7_20_0 .C_ON=1'b1;
    defparam \pid_alt.error_cry_7_c_RNI9LEM_LC_7_20_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_7_c_RNI9LEM_LC_7_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_cry_7_c_RNI9LEM_LC_7_20_0  (
            .in0(_gnd_net_),
            .in1(N__22098),
            .in2(N__24747),
            .in3(N__21729),
            .lcout(\pid_alt.error_8 ),
            .ltout(),
            .carryin(bfn_7_20_0_),
            .carryout(\pid_alt.error_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_8_c_RNICPFM_LC_7_20_1 .C_ON=1'b1;
    defparam \pid_alt.error_cry_8_c_RNICPFM_LC_7_20_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_8_c_RNICPFM_LC_7_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_cry_8_c_RNICPFM_LC_7_20_1  (
            .in0(_gnd_net_),
            .in1(N__22092),
            .in2(N__23373),
            .in3(N__21675),
            .lcout(\pid_alt.error_9 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_8 ),
            .carryout(\pid_alt.error_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_9_c_RNIMMUJ_LC_7_20_2 .C_ON=1'b1;
    defparam \pid_alt.error_cry_9_c_RNIMMUJ_LC_7_20_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_9_c_RNIMMUJ_LC_7_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_cry_9_c_RNIMMUJ_LC_7_20_2  (
            .in0(_gnd_net_),
            .in1(N__22083),
            .in2(N__23220),
            .in3(N__21630),
            .lcout(\pid_alt.error_10 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_9 ),
            .carryout(\pid_alt.error_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_10_c_RNI0SDO_LC_7_20_3 .C_ON=1'b1;
    defparam \pid_alt.error_cry_10_c_RNI0SDO_LC_7_20_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_10_c_RNI0SDO_LC_7_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_cry_10_c_RNI0SDO_LC_7_20_3  (
            .in0(_gnd_net_),
            .in1(N__22074),
            .in2(N__23211),
            .in3(N__21582),
            .lcout(\pid_alt.error_11 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_10 ),
            .carryout(\pid_alt.error_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_11_c_RNI5JAH_LC_7_20_4 .C_ON=1'b1;
    defparam \pid_alt.error_cry_11_c_RNI5JAH_LC_7_20_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_11_c_RNI5JAH_LC_7_20_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pid_alt.error_cry_11_c_RNI5JAH_LC_7_20_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23427),
            .in3(N__21528),
            .lcout(\pid_alt.error_12 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_11 ),
            .carryout(\pid_alt.error_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_12_c_RNI7MBH_LC_7_20_5 .C_ON=1'b1;
    defparam \pid_alt.error_cry_12_c_RNI7MBH_LC_7_20_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_12_c_RNI7MBH_LC_7_20_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pid_alt.error_cry_12_c_RNI7MBH_LC_7_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23418),
            .in3(N__22209),
            .lcout(\pid_alt.error_13 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_12 ),
            .carryout(\pid_alt.error_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_13_c_RNI9PCH_LC_7_20_6 .C_ON=1'b1;
    defparam \pid_alt.error_cry_13_c_RNI9PCH_LC_7_20_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_13_c_RNI9PCH_LC_7_20_6 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pid_alt.error_cry_13_c_RNI9PCH_LC_7_20_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23409),
            .in3(N__22155),
            .lcout(\pid_alt.error_14 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_13 ),
            .carryout(\pid_alt.error_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_14_c_RNIBSDH_LC_7_20_7 .C_ON=1'b0;
    defparam \pid_alt.error_cry_14_c_RNIBSDH_LC_7_20_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_14_c_RNIBSDH_LC_7_20_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \pid_alt.error_cry_14_c_RNIBSDH_LC_7_20_7  (
            .in0(_gnd_net_),
            .in1(N__25062),
            .in2(_gnd_net_),
            .in3(N__22152),
            .lcout(\pid_alt.error_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_CH1data_esr_4_LC_7_21_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH1data_esr_4_LC_7_21_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH1data_esr_4_LC_7_21_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH1data_esr_4_LC_7_21_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45362),
            .lcout(alt_command_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47294),
            .ce(N__31791),
            .sr(N__43864));
    defparam \Commands_frame_decoder.source_CH1data_esr_5_LC_7_21_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH1data_esr_5_LC_7_21_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH1data_esr_5_LC_7_21_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH1data_esr_5_LC_7_21_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44290),
            .lcout(alt_command_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47294),
            .ce(N__31791),
            .sr(N__43864));
    defparam \Commands_frame_decoder.source_CH1data_esr_6_LC_7_21_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH1data_esr_6_LC_7_21_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH1data_esr_6_LC_7_21_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH1data_esr_6_LC_7_21_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33441),
            .lcout(alt_command_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47294),
            .ce(N__31791),
            .sr(N__43864));
    defparam \Commands_frame_decoder.source_CH1data_esr_7_LC_7_21_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH1data_esr_7_LC_7_21_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH1data_esr_7_LC_7_21_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH1data_esr_7_LC_7_21_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45014),
            .lcout(alt_command_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47294),
            .ce(N__31791),
            .sr(N__43864));
    defparam \pid_alt.error_d_reg_prev_esr_RNIOTU12_27_LC_7_22_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIOTU12_27_LC_7_22_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIOTU12_27_LC_7_22_7 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIOTU12_27_LC_7_22_7  (
            .in0(N__22052),
            .in1(N__22023),
            .in2(_gnd_net_),
            .in3(N__30706),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIOTU12Z0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIOTU12_0_27_LC_7_23_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIOTU12_0_27_LC_7_23_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIOTU12_0_27_LC_7_23_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIOTU12_0_27_LC_7_23_2  (
            .in0(N__22051),
            .in1(N__22022),
            .in2(_gnd_net_),
            .in3(N__30651),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIOTU12_0Z0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.state_RNICP2N1_0_LC_7_29_0 .C_ON=1'b0;
    defparam \pid_alt.state_RNICP2N1_0_LC_7_29_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.state_RNICP2N1_0_LC_7_29_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \pid_alt.state_RNICP2N1_0_LC_7_29_0  (
            .in0(_gnd_net_),
            .in1(N__24135),
            .in2(_gnd_net_),
            .in3(N__46674),
            .lcout(\pid_alt.N_410_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone_sync.aux_2__0__0_LC_8_4_4 .C_ON=1'b0;
    defparam \uart_drone_sync.aux_2__0__0_LC_8_4_4 .SEQ_MODE=4'b1000;
    defparam \uart_drone_sync.aux_2__0__0_LC_8_4_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone_sync.aux_2__0__0_LC_8_4_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22281),
            .lcout(\uart_drone_sync.aux_2__0__0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47469),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone_sync.aux_1__0__0_LC_8_4_5 .C_ON=1'b0;
    defparam \uart_drone_sync.aux_1__0__0_LC_8_4_5 .SEQ_MODE=4'b1000;
    defparam \uart_drone_sync.aux_1__0__0_LC_8_4_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone_sync.aux_1__0__0_LC_8_4_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22266),
            .lcout(\uart_drone_sync.aux_1__0__0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47469),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone_sync.aux_0__0__0_LC_8_4_6 .C_ON=1'b0;
    defparam \uart_drone_sync.aux_0__0__0_LC_8_4_6 .SEQ_MODE=4'b1000;
    defparam \uart_drone_sync.aux_0__0__0_LC_8_4_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uart_drone_sync.aux_0__0__0_LC_8_4_6  (
            .in0(N__22275),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\uart_drone_sync.aux_0__0__0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47469),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.WDT_RNID7P31_6_LC_8_5_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.WDT_RNID7P31_6_LC_8_5_1 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.WDT_RNID7P31_6_LC_8_5_1 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \Commands_frame_decoder.WDT_RNID7P31_6_LC_8_5_1  (
            .in0(N__23476),
            .in1(N__25406),
            .in2(_gnd_net_),
            .in3(N__25382),
            .lcout(),
            .ltout(\Commands_frame_decoder.WDT8lto13_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.WDT_RNIUG2B4_7_LC_8_5_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.WDT_RNIUG2B4_7_LC_8_5_2 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.WDT_RNIUG2B4_7_LC_8_5_2 .LUT_INIT=16'b0010001100110011;
    LogicCell40 \Commands_frame_decoder.WDT_RNIUG2B4_7_LC_8_5_2  (
            .in0(N__23456),
            .in1(N__22257),
            .in2(N__22260),
            .in3(N__22344),
            .lcout(\Commands_frame_decoder.WDT8lt14_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.WDT_RNI2VDI1_10_LC_8_6_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.WDT_RNI2VDI1_10_LC_8_6_0 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.WDT_RNI2VDI1_10_LC_8_6_0 .LUT_INIT=16'b0101010101010111;
    LogicCell40 \Commands_frame_decoder.WDT_RNI2VDI1_10_LC_8_6_0  (
            .in0(N__25427),
            .in1(N__25405),
            .in2(N__23607),
            .in3(N__25381),
            .lcout(\Commands_frame_decoder.WDT_RNI2VDI1Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.WDT_RNII19A1_0_4_LC_8_6_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.WDT_RNII19A1_0_4_LC_8_6_2 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.WDT_RNII19A1_0_4_LC_8_6_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \Commands_frame_decoder.WDT_RNII19A1_0_4_LC_8_6_2  (
            .in0(N__23647),
            .in1(N__23494),
            .in2(N__23630),
            .in3(N__23512),
            .lcout(),
            .ltout(\Commands_frame_decoder.WDT8lto9_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.WDT_RNII01C2_6_LC_8_6_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.WDT_RNII01C2_6_LC_8_6_3 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.WDT_RNII01C2_6_LC_8_6_3 .LUT_INIT=16'b1110111100000000;
    LogicCell40 \Commands_frame_decoder.WDT_RNII01C2_6_LC_8_6_3  (
            .in0(N__23455),
            .in1(N__23477),
            .in2(N__22251),
            .in3(N__23605),
            .lcout(),
            .ltout(\Commands_frame_decoder.WDT8lt12_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.WDT_RNIPJEG6_6_LC_8_6_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.WDT_RNIPJEG6_6_LC_8_6_4 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.WDT_RNIPJEG6_6_LC_8_6_4 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \Commands_frame_decoder.WDT_RNIPJEG6_6_LC_8_6_4  (
            .in0(_gnd_net_),
            .in1(N__22350),
            .in2(N__22353),
            .in3(N__25284),
            .lcout(\Commands_frame_decoder.state_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.preinit_RNIR9JL1_LC_8_6_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.preinit_RNIR9JL1_LC_8_6_5 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.preinit_RNIR9JL1_LC_8_6_5 .LUT_INIT=16'b0000010100000111;
    LogicCell40 \Commands_frame_decoder.preinit_RNIR9JL1_LC_8_6_5  (
            .in0(N__25347),
            .in1(N__25308),
            .in2(N__25275),
            .in3(N__25426),
            .lcout(\Commands_frame_decoder.state_0_sqmuxacf1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.WDT_RNII19A1_4_LC_8_6_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.WDT_RNII19A1_4_LC_8_6_6 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.WDT_RNII19A1_4_LC_8_6_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \Commands_frame_decoder.WDT_RNII19A1_4_LC_8_6_6  (
            .in0(N__23648),
            .in1(N__23495),
            .in2(N__23631),
            .in3(N__23513),
            .lcout(\Commands_frame_decoder.WDT_RNII19A1Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone_sync.aux_3__0__0_LC_8_6_7 .C_ON=1'b0;
    defparam \uart_drone_sync.aux_3__0__0_LC_8_6_7 .SEQ_MODE=4'b1000;
    defparam \uart_drone_sync.aux_3__0__0_LC_8_6_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone_sync.aux_3__0__0_LC_8_6_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22338),
            .lcout(\uart_drone_sync.aux_3__0__0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47457),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_data_valid_2_sqmuxa_i_LC_8_8_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_data_valid_2_sqmuxa_i_LC_8_8_3 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_data_valid_2_sqmuxa_i_LC_8_8_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \dron_frame_decoder_1.source_data_valid_2_sqmuxa_i_LC_8_8_3  (
            .in0(_gnd_net_),
            .in1(N__29668),
            .in2(_gnd_net_),
            .in3(N__44086),
            .lcout(\dron_frame_decoder_1.source_data_valid_2_sqmuxa_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNIJN1J_7_LC_8_8_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIJN1J_7_LC_8_8_4 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIJN1J_7_LC_8_8_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \Commands_frame_decoder.state_RNIJN1J_7_LC_8_8_4  (
            .in0(N__27035),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23678),
            .lcout(\Commands_frame_decoder.source_offset2data_1_sqmuxa ),
            .ltout(\Commands_frame_decoder.source_offset2data_1_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNIG48S_7_LC_8_8_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIG48S_7_LC_8_8_5 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIG48S_7_LC_8_8_5 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \Commands_frame_decoder.state_RNIG48S_7_LC_8_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22299),
            .in3(N__44087),
            .lcout(\Commands_frame_decoder.source_offset2data_1_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNO_2_0_LC_8_8_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNO_2_0_LC_8_8_6 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNO_2_0_LC_8_8_6 .LUT_INIT=16'b0000101000001000;
    LogicCell40 \Commands_frame_decoder.state_RNO_2_0_LC_8_8_6  (
            .in0(N__25359),
            .in1(N__25316),
            .in2(N__27044),
            .in3(N__23663),
            .lcout(),
            .ltout(\Commands_frame_decoder.N_322_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNO_0_0_LC_8_8_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNO_0_0_LC_8_8_7 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNO_0_0_LC_8_8_7 .LUT_INIT=16'b0000001100000000;
    LogicCell40 \Commands_frame_decoder.state_RNO_0_0_LC_8_8_7  (
            .in0(_gnd_net_),
            .in1(N__25238),
            .in2(N__22296),
            .in3(N__25616),
            .lcout(\Commands_frame_decoder.N_327 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNIF38S_6_LC_8_9_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIF38S_6_LC_8_9_0 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIF38S_6_LC_8_9_0 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \Commands_frame_decoder.state_RNIF38S_6_LC_8_9_0  (
            .in0(N__27009),
            .in1(N__25524),
            .in2(_gnd_net_),
            .in3(N__44068),
            .lcout(\Commands_frame_decoder.state_RNIF38SZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNIQRI31_10_LC_8_9_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIQRI31_10_LC_8_9_2 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIQRI31_10_LC_8_9_2 .LUT_INIT=16'b1111111110100000;
    LogicCell40 \Commands_frame_decoder.state_RNIQRI31_10_LC_8_9_2  (
            .in0(N__27010),
            .in1(_gnd_net_),
            .in2(N__23777),
            .in3(N__44067),
            .lcout(\Commands_frame_decoder.state_RNIQRI31Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_12_LC_8_9_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_12_LC_8_9_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_12_LC_8_9_5 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \Commands_frame_decoder.state_12_LC_8_9_5  (
            .in0(N__24863),
            .in1(N__26448),
            .in2(N__22431),
            .in3(N__26466),
            .lcout(\Commands_frame_decoder.stateZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47431),
            .ce(),
            .sr(N__43801));
    defparam \Commands_frame_decoder.state_8_LC_8_9_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_8_LC_8_9_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_8_LC_8_9_6 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \Commands_frame_decoder.state_8_LC_8_9_6  (
            .in0(N__22413),
            .in1(N__22419),
            .in2(_gnd_net_),
            .in3(N__24862),
            .lcout(\Commands_frame_decoder.stateZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47431),
            .ce(),
            .sr(N__43801));
    defparam \Commands_frame_decoder.state_RNIKO1J_8_LC_8_9_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIKO1J_8_LC_8_9_7 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIKO1J_8_LC_8_9_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Commands_frame_decoder.state_RNIKO1J_8_LC_8_9_7  (
            .in0(_gnd_net_),
            .in1(N__22412),
            .in2(_gnd_net_),
            .in3(N__27008),
            .lcout(\Commands_frame_decoder.source_offset3data_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_RNI0TLI1_5_LC_8_10_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNI0TLI1_5_LC_8_10_0 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNI0TLI1_5_LC_8_10_0 .LUT_INIT=16'b1111111100000100;
    LogicCell40 \dron_frame_decoder_1.state_RNI0TLI1_5_LC_8_10_0  (
            .in0(N__22391),
            .in1(N__29705),
            .in2(N__22404),
            .in3(N__44082),
            .lcout(\dron_frame_decoder_1.N_392_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_RNI6P6K_4_LC_8_10_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNI6P6K_4_LC_8_10_1 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNI6P6K_4_LC_8_10_1 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \dron_frame_decoder_1.state_RNI6P6K_4_LC_8_10_1  (
            .in0(_gnd_net_),
            .in1(N__29642),
            .in2(_gnd_net_),
            .in3(N__22366),
            .lcout(\dron_frame_decoder_1.un1_sink_data_valid_5_i_0 ),
            .ltout(\dron_frame_decoder_1.un1_sink_data_valid_5_i_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_RNI3T3K1_7_LC_8_10_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNI3T3K1_7_LC_8_10_2 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNI3T3K1_7_LC_8_10_2 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \dron_frame_decoder_1.state_RNI3T3K1_7_LC_8_10_2  (
            .in0(N__22492),
            .in1(N__22389),
            .in2(N__22395),
            .in3(N__29704),
            .lcout(\dron_frame_decoder_1.state_RNI3T3K1Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_4_LC_8_10_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_4_LC_8_10_4 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.state_4_LC_8_10_4 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \dron_frame_decoder_1.state_4_LC_8_10_4  (
            .in0(N__22367),
            .in1(N__22390),
            .in2(N__29663),
            .in3(N__22531),
            .lcout(\dron_frame_decoder_1.stateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47422),
            .ce(),
            .sr(N__43805));
    defparam \dron_frame_decoder_1.state_7_LC_8_10_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_7_LC_8_10_5 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.state_7_LC_8_10_5 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \dron_frame_decoder_1.state_7_LC_8_10_5  (
            .in0(N__22533),
            .in1(N__29643),
            .in2(N__22371),
            .in3(N__22494),
            .lcout(\dron_frame_decoder_1.stateZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47422),
            .ce(),
            .sr(N__43805));
    defparam \uart_drone.data_rdy_LC_8_10_6 .C_ON=1'b0;
    defparam \uart_drone.data_rdy_LC_8_10_6 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_rdy_LC_8_10_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uart_drone.data_rdy_LC_8_10_6  (
            .in0(N__31371),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31647),
            .lcout(uart_drone_data_rdy),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47422),
            .ce(),
            .sr(N__43805));
    defparam \dron_frame_decoder_1.state_6_LC_8_10_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_6_LC_8_10_7 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.state_6_LC_8_10_7 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \dron_frame_decoder_1.state_6_LC_8_10_7  (
            .in0(N__22532),
            .in1(N__22493),
            .in2(N__29714),
            .in3(N__29647),
            .lcout(\dron_frame_decoder_1.stateZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47422),
            .ce(),
            .sr(N__43805));
    defparam \pid_alt.un9lto29_i_a2_0_c_LC_8_11_0 .C_ON=1'b1;
    defparam \pid_alt.un9lto29_i_a2_0_c_LC_8_11_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un9lto29_i_a2_0_c_LC_8_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_alt.un9lto29_i_a2_0_c_LC_8_11_0  (
            .in0(_gnd_net_),
            .in1(N__22584),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_11_0_),
            .carryout(\pid_alt.un9lto29_i_a2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un9lto29_i_a2_1_c_LC_8_11_1 .C_ON=1'b1;
    defparam \pid_alt.un9lto29_i_a2_1_c_LC_8_11_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un9lto29_i_a2_1_c_LC_8_11_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_alt.un9lto29_i_a2_1_c_LC_8_11_1  (
            .in0(_gnd_net_),
            .in1(N__24216),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pid_alt.un9lto29_i_a2 ),
            .carryout(\pid_alt.un9lto29_i_a2_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un9lto29_i_a2_2_c_LC_8_11_2 .C_ON=1'b1;
    defparam \pid_alt.un9lto29_i_a2_2_c_LC_8_11_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un9lto29_i_a2_2_c_LC_8_11_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_alt.un9lto29_i_a2_2_c_LC_8_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23904),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pid_alt.un9lto29_i_a2_0 ),
            .carryout(\pid_alt.un9lto29_i_a2_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un9lto29_i_a2_3_c_LC_8_11_3 .C_ON=1'b1;
    defparam \pid_alt.un9lto29_i_a2_3_c_LC_8_11_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un9lto29_i_a2_3_c_LC_8_11_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_alt.un9lto29_i_a2_3_c_LC_8_11_3  (
            .in0(_gnd_net_),
            .in1(N__22575),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pid_alt.un9lto29_i_a2_1 ),
            .carryout(\pid_alt.un9lto29_i_a2_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un9lto29_i_a2_4_c_LC_8_11_4 .C_ON=1'b1;
    defparam \pid_alt.un9lto29_i_a2_4_c_LC_8_11_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un9lto29_i_a2_4_c_LC_8_11_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_alt.un9lto29_i_a2_4_c_LC_8_11_4  (
            .in0(_gnd_net_),
            .in1(N__23891),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pid_alt.un9lto29_i_a2_2 ),
            .carryout(\pid_alt.un9lto29_i_a2_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un9lto29_i_a2_5_c_LC_8_11_5 .C_ON=1'b1;
    defparam \pid_alt.un9lto29_i_a2_5_c_LC_8_11_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un9lto29_i_a2_5_c_LC_8_11_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_alt.un9lto29_i_a2_5_c_LC_8_11_5  (
            .in0(_gnd_net_),
            .in1(N__23865),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pid_alt.un9lto29_i_a2_3 ),
            .carryout(\pid_alt.un9lto29_i_a2_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un9lto29_i_a2_6_c_LC_8_11_6 .C_ON=1'b1;
    defparam \pid_alt.un9lto29_i_a2_6_c_LC_8_11_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un9lto29_i_a2_6_c_LC_8_11_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_alt.un9lto29_i_a2_6_c_LC_8_11_6  (
            .in0(_gnd_net_),
            .in1(N__23994),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pid_alt.un9lto29_i_a2_4 ),
            .carryout(\pid_alt.un9lto29_i_a2_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un9lto29_i_a2_7_c_LC_8_11_7 .C_ON=1'b1;
    defparam \pid_alt.un9lto29_i_a2_7_c_LC_8_11_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un9lto29_i_a2_7_c_LC_8_11_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_alt.un9lto29_i_a2_7_c_LC_8_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22662),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pid_alt.un9lto29_i_a2_5 ),
            .carryout(\pid_alt.un9lto29_i_a2_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un9lto29_i_a2_7_c_RNIOG6V_LC_8_12_0 .C_ON=1'b0;
    defparam \pid_alt.un9lto29_i_a2_7_c_RNIOG6V_LC_8_12_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un9lto29_i_a2_7_c_RNIOG6V_LC_8_12_0 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \pid_alt.un9lto29_i_a2_7_c_RNIOG6V_LC_8_12_0  (
            .in0(N__33173),
            .in1(N__28043),
            .in2(_gnd_net_),
            .in3(N__22653),
            .lcout(\pid_alt.source_pid_1_sqmuxa_0_a2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.state_0_LC_8_12_1 .C_ON=1'b0;
    defparam \pid_alt.state_0_LC_8_12_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.state_0_LC_8_12_1 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \pid_alt.state_0_LC_8_12_1  (
            .in0(N__24950),
            .in1(N__29601),
            .in2(_gnd_net_),
            .in3(N__33174),
            .lcout(\pid_alt.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47398),
            .ce(),
            .sr(N__43811));
    defparam \dron_frame_decoder_1.state_RNO_2_0_LC_8_12_6 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNO_2_0_LC_8_12_6 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNO_2_0_LC_8_12_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \dron_frame_decoder_1.state_RNO_2_0_LC_8_12_6  (
            .in0(_gnd_net_),
            .in1(N__29712),
            .in2(_gnd_net_),
            .in3(N__22649),
            .lcout(\dron_frame_decoder_1.state_ns_i_i_a2_2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNI2K0N_20_LC_8_13_0 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNI2K0N_20_LC_8_13_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNI2K0N_20_LC_8_13_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_alt.pid_prereg_esr_RNI2K0N_20_LC_8_13_0  (
            .in0(N__22623),
            .in1(N__22614),
            .in2(N__22605),
            .in3(N__22593),
            .lcout(\pid_alt.un9lto29_i_a2_4_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNIDJJA1_1_LC_8_13_1 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNIDJJA1_1_LC_8_13_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNIDJJA1_1_LC_8_13_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_alt.pid_prereg_esr_RNIDJJA1_1_LC_8_13_1  (
            .in0(N__25951),
            .in1(N__23830),
            .in2(N__25886),
            .in3(N__25928),
            .lcout(\pid_alt.source_pid_1_sqmuxa_0_a2_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un9lto29_i_a2_0_c_RNO_LC_8_13_2 .C_ON=1'b0;
    defparam \pid_alt.un9lto29_i_a2_0_c_RNO_LC_8_13_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un9lto29_i_a2_0_c_RNO_LC_8_13_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_alt.un9lto29_i_a2_0_c_RNO_LC_8_13_2  (
            .in0(N__25927),
            .in1(N__25975),
            .in2(N__25958),
            .in3(N__25879),
            .lcout(\pid_alt.source_pid10lt4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un9lto29_i_a2_3_c_RNO_LC_8_13_3 .C_ON=1'b0;
    defparam \pid_alt.un9lto29_i_a2_3_c_RNO_LC_8_13_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un9lto29_i_a2_3_c_RNO_LC_8_13_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_alt.un9lto29_i_a2_3_c_RNO_LC_8_13_3  (
            .in0(N__22716),
            .in1(N__23973),
            .in2(N__22548),
            .in3(N__23829),
            .lcout(\pid_alt.un9lto29_i_a2_2_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNIK4VM_14_LC_8_13_4 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNIK4VM_14_LC_8_13_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNIK4VM_14_LC_8_13_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_alt.pid_prereg_esr_RNIK4VM_14_LC_8_13_4  (
            .in0(N__22565),
            .in1(N__22544),
            .in2(N__22740),
            .in3(N__22715),
            .lcout(\pid_alt.source_pid_1_sqmuxa_0_a2_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.source_pid_1_esr_12_LC_8_13_6 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_esr_12_LC_8_13_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_esr_12_LC_8_13_6 .LUT_INIT=16'b1010001010100000;
    LogicCell40 \pid_alt.source_pid_1_esr_12_LC_8_13_6  (
            .in0(N__23831),
            .in1(N__23972),
            .in2(N__28067),
            .in3(N__23813),
            .lcout(throttle_command_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47384),
            .ce(N__27913),
            .sr(N__27865));
    defparam \pid_alt.source_pid_1_esr_13_LC_8_13_7 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_esr_13_LC_8_13_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_esr_13_LC_8_13_7 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \pid_alt.source_pid_1_esr_13_LC_8_13_7  (
            .in0(N__23814),
            .in1(N__28047),
            .in2(_gnd_net_),
            .in3(N__23974),
            .lcout(throttle_command_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47384),
            .ce(N__27913),
            .sr(N__27865));
    defparam \pid_alt.error_d_reg_prev_esr_5_LC_8_14_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_5_LC_8_14_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_5_LC_8_14_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_5_LC_8_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25809),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47371),
            .ce(N__33601),
            .sr(N__43821));
    defparam \pid_alt.error_d_reg_prev_esr_RNIL81T2_5_LC_8_14_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIL81T2_5_LC_8_14_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIL81T2_5_LC_8_14_2 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIL81T2_5_LC_8_14_2  (
            .in0(N__22707),
            .in1(N__25782),
            .in2(_gnd_net_),
            .in3(N__29880),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIL81T2Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNICV511_0_6_LC_8_14_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNICV511_0_6_LC_8_14_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNICV511_0_6_LC_8_14_3 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNICV511_0_6_LC_8_14_3  (
            .in0(N__24539),
            .in1(N__24510),
            .in2(_gnd_net_),
            .in3(N__24487),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNICV511_0Z0Z_6 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNICV511_0Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI171A6_5_LC_8_14_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI171A6_5_LC_8_14_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI171A6_5_LC_8_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI171A6_5_LC_8_14_4  (
            .in0(N__22691),
            .in1(N__25781),
            .in2(N__22701),
            .in3(N__29879),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI171A6Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNICUVC3_4_LC_8_14_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNICUVC3_4_LC_8_14_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNICUVC3_4_LC_8_14_5 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNICUVC3_4_LC_8_14_5  (
            .in0(N__24072),
            .in1(N__22677),
            .in2(_gnd_net_),
            .in3(N__29906),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNICUVC3Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI9S511_0_5_LC_8_14_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI9S511_0_5_LC_8_14_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI9S511_0_5_LC_8_14_6 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI9S511_0_5_LC_8_14_6  (
            .in0(N__25848),
            .in1(N__25824),
            .in2(_gnd_net_),
            .in3(N__25808),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI9S511_0Z0Z_5 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNI9S511_0Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIOGSO6_4_LC_8_14_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIOGSO6_4_LC_8_14_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIOGSO6_4_LC_8_14_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIOGSO6_4_LC_8_14_7  (
            .in0(N__24071),
            .in1(N__26048),
            .in2(N__22671),
            .in3(N__29905),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIOGSO6Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIL8611_9_LC_8_15_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIL8611_9_LC_8_15_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIL8611_9_LC_8_15_1 .LUT_INIT=16'b1010111100001010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIL8611_9_LC_8_15_1  (
            .in0(N__22853),
            .in1(_gnd_net_),
            .in2(N__22866),
            .in3(N__22887),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIL8611Z0Z_9 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNIL8611Z0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNICI045_9_LC_8_15_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNICI045_9_LC_8_15_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNICI045_9_LC_8_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNICI045_9_LC_8_15_2  (
            .in0(N__22901),
            .in1(N__23093),
            .in2(N__22983),
            .in3(N__30339),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNICI045Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIDAHM_0_10_LC_8_15_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIDAHM_0_10_LC_8_15_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIDAHM_0_10_LC_8_15_3 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIDAHM_0_10_LC_8_15_3  (
            .in0(N__22970),
            .in1(N__22950),
            .in2(_gnd_net_),
            .in3(N__22932),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIDAHM_0Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_9_LC_8_15_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_9_LC_8_15_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_9_LC_8_15_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_9_LC_8_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22854),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47358),
            .ce(N__33604),
            .sr(N__43827));
    defparam \pid_alt.error_d_reg_prev_esr_RNIG75T2_8_LC_8_15_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIG75T2_8_LC_8_15_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIG75T2_8_LC_8_15_5 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIG75T2_8_LC_8_15_5  (
            .in0(N__22824),
            .in1(N__22830),
            .in2(_gnd_net_),
            .in3(N__30378),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIG75T2Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIL8611_0_9_LC_8_15_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIL8611_0_9_LC_8_15_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIL8611_0_9_LC_8_15_6 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIL8611_0_9_LC_8_15_6  (
            .in0(N__22886),
            .in1(N__22862),
            .in2(_gnd_net_),
            .in3(N__22852),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIL8611_0Z0Z_9 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNIL8611_0Z0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIN49Q5_8_LC_8_15_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIN49Q5_8_LC_8_15_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIN49Q5_8_LC_8_15_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIN49Q5_8_LC_8_15_7  (
            .in0(N__22823),
            .in1(N__22809),
            .in2(N__22782),
            .in3(N__30377),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIN49Q5Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIJR3Q5_6_LC_8_16_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIJR3Q5_6_LC_8_16_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIJR3Q5_6_LC_8_16_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIJR3Q5_6_LC_8_16_0  (
            .in0(N__26345),
            .in1(N__26327),
            .in2(N__22773),
            .in3(N__30480),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIJR3Q5Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIS5212_19_LC_8_16_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIS5212_19_LC_8_16_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIS5212_19_LC_8_16_1 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIS5212_19_LC_8_16_1  (
            .in0(N__23202),
            .in1(N__23184),
            .in2(_gnd_net_),
            .in3(N__30770),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIS5212Z0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_RNI0AAT1_7_LC_8_16_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNI0AAT1_7_LC_8_16_2 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNI0AAT1_7_LC_8_16_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \dron_frame_decoder_1.state_RNI0AAT1_7_LC_8_16_2  (
            .in0(_gnd_net_),
            .in1(N__23163),
            .in2(_gnd_net_),
            .in3(N__44083),
            .lcout(\dron_frame_decoder_1.N_384_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNISSKM_0_26_LC_8_16_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNISSKM_0_26_LC_8_16_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNISSKM_0_26_LC_8_16_4 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNISSKM_0_26_LC_8_16_4  (
            .in0(N__23154),
            .in1(N__23132),
            .in2(_gnd_net_),
            .in3(N__24663),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNISSKM_0Z0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNISAR62_9_LC_8_16_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNISAR62_9_LC_8_16_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNISAR62_9_LC_8_16_7 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNISAR62_9_LC_8_16_7  (
            .in0(N__23100),
            .in1(N__23094),
            .in2(_gnd_net_),
            .in3(N__30338),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNISAR62Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_21_LC_8_17_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_21_LC_8_17_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_21_LC_8_17_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_21_LC_8_17_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23322),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47330),
            .ce(N__33613),
            .sr(N__43843));
    defparam \pid_alt.error_d_reg_prev_esr_RNI27U12_21_LC_8_17_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI27U12_21_LC_8_17_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI27U12_21_LC_8_17_2 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI27U12_21_LC_8_17_2  (
            .in0(N__30697),
            .in1(N__23034),
            .in2(_gnd_net_),
            .in3(N__23028),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI27U12Z0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIIIKM_21_LC_8_17_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIIIKM_21_LC_8_17_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIIIKM_21_LC_8_17_3 .LUT_INIT=16'b1010111100001010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIIIKM_21_LC_8_17_3  (
            .in0(N__23321),
            .in1(_gnd_net_),
            .in2(N__23334),
            .in3(N__24658),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIIIKMZ0Z_21 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNIIIKMZ0Z_21_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI0AS34_21_LC_8_17_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI0AS34_21_LC_8_17_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI0AS34_21_LC_8_17_4 .LUT_INIT=16'b1001011010010110;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI0AS34_21_LC_8_17_4  (
            .in0(N__30696),
            .in1(N__23027),
            .in2(N__23013),
            .in3(N__22997),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI0AS34Z0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIU2U12_20_LC_8_17_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIU2U12_20_LC_8_17_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIU2U12_20_LC_8_17_5 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIU2U12_20_LC_8_17_5  (
            .in0(N__23298),
            .in1(N__23277),
            .in2(_gnd_net_),
            .in3(N__30695),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIU2U12Z0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIIIKM_0_21_LC_8_17_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIIIKM_0_21_LC_8_17_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIIIKM_0_21_LC_8_17_6 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIIIKM_0_21_LC_8_17_6  (
            .in0(N__24657),
            .in1(N__23330),
            .in2(_gnd_net_),
            .in3(N__23320),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIIIKM_0Z0Z_21 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNIIIKM_0Z0Z_21_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIQ8034_20_LC_8_17_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIQ8034_20_LC_8_17_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIQ8034_20_LC_8_17_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIQ8034_20_LC_8_17_7  (
            .in0(N__23291),
            .in1(N__23276),
            .in2(N__23259),
            .in3(N__30694),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIQ8034Z0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_0_c_inv_LC_8_18_2 .C_ON=1'b0;
    defparam \pid_alt.error_cry_0_c_inv_LC_8_18_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_0_c_inv_LC_8_18_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_alt.error_cry_0_c_inv_LC_8_18_2  (
            .in0(N__23243),
            .in1(N__42886),
            .in2(_gnd_net_),
            .in3(N__24418),
            .lcout(\pid_alt.drone_altitude_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_axb_3_LC_8_18_3 .C_ON=1'b0;
    defparam \pid_alt.error_axb_3_LC_8_18_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_axb_3_LC_8_18_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_alt.error_axb_3_LC_8_18_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24390),
            .lcout(\pid_alt.error_axbZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_6_LC_8_18_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_6_LC_8_18_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_6_LC_8_18_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_6_LC_8_18_5  (
            .in0(N__24495),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47314),
            .ce(N__33617),
            .sr(N__43850));
    defparam \pid_alt.error_i_acumm_prereg_esr_3_LC_8_18_6 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_3_LC_8_18_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_3_LC_8_18_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_3_LC_8_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29989),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47314),
            .ce(N__33617),
            .sr(N__43850));
    defparam \pid_alt.error_i_acumm_prereg_esr_13_LC_8_18_7 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_13_LC_8_18_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_13_LC_8_18_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_13_LC_8_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30219),
            .lcout(\pid_alt.error_i_acumm7lto13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47314),
            .ce(N__33617),
            .sr(N__43850));
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIUHR9_10_LC_8_19_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIUHR9_10_LC_8_19_1 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIUHR9_10_LC_8_19_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_RNIUHR9_10_LC_8_19_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24705),
            .lcout(drone_altitude_i_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIVIR9_11_LC_8_19_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIVIR9_11_LC_8_19_2 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIVIR9_11_LC_8_19_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_RNIVIR9_11_LC_8_19_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26157),
            .lcout(drone_altitude_i_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_axb_1_LC_8_19_3 .C_ON=1'b0;
    defparam \pid_alt.error_axb_1_LC_8_19_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_axb_1_LC_8_19_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_alt.error_axb_1_LC_8_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24402),
            .lcout(\pid_alt.error_axbZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_axb_12_LC_8_19_4 .C_ON=1'b0;
    defparam \pid_alt.error_axb_12_LC_8_19_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_axb_12_LC_8_19_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_alt.error_axb_12_LC_8_19_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25182),
            .lcout(\pid_alt.error_axbZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_axb_13_LC_8_19_5 .C_ON=1'b0;
    defparam \pid_alt.error_axb_13_LC_8_19_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_axb_13_LC_8_19_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_alt.error_axb_13_LC_8_19_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25146),
            .lcout(\pid_alt.error_axbZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_axb_14_LC_8_19_6 .C_ON=1'b0;
    defparam \pid_alt.error_axb_14_LC_8_19_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_axb_14_LC_8_19_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_alt.error_axb_14_LC_8_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25098),
            .lcout(\pid_alt.error_axbZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_axb_2_LC_8_19_7 .C_ON=1'b0;
    defparam \pid_alt.error_axb_2_LC_8_19_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_axb_2_LC_8_19_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_alt.error_axb_2_LC_8_19_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24396),
            .lcout(\pid_alt.error_axbZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_ki_0_LC_8_20_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_ki_0_LC_8_20_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_ki_0_LC_8_20_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_ki_0_LC_8_20_0  (
            .in0(_gnd_net_),
            .in1(N__27662),
            .in2(_gnd_net_),
            .in3(N__46682),
            .lcout(alt_ki_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47295),
            .ce(N__44821),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIMNDC_9_LC_8_20_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIMNDC_9_LC_8_20_7 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIMNDC_9_LC_8_20_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_RNIMNDC_9_LC_8_20_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24972),
            .lcout(drone_altitude_i_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_CH1data_0_LC_8_21_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH1data_0_LC_8_21_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH1data_0_LC_8_21_2 .LUT_INIT=16'b0100111101000000;
    LogicCell40 \Commands_frame_decoder.source_CH1data_0_LC_8_21_2  (
            .in0(N__24102),
            .in1(N__27673),
            .in2(N__31851),
            .in3(N__23363),
            .lcout(alt_command_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47288),
            .ce(),
            .sr(N__43873));
    defparam \pid_alt.error_p_reg_esr_5_LC_8_22_7 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_5_LC_8_22_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_5_LC_8_22_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_5_LC_8_22_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23349),
            .lcout(\pid_alt.error_p_regZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47280),
            .ce(N__46784),
            .sr(N__46598));
    defparam \uart_pc_sync.aux_0__0__0_LC_9_1_6 .C_ON=1'b0;
    defparam \uart_pc_sync.aux_0__0__0_LC_9_1_6 .SEQ_MODE=4'b1000;
    defparam \uart_pc_sync.aux_0__0__0_LC_9_1_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_pc_sync.aux_0__0__0_LC_9_1_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23571),
            .lcout(\uart_pc_sync.aux_0__0_Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47475),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.WDT_0_LC_9_5_0 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_0_LC_9_5_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_0_LC_9_5_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_0_LC_9_5_0  (
            .in0(_gnd_net_),
            .in1(N__23547),
            .in2(N__23564),
            .in3(N__23565),
            .lcout(\Commands_frame_decoder.WDTZ0Z_0 ),
            .ltout(),
            .carryin(bfn_9_5_0_),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_0 ),
            .clk(N__47458),
            .ce(),
            .sr(N__25439));
    defparam \Commands_frame_decoder.WDT_1_LC_9_5_1 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_1_LC_9_5_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_1_LC_9_5_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_1_LC_9_5_1  (
            .in0(_gnd_net_),
            .in1(N__23541),
            .in2(_gnd_net_),
            .in3(N__23535),
            .lcout(\Commands_frame_decoder.WDTZ0Z_1 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_0 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_1 ),
            .clk(N__47458),
            .ce(),
            .sr(N__25439));
    defparam \Commands_frame_decoder.WDT_2_LC_9_5_2 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_2_LC_9_5_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_2_LC_9_5_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_2_LC_9_5_2  (
            .in0(_gnd_net_),
            .in1(N__23532),
            .in2(_gnd_net_),
            .in3(N__23526),
            .lcout(\Commands_frame_decoder.WDTZ0Z_2 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_1 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_2 ),
            .clk(N__47458),
            .ce(),
            .sr(N__25439));
    defparam \Commands_frame_decoder.WDT_3_LC_9_5_3 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_3_LC_9_5_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_3_LC_9_5_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_3_LC_9_5_3  (
            .in0(_gnd_net_),
            .in1(N__23523),
            .in2(_gnd_net_),
            .in3(N__23517),
            .lcout(\Commands_frame_decoder.WDTZ0Z_3 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_2 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_3 ),
            .clk(N__47458),
            .ce(),
            .sr(N__25439));
    defparam \Commands_frame_decoder.WDT_4_LC_9_5_4 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_4_LC_9_5_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_4_LC_9_5_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_4_LC_9_5_4  (
            .in0(_gnd_net_),
            .in1(N__23514),
            .in2(_gnd_net_),
            .in3(N__23499),
            .lcout(\Commands_frame_decoder.WDTZ0Z_4 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_3 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_4 ),
            .clk(N__47458),
            .ce(),
            .sr(N__25439));
    defparam \Commands_frame_decoder.WDT_5_LC_9_5_5 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_5_LC_9_5_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_5_LC_9_5_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_5_LC_9_5_5  (
            .in0(_gnd_net_),
            .in1(N__23496),
            .in2(_gnd_net_),
            .in3(N__23481),
            .lcout(\Commands_frame_decoder.WDTZ0Z_5 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_4 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_5 ),
            .clk(N__47458),
            .ce(),
            .sr(N__25439));
    defparam \Commands_frame_decoder.WDT_6_LC_9_5_6 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_6_LC_9_5_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_6_LC_9_5_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_6_LC_9_5_6  (
            .in0(_gnd_net_),
            .in1(N__23478),
            .in2(_gnd_net_),
            .in3(N__23460),
            .lcout(\Commands_frame_decoder.WDTZ0Z_6 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_5 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_6 ),
            .clk(N__47458),
            .ce(),
            .sr(N__25439));
    defparam \Commands_frame_decoder.WDT_7_LC_9_5_7 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_7_LC_9_5_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_7_LC_9_5_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_7_LC_9_5_7  (
            .in0(_gnd_net_),
            .in1(N__23457),
            .in2(_gnd_net_),
            .in3(N__23439),
            .lcout(\Commands_frame_decoder.WDTZ0Z_7 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_6 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_7 ),
            .clk(N__47458),
            .ce(),
            .sr(N__25439));
    defparam \Commands_frame_decoder.WDT_8_LC_9_6_0 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_8_LC_9_6_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_8_LC_9_6_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_8_LC_9_6_0  (
            .in0(_gnd_net_),
            .in1(N__23649),
            .in2(_gnd_net_),
            .in3(N__23634),
            .lcout(\Commands_frame_decoder.WDTZ0Z_8 ),
            .ltout(),
            .carryin(bfn_9_6_0_),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_8 ),
            .clk(N__47449),
            .ce(),
            .sr(N__25440));
    defparam \Commands_frame_decoder.WDT_9_LC_9_6_1 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_9_LC_9_6_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_9_LC_9_6_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_9_LC_9_6_1  (
            .in0(_gnd_net_),
            .in1(N__23629),
            .in2(_gnd_net_),
            .in3(N__23610),
            .lcout(\Commands_frame_decoder.WDTZ0Z_9 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_8 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_9 ),
            .clk(N__47449),
            .ce(),
            .sr(N__25440));
    defparam \Commands_frame_decoder.WDT_10_LC_9_6_2 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_10_LC_9_6_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_10_LC_9_6_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_10_LC_9_6_2  (
            .in0(_gnd_net_),
            .in1(N__23606),
            .in2(_gnd_net_),
            .in3(N__23589),
            .lcout(\Commands_frame_decoder.WDTZ0Z_10 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_9 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_10 ),
            .clk(N__47449),
            .ce(),
            .sr(N__25440));
    defparam \Commands_frame_decoder.WDT_11_LC_9_6_3 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_11_LC_9_6_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_11_LC_9_6_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_11_LC_9_6_3  (
            .in0(_gnd_net_),
            .in1(N__25383),
            .in2(_gnd_net_),
            .in3(N__23586),
            .lcout(\Commands_frame_decoder.WDTZ0Z_11 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_10 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_11 ),
            .clk(N__47449),
            .ce(),
            .sr(N__25440));
    defparam \Commands_frame_decoder.WDT_12_LC_9_6_4 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_12_LC_9_6_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_12_LC_9_6_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_12_LC_9_6_4  (
            .in0(_gnd_net_),
            .in1(N__25407),
            .in2(_gnd_net_),
            .in3(N__23583),
            .lcout(\Commands_frame_decoder.WDTZ0Z_12 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_11 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_12 ),
            .clk(N__47449),
            .ce(),
            .sr(N__25440));
    defparam \Commands_frame_decoder.WDT_13_LC_9_6_5 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_13_LC_9_6_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_13_LC_9_6_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_13_LC_9_6_5  (
            .in0(_gnd_net_),
            .in1(N__25428),
            .in2(_gnd_net_),
            .in3(N__23580),
            .lcout(\Commands_frame_decoder.WDTZ0Z_13 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_12 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_13 ),
            .clk(N__47449),
            .ce(),
            .sr(N__25440));
    defparam \Commands_frame_decoder.WDT_14_LC_9_6_6 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_14_LC_9_6_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_14_LC_9_6_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_14_LC_9_6_6  (
            .in0(_gnd_net_),
            .in1(N__25315),
            .in2(_gnd_net_),
            .in3(N__23577),
            .lcout(\Commands_frame_decoder.WDTZ0Z_14 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_13 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_14 ),
            .clk(N__47449),
            .ce(),
            .sr(N__25440));
    defparam \Commands_frame_decoder.WDT_15_LC_9_6_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.WDT_15_LC_9_6_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_15_LC_9_6_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \Commands_frame_decoder.WDT_15_LC_9_6_7  (
            .in0(_gnd_net_),
            .in1(N__25354),
            .in2(_gnd_net_),
            .in3(N__23574),
            .lcout(\Commands_frame_decoder.WDTZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47449),
            .ce(),
            .sr(N__25440));
    defparam \Commands_frame_decoder.state_RNI4OPK_1_LC_9_7_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNI4OPK_1_LC_9_7_1 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNI4OPK_1_LC_9_7_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \Commands_frame_decoder.state_RNI4OPK_1_LC_9_7_1  (
            .in0(_gnd_net_),
            .in1(N__26476),
            .in2(_gnd_net_),
            .in3(N__25581),
            .lcout(\Commands_frame_decoder.N_320_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_ns_i_a2_2_0_LC_9_7_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_ns_i_a2_2_0_LC_9_7_4 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_ns_i_a2_2_0_LC_9_7_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Commands_frame_decoder.state_ns_i_a2_2_0_LC_9_7_4  (
            .in0(N__27041),
            .in1(N__43286),
            .in2(N__33404),
            .in3(N__25599),
            .lcout(\Commands_frame_decoder.N_364 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_0_LC_9_8_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_0_LC_9_8_0 .SEQ_MODE=4'b1001;
    defparam \Commands_frame_decoder.state_0_LC_9_8_0 .LUT_INIT=16'b0000000010110000;
    LogicCell40 \Commands_frame_decoder.state_0_LC_9_8_0  (
            .in0(N__25617),
            .in1(N__24861),
            .in2(N__25539),
            .in3(N__23727),
            .lcout(\Commands_frame_decoder.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47432),
            .ce(),
            .sr(N__43802));
    defparam \Commands_frame_decoder.state_1_LC_9_8_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_1_LC_9_8_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_1_LC_9_8_2 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \Commands_frame_decoder.state_1_LC_9_8_2  (
            .in0(N__25562),
            .in1(N__25584),
            .in2(N__25227),
            .in3(N__24859),
            .lcout(\Commands_frame_decoder.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47432),
            .ce(),
            .sr(N__43802));
    defparam \Commands_frame_decoder.state_2_LC_9_8_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_2_LC_9_8_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_2_LC_9_8_4 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \Commands_frame_decoder.state_2_LC_9_8_4  (
            .in0(N__25563),
            .in1(N__25590),
            .in2(N__23721),
            .in3(N__24860),
            .lcout(\Commands_frame_decoder.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47432),
            .ce(),
            .sr(N__43802));
    defparam \Commands_frame_decoder.state_RNIEI1J_2_LC_9_8_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIEI1J_2_LC_9_8_7 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIEI1J_2_LC_9_8_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Commands_frame_decoder.state_RNIEI1J_2_LC_9_8_7  (
            .in0(_gnd_net_),
            .in1(N__23717),
            .in2(_gnd_net_),
            .in3(N__26972),
            .lcout(\Commands_frame_decoder.un1_sink_data_valid_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_11_LC_9_9_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_11_LC_9_9_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_11_LC_9_9_0 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \Commands_frame_decoder.state_11_LC_9_9_0  (
            .in0(N__23701),
            .in1(N__26989),
            .in2(N__23778),
            .in3(N__24853),
            .lcout(\Commands_frame_decoder.stateZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47423),
            .ce(),
            .sr(N__43806));
    defparam \Commands_frame_decoder.state_7_LC_9_9_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_7_LC_9_9_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_7_LC_9_9_1 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \Commands_frame_decoder.state_7_LC_9_9_1  (
            .in0(N__24858),
            .in1(N__25528),
            .in2(N__23682),
            .in3(N__26998),
            .lcout(\Commands_frame_decoder.stateZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47423),
            .ce(),
            .sr(N__43806));
    defparam \Commands_frame_decoder.state_6_LC_9_9_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_6_LC_9_9_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_6_LC_9_9_2 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \Commands_frame_decoder.state_6_LC_9_9_2  (
            .in0(N__25529),
            .in1(N__25716),
            .in2(_gnd_net_),
            .in3(N__24857),
            .lcout(\Commands_frame_decoder.stateZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47423),
            .ce(),
            .sr(N__43806));
    defparam \Commands_frame_decoder.WDT_RNIPRJG5_15_LC_9_9_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.WDT_RNIPRJG5_15_LC_9_9_3 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.WDT_RNIPRJG5_15_LC_9_9_3 .LUT_INIT=16'b0000010100000111;
    LogicCell40 \Commands_frame_decoder.WDT_RNIPRJG5_15_LC_9_9_3  (
            .in0(N__25358),
            .in1(N__25317),
            .in2(N__27026),
            .in3(N__23667),
            .lcout(\Commands_frame_decoder.N_358 ),
            .ltout(\Commands_frame_decoder.N_358_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_10_LC_9_9_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_10_LC_9_9_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_10_LC_9_9_4 .LUT_INIT=16'b1111111110100000;
    LogicCell40 \Commands_frame_decoder.state_10_LC_9_9_4  (
            .in0(N__23776),
            .in1(_gnd_net_),
            .in2(N__23781),
            .in3(N__27348),
            .lcout(\Commands_frame_decoder.stateZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47423),
            .ce(),
            .sr(N__43806));
    defparam \Commands_frame_decoder.state_3_LC_9_9_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_3_LC_9_9_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_3_LC_9_9_5 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \Commands_frame_decoder.state_3_LC_9_9_5  (
            .in0(N__24854),
            .in1(N__23753),
            .in2(_gnd_net_),
            .in3(N__31810),
            .lcout(\Commands_frame_decoder.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47423),
            .ce(),
            .sr(N__43806));
    defparam \Commands_frame_decoder.state_4_LC_9_9_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_4_LC_9_9_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_4_LC_9_9_6 .LUT_INIT=16'b1110111010101010;
    LogicCell40 \Commands_frame_decoder.state_4_LC_9_9_6  (
            .in0(N__23739),
            .in1(N__25479),
            .in2(_gnd_net_),
            .in3(N__24855),
            .lcout(\Commands_frame_decoder.stateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47423),
            .ce(),
            .sr(N__43806));
    defparam \Commands_frame_decoder.state_5_LC_9_9_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_5_LC_9_9_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_5_LC_9_9_7 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \Commands_frame_decoder.state_5_LC_9_9_7  (
            .in0(N__24856),
            .in1(N__25467),
            .in2(_gnd_net_),
            .in3(N__25728),
            .lcout(\Commands_frame_decoder.stateZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47423),
            .ce(),
            .sr(N__43806));
    defparam \uart_drone.data_esr_0_LC_9_10_0 .C_ON=1'b0;
    defparam \uart_drone.data_esr_0_LC_9_10_0 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_esr_0_LC_9_10_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone.data_esr_0_LC_9_10_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25703),
            .lcout(uart_drone_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47411),
            .ce(N__26601),
            .sr(N__26619));
    defparam \uart_drone.data_esr_1_LC_9_10_1 .C_ON=1'b0;
    defparam \uart_drone.data_esr_1_LC_9_10_1 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_esr_1_LC_9_10_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone.data_esr_1_LC_9_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25688),
            .lcout(uart_drone_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47411),
            .ce(N__26601),
            .sr(N__26619));
    defparam \uart_drone.data_esr_2_LC_9_10_2 .C_ON=1'b0;
    defparam \uart_drone.data_esr_2_LC_9_10_2 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_esr_2_LC_9_10_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone.data_esr_2_LC_9_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25673),
            .lcout(uart_drone_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47411),
            .ce(N__26601),
            .sr(N__26619));
    defparam \uart_drone.data_esr_3_LC_9_10_3 .C_ON=1'b0;
    defparam \uart_drone.data_esr_3_LC_9_10_3 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_esr_3_LC_9_10_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uart_drone.data_esr_3_LC_9_10_3  (
            .in0(N__25658),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(uart_drone_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47411),
            .ce(N__26601),
            .sr(N__26619));
    defparam \uart_drone.data_esr_4_LC_9_10_4 .C_ON=1'b0;
    defparam \uart_drone.data_esr_4_LC_9_10_4 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_esr_4_LC_9_10_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone.data_esr_4_LC_9_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25644),
            .lcout(uart_drone_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47411),
            .ce(N__26601),
            .sr(N__26619));
    defparam \uart_drone.data_esr_5_LC_9_10_5 .C_ON=1'b0;
    defparam \uart_drone.data_esr_5_LC_9_10_5 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_esr_5_LC_9_10_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uart_drone.data_esr_5_LC_9_10_5  (
            .in0(N__25631),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(uart_drone_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47411),
            .ce(N__26601),
            .sr(N__26619));
    defparam \uart_drone.data_esr_6_LC_9_10_6 .C_ON=1'b0;
    defparam \uart_drone.data_esr_6_LC_9_10_6 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_esr_6_LC_9_10_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone.data_esr_6_LC_9_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25769),
            .lcout(uart_drone_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47411),
            .ce(N__26601),
            .sr(N__26619));
    defparam \uart_drone.data_esr_7_LC_9_10_7 .C_ON=1'b0;
    defparam \uart_drone.data_esr_7_LC_9_10_7 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_esr_7_LC_9_10_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone.data_esr_7_LC_9_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25754),
            .lcout(uart_drone_data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47411),
            .ce(N__26601),
            .sr(N__26619));
    defparam \Commands_frame_decoder.source_offset3data_ess_7_LC_9_11_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset3data_ess_7_LC_9_11_7 .SEQ_MODE=4'b1001;
    defparam \Commands_frame_decoder.source_offset3data_ess_7_LC_9_11_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset3data_ess_7_LC_9_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44984),
            .lcout(frame_decoder_OFF3data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47399),
            .ce(N__26744),
            .sr(N__43812));
    defparam \pid_alt.pid_prereg_esr_RNIU1UR2_14_LC_9_12_0 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNIU1UR2_14_LC_9_12_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNIU1UR2_14_LC_9_12_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \pid_alt.pid_prereg_esr_RNIU1UR2_14_LC_9_12_0  (
            .in0(N__23990),
            .in1(N__23892),
            .in2(N__23877),
            .in3(N__23864),
            .lcout(\pid_alt.N_123 ),
            .ltout(\pid_alt.N_123_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNI0T1S7_0_LC_9_12_1 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNI0T1S7_0_LC_9_12_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNI0T1S7_0_LC_9_12_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \pid_alt.pid_prereg_esr_RNI0T1S7_0_LC_9_12_1  (
            .in0(N__23850),
            .in1(N__24144),
            .in2(N__23841),
            .in3(N__23942),
            .lcout(\pid_alt.N_100 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNIH58S_8_LC_9_12_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIH58S_8_LC_9_12_2 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIH58S_8_LC_9_12_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \Commands_frame_decoder.state_RNIH58S_8_LC_9_12_2  (
            .in0(_gnd_net_),
            .in1(N__24881),
            .in2(_gnd_net_),
            .in3(N__44085),
            .lcout(\Commands_frame_decoder.source_offset3data_1_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNIV9C73_12_LC_9_12_3 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNIV9C73_12_LC_9_12_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNIV9C73_12_LC_9_12_3 .LUT_INIT=16'b0111011100000000;
    LogicCell40 \pid_alt.pid_prereg_esr_RNIV9C73_12_LC_9_12_3  (
            .in0(N__23979),
            .in1(N__23838),
            .in2(_gnd_net_),
            .in3(N__23812),
            .lcout(\pid_alt.N_106 ),
            .ltout(\pid_alt.N_106_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNIIJ486_30_LC_9_12_4 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNIIJ486_30_LC_9_12_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNIIJ486_30_LC_9_12_4 .LUT_INIT=16'b0010001100000011;
    LogicCell40 \pid_alt.pid_prereg_esr_RNIIJ486_30_LC_9_12_4  (
            .in0(N__23943),
            .in1(N__28068),
            .in2(N__23799),
            .in3(N__24207),
            .lcout(\pid_alt.N_91_1 ),
            .ltout(\pid_alt.N_91_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un9lto29_i_a2_7_c_RNI7EJCF_LC_9_12_5 .C_ON=1'b0;
    defparam \pid_alt.un9lto29_i_a2_7_c_RNI7EJCF_LC_9_12_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un9lto29_i_a2_7_c_RNI7EJCF_LC_9_12_5 .LUT_INIT=16'b1111111111001110;
    LogicCell40 \pid_alt.un9lto29_i_a2_7_c_RNI7EJCF_LC_9_12_5  (
            .in0(N__23796),
            .in1(N__23790),
            .in2(N__23784),
            .in3(N__32928),
            .lcout(\pid_alt.un1_reset_0_i ),
            .ltout(\pid_alt.un1_reset_0_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.state_RNIS3RQF_1_LC_9_12_6 .C_ON=1'b0;
    defparam \pid_alt.state_RNIS3RQF_1_LC_9_12_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.state_RNIS3RQF_1_LC_9_12_6 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \pid_alt.state_RNIS3RQF_1_LC_9_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__24048),
            .in3(N__33181),
            .lcout(\pid_alt.N_96_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNII41N_24_LC_9_13_0 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNII41N_24_LC_9_13_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNII41N_24_LC_9_13_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_alt.pid_prereg_esr_RNII41N_24_LC_9_13_0  (
            .in0(N__24045),
            .in1(N__24033),
            .in2(N__24021),
            .in3(N__24006),
            .lcout(\pid_alt.un9lto29_i_a2_5_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.source_pid_1_esr_5_LC_9_13_2 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_esr_5_LC_9_13_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_esr_5_LC_9_13_2 .LUT_INIT=16'b1111000000100000;
    LogicCell40 \pid_alt.source_pid_1_esr_5_LC_9_13_2  (
            .in0(N__27977),
            .in1(N__23941),
            .in2(N__24198),
            .in3(N__28065),
            .lcout(throttle_command_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47372),
            .ce(N__27912),
            .sr(N__27863));
    defparam \pid_alt.source_pid_1_esr_10_LC_9_13_3 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_esr_10_LC_9_13_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_esr_10_LC_9_13_3 .LUT_INIT=16'b1010101010101111;
    LogicCell40 \pid_alt.source_pid_1_esr_10_LC_9_13_3  (
            .in0(N__27105),
            .in1(_gnd_net_),
            .in2(N__28072),
            .in3(N__27975),
            .lcout(throttle_command_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47372),
            .ce(N__27912),
            .sr(N__27863));
    defparam \pid_alt.source_pid_1_esr_11_LC_9_13_4 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_esr_11_LC_9_13_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_esr_11_LC_9_13_4 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \pid_alt.source_pid_1_esr_11_LC_9_13_4  (
            .in0(N__27976),
            .in1(N__28057),
            .in2(_gnd_net_),
            .in3(N__27140),
            .lcout(throttle_command_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47372),
            .ce(N__27912),
            .sr(N__27863));
    defparam \pid_alt.source_pid_1_esr_7_LC_9_13_6 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_esr_7_LC_9_13_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_esr_7_LC_9_13_6 .LUT_INIT=16'b1111000011110101;
    LogicCell40 \pid_alt.source_pid_1_esr_7_LC_9_13_6  (
            .in0(N__27978),
            .in1(_gnd_net_),
            .in2(N__27177),
            .in3(N__28058),
            .lcout(throttle_command_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47372),
            .ce(N__27912),
            .sr(N__27863));
    defparam \pid_alt.source_pid_1_esr_8_LC_9_13_7 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_esr_8_LC_9_13_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_esr_8_LC_9_13_7 .LUT_INIT=16'b1010101010101111;
    LogicCell40 \pid_alt.source_pid_1_esr_8_LC_9_13_7  (
            .in0(N__23925),
            .in1(_gnd_net_),
            .in2(N__28073),
            .in3(N__27979),
            .lcout(throttle_command_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47372),
            .ce(N__27912),
            .sr(N__27863));
    defparam \pid_alt.pid_prereg_esr_RNI0VB22_6_LC_9_14_0 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNI0VB22_6_LC_9_14_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNI0VB22_6_LC_9_14_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \pid_alt.pid_prereg_esr_RNI0VB22_6_LC_9_14_0  (
            .in0(N__26006),
            .in1(N__23975),
            .in2(N__27078),
            .in3(N__23921),
            .lcout(\pid_alt.N_124 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un9lto29_i_a2_2_c_RNO_LC_9_14_2 .C_ON=1'b0;
    defparam \pid_alt.un9lto29_i_a2_2_c_RNO_LC_9_14_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un9lto29_i_a2_2_c_RNO_LC_9_14_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_alt.un9lto29_i_a2_2_c_RNO_LC_9_14_2  (
            .in0(N__27940),
            .in1(N__27097),
            .in2(N__27136),
            .in3(N__23920),
            .lcout(\pid_alt.N_12_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un9lto29_i_a2_1_c_RNO_LC_9_14_3 .C_ON=1'b0;
    defparam \pid_alt.un9lto29_i_a2_1_c_RNO_LC_9_14_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un9lto29_i_a2_1_c_RNO_LC_9_14_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_alt.un9lto29_i_a2_1_c_RNO_LC_9_14_3  (
            .in0(N__24195),
            .in1(N__26005),
            .in2(N__27170),
            .in3(N__24166),
            .lcout(\pid_alt.un9lto29_i_a2_0_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNI35JO_4_LC_9_14_4 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNI35JO_4_LC_9_14_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNI35JO_4_LC_9_14_4 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \pid_alt.pid_prereg_esr_RNI35JO_4_LC_9_14_4  (
            .in0(N__24168),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24197),
            .lcout(\pid_alt.N_96 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNIL84J1_0_LC_9_14_5 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNIL84J1_0_LC_9_14_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNIL84J1_0_LC_9_14_5 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \pid_alt.pid_prereg_esr_RNIL84J1_0_LC_9_14_5  (
            .in0(N__24196),
            .in1(N__24167),
            .in2(N__33172),
            .in3(N__25986),
            .lcout(\pid_alt.source_pid_1_sqmuxa_0_a2_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.state_1_LC_9_14_6 .C_ON=1'b0;
    defparam \pid_alt.state_1_LC_9_14_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.state_1_LC_9_14_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.state_1_LC_9_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24957),
            .lcout(\pid_alt.N_96_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47359),
            .ce(),
            .sr(N__43828));
    defparam \pid_alt.state_RNIFCSD1_0_LC_9_14_7 .C_ON=1'b0;
    defparam \pid_alt.state_RNIFCSD1_0_LC_9_14_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.state_RNIFCSD1_0_LC_9_14_7 .LUT_INIT=16'b1111111100000100;
    LogicCell40 \pid_alt.state_RNIFCSD1_0_LC_9_14_7  (
            .in0(N__33146),
            .in1(N__29590),
            .in2(N__24962),
            .in3(N__44066),
            .lcout(\pid_alt.state_RNIFCSD1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_CH1data8lto7_LC_9_15_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH1data8lto7_LC_9_15_1 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.source_CH1data8lto7_LC_9_15_1 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \Commands_frame_decoder.source_CH1data8lto7_LC_9_15_1  (
            .in0(N__26361),
            .in1(N__25862),
            .in2(N__45351),
            .in3(N__33405),
            .lcout(\Commands_frame_decoder.source_CH1data8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI6P511_4_LC_9_15_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI6P511_4_LC_9_15_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI6P511_4_LC_9_15_3 .LUT_INIT=16'b1010111100001010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI6P511_4_LC_9_15_3  (
            .in0(N__45494),
            .in1(_gnd_net_),
            .in2(N__26022),
            .in3(N__24063),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI6P511Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI6P511_0_4_LC_9_15_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI6P511_0_4_LC_9_15_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI6P511_0_4_LC_9_15_4 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI6P511_0_4_LC_9_15_4  (
            .in0(N__24062),
            .in1(N__26018),
            .in2(_gnd_net_),
            .in3(N__45493),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI6P511_0Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIQQKM_25_LC_9_15_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIQQKM_25_LC_9_15_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIQQKM_25_LC_9_15_7 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIQQKM_25_LC_9_15_7  (
            .in0(N__24300),
            .in1(N__24312),
            .in2(_gnd_net_),
            .in3(N__24662),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIQQKMZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI0BT34_25_LC_9_16_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI0BT34_25_LC_9_16_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI0BT34_25_LC_9_16_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI0BT34_25_LC_9_16_0  (
            .in0(N__30699),
            .in1(N__24359),
            .in2(N__24261),
            .in3(N__24368),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI0BT34Z0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIINU12_25_LC_9_16_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIINU12_25_LC_9_16_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIINU12_25_LC_9_16_2 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIINU12_25_LC_9_16_2  (
            .in0(N__30702),
            .in1(N__24369),
            .in2(_gnd_net_),
            .in3(N__24360),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIINU12Z0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_25_LC_9_16_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_25_LC_9_16_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_25_LC_9_16_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_25_LC_9_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24299),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47331),
            .ce(N__33605),
            .sr(N__43844));
    defparam \pid_alt.error_d_reg_prev_esr_RNIO2T34_24_LC_9_16_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIO2T34_24_LC_9_16_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIO2T34_24_LC_9_16_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIO2T34_24_LC_9_16_5  (
            .in0(N__24548),
            .in1(N__24270),
            .in2(N__24240),
            .in3(N__30701),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIO2T34Z0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIQQKM_0_25_LC_9_16_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIQQKM_0_25_LC_9_16_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIQQKM_0_25_LC_9_16_6 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIQQKM_0_25_LC_9_16_6  (
            .in0(N__24311),
            .in1(N__24298),
            .in2(_gnd_net_),
            .in3(N__24661),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIQQKM_0Z0Z_25 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNIQQKM_0Z0Z_25_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIEJU12_24_LC_9_16_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIEJU12_24_LC_9_16_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIEJU12_24_LC_9_16_7 .LUT_INIT=16'b1111101010100000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIEJU12_24_LC_9_16_7  (
            .in0(N__24549),
            .in1(_gnd_net_),
            .in2(N__24264),
            .in3(N__30700),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIEJU12Z0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_24_LC_9_17_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_24_LC_9_17_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_24_LC_9_17_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_24_LC_9_17_0  (
            .in0(N__24690),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47315),
            .ce(N__33608),
            .sr(N__43851));
    defparam \pid_alt.error_d_reg_prev_esr_RNIOOKM_0_24_LC_9_17_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIOOKM_0_24_LC_9_17_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIOOKM_0_24_LC_9_17_1 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIOOKM_0_24_LC_9_17_1  (
            .in0(N__24698),
            .in1(N__24688),
            .in2(_gnd_net_),
            .in3(N__24659),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIOOKM_0Z0Z_24 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNIOOKM_0Z0Z_24_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIAFU12_23_LC_9_17_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIAFU12_23_LC_9_17_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIAFU12_23_LC_9_17_2 .LUT_INIT=16'b1111110011000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIAFU12_23_LC_9_17_2  (
            .in0(_gnd_net_),
            .in1(N__26280),
            .in2(N__24243),
            .in3(N__30698),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIAFU12Z0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIOOKM_24_LC_9_17_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIOOKM_24_LC_9_17_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIOOKM_24_LC_9_17_3 .LUT_INIT=16'b1101110101000100;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIOOKM_24_LC_9_17_3  (
            .in0(N__24699),
            .in1(N__24689),
            .in2(_gnd_net_),
            .in3(N__24660),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIOOKMZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNICV511_6_LC_9_17_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNICV511_6_LC_9_17_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNICV511_6_LC_9_17_7 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNICV511_6_LC_9_17_7  (
            .in0(N__24540),
            .in1(N__24509),
            .in2(_gnd_net_),
            .in3(N__24494),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNICV511Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_0_LC_9_18_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_0_LC_9_18_0 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_0_LC_9_18_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_0_LC_9_18_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25049),
            .lcout(drone_altitude_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47304),
            .ce(N__24900),
            .sr(N__43857));
    defparam \dron_frame_decoder_1.source_Altitude_esr_1_LC_9_18_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_1_LC_9_18_1 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_1_LC_9_18_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_1_LC_9_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25010),
            .lcout(drone_altitude_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47304),
            .ce(N__24900),
            .sr(N__43857));
    defparam \dron_frame_decoder_1.source_Altitude_esr_2_LC_9_18_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_2_LC_9_18_2 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_2_LC_9_18_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_2_LC_9_18_2  (
            .in0(N__24730),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(drone_altitude_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47304),
            .ce(N__24900),
            .sr(N__43857));
    defparam \dron_frame_decoder_1.source_Altitude_esr_3_LC_9_18_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_3_LC_9_18_3 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_3_LC_9_18_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_3_LC_9_18_3  (
            .in0(N__26201),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(drone_altitude_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47304),
            .ce(N__24900),
            .sr(N__43857));
    defparam \dron_frame_decoder_1.source_Altitude_esr_4_LC_9_18_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_4_LC_9_18_4 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_4_LC_9_18_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_4_LC_9_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25217),
            .lcout(\dron_frame_decoder_1.drone_altitude_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47304),
            .ce(N__24900),
            .sr(N__43857));
    defparam \dron_frame_decoder_1.source_Altitude_esr_5_LC_9_18_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_5_LC_9_18_5 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_5_LC_9_18_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_5_LC_9_18_5  (
            .in0(N__25175),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\dron_frame_decoder_1.drone_altitude_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47304),
            .ce(N__24900),
            .sr(N__43857));
    defparam \dron_frame_decoder_1.source_Altitude_esr_6_LC_9_18_6 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_6_LC_9_18_6 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_6_LC_9_18_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_6_LC_9_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25139),
            .lcout(\dron_frame_decoder_1.drone_altitude_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47304),
            .ce(N__24900),
            .sr(N__43857));
    defparam \dron_frame_decoder_1.source_Altitude_esr_7_LC_9_18_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_7_LC_9_18_7 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_7_LC_9_18_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_7_LC_9_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25091),
            .lcout(\dron_frame_decoder_1.drone_altitude_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47304),
            .ce(N__24900),
            .sr(N__43857));
    defparam \Commands_frame_decoder.state_9_LC_9_19_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_9_LC_9_19_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_9_LC_9_19_0 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \Commands_frame_decoder.state_9_LC_9_19_0  (
            .in0(N__27059),
            .in1(N__24888),
            .in2(_gnd_net_),
            .in3(N__24867),
            .lcout(\Commands_frame_decoder.stateZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47296),
            .ce(),
            .sr(N__43865));
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIHIDC_4_LC_9_19_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIHIDC_4_LC_9_19_3 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIHIDC_4_LC_9_19_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_RNIHIDC_4_LC_9_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24816),
            .lcout(drone_altitude_i_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIIJDC_5_LC_9_19_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIIJDC_5_LC_9_19_4 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIIJDC_5_LC_9_19_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_RNIIJDC_5_LC_9_19_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24798),
            .lcout(drone_altitude_i_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIJKDC_6_LC_9_19_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIJKDC_6_LC_9_19_5 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIJKDC_6_LC_9_19_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_RNIJKDC_6_LC_9_19_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24780),
            .lcout(drone_altitude_i_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIKLDC_7_LC_9_19_6 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIKLDC_7_LC_9_19_6 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIKLDC_7_LC_9_19_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_RNIKLDC_7_LC_9_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24765),
            .lcout(drone_altitude_i_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNILMDC_8_LC_9_19_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNILMDC_8_LC_9_19_7 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNILMDC_8_LC_9_19_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_RNILMDC_8_LC_9_19_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__25020),
            .in3(_gnd_net_),
            .lcout(drone_altitude_i_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_10_LC_9_20_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_10_LC_9_20_0 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_10_LC_9_20_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_10_LC_9_20_0  (
            .in0(N__24731),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\dron_frame_decoder_1.drone_altitude_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47289),
            .ce(N__26148),
            .sr(N__43874));
    defparam \dron_frame_decoder_1.source_Altitude_esr_12_LC_9_20_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_12_LC_9_20_2 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_12_LC_9_20_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_12_LC_9_20_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25218),
            .lcout(drone_altitude_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47289),
            .ce(N__26148),
            .sr(N__43874));
    defparam \dron_frame_decoder_1.source_Altitude_esr_13_LC_9_20_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_13_LC_9_20_3 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_13_LC_9_20_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_13_LC_9_20_3  (
            .in0(N__25176),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(drone_altitude_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47289),
            .ce(N__26148),
            .sr(N__43874));
    defparam \dron_frame_decoder_1.source_Altitude_esr_14_LC_9_20_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_14_LC_9_20_4 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_14_LC_9_20_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_14_LC_9_20_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25140),
            .lcout(drone_altitude_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47289),
            .ce(N__26148),
            .sr(N__43874));
    defparam \dron_frame_decoder_1.source_Altitude_esr_15_LC_9_20_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_15_LC_9_20_5 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_15_LC_9_20_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_15_LC_9_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25092),
            .lcout(drone_altitude_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47289),
            .ce(N__26148),
            .sr(N__43874));
    defparam \dron_frame_decoder_1.source_Altitude_esr_8_LC_9_20_6 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_8_LC_9_20_6 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_8_LC_9_20_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_8_LC_9_20_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25053),
            .lcout(\dron_frame_decoder_1.drone_altitude_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47289),
            .ce(N__26148),
            .sr(N__43874));
    defparam \dron_frame_decoder_1.source_Altitude_esr_9_LC_9_20_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_9_LC_9_20_7 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_9_LC_9_20_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_9_LC_9_20_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25011),
            .lcout(\dron_frame_decoder_1.drone_altitude_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47289),
            .ce(N__26148),
            .sr(N__43874));
    defparam \Commands_frame_decoder.source_CH4data_esr_4_LC_9_21_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH4data_esr_4_LC_9_21_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH4data_esr_4_LC_9_21_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH4data_esr_4_LC_9_21_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45358),
            .lcout(frame_decoder_CH4data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47281),
            .ce(N__26396),
            .sr(N__43879));
    defparam \pid_alt.state_RNIH1EN_0_LC_10_3_4 .C_ON=1'b0;
    defparam \pid_alt.state_RNIH1EN_0_LC_10_3_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.state_RNIH1EN_0_LC_10_3_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \pid_alt.state_RNIH1EN_0_LC_10_3_4  (
            .in0(_gnd_net_),
            .in1(N__24966),
            .in2(_gnd_net_),
            .in3(N__44069),
            .lcout(\pid_alt.state_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc_sync.aux_3__0__0_LC_10_4_2 .C_ON=1'b0;
    defparam \uart_pc_sync.aux_3__0__0_LC_10_4_2 .SEQ_MODE=4'b1000;
    defparam \uart_pc_sync.aux_3__0__0_LC_10_4_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_pc_sync.aux_3__0__0_LC_10_4_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25461),
            .lcout(\uart_pc_sync.aux_3__0_Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47450),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc_sync.aux_2__0__0_LC_10_4_6 .C_ON=1'b0;
    defparam \uart_pc_sync.aux_2__0__0_LC_10_4_6 .SEQ_MODE=4'b1000;
    defparam \uart_pc_sync.aux_2__0__0_LC_10_4_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_pc_sync.aux_2__0__0_LC_10_4_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25446),
            .lcout(\uart_pc_sync.aux_2__0_Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47450),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc_sync.aux_1__0__0_LC_10_4_7 .C_ON=1'b0;
    defparam \uart_pc_sync.aux_1__0__0_LC_10_4_7 .SEQ_MODE=4'b1000;
    defparam \uart_pc_sync.aux_1__0__0_LC_10_4_7 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \uart_pc_sync.aux_1__0__0_LC_10_4_7  (
            .in0(_gnd_net_),
            .in1(N__25455),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\uart_pc_sync.aux_1__0_Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47450),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.un1_state53_i_LC_10_5_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.un1_state53_i_LC_10_5_5 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.un1_state53_i_LC_10_5_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \Commands_frame_decoder.un1_state53_i_LC_10_5_5  (
            .in0(_gnd_net_),
            .in1(N__27027),
            .in2(_gnd_net_),
            .in3(N__44099),
            .lcout(\Commands_frame_decoder.un1_state53_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.WDT_RNIRGQ51_11_LC_10_6_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.WDT_RNIRGQ51_11_LC_10_6_2 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.WDT_RNIRGQ51_11_LC_10_6_2 .LUT_INIT=16'b0101010101110111;
    LogicCell40 \Commands_frame_decoder.WDT_RNIRGQ51_11_LC_10_6_2  (
            .in0(N__25425),
            .in1(N__25404),
            .in2(_gnd_net_),
            .in3(N__25380),
            .lcout(),
            .ltout(\Commands_frame_decoder.state_0_sqmuxacf0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.preinit_RNIC9QE2_LC_10_6_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.preinit_RNIC9QE2_LC_10_6_3 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.preinit_RNIC9QE2_LC_10_6_3 .LUT_INIT=16'b0001000101010001;
    LogicCell40 \Commands_frame_decoder.preinit_RNIC9QE2_LC_10_6_3  (
            .in0(N__25266),
            .in1(N__25346),
            .in2(N__25320),
            .in3(N__25307),
            .lcout(\Commands_frame_decoder.state_0_sqmuxacf0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.preinit_LC_10_6_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.preinit_LC_10_6_6 .SEQ_MODE=4'b1001;
    defparam \Commands_frame_decoder.preinit_LC_10_6_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Commands_frame_decoder.preinit_LC_10_6_6  (
            .in0(_gnd_net_),
            .in1(N__27028),
            .in2(_gnd_net_),
            .in3(N__25267),
            .lcout(\Commands_frame_decoder.preinitZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47433),
            .ce(),
            .sr(N__43799));
    defparam \Commands_frame_decoder.source_data_valid_LC_10_6_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_data_valid_LC_10_6_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_data_valid_LC_10_6_7 .LUT_INIT=16'b1111101011001010;
    LogicCell40 \Commands_frame_decoder.source_data_valid_LC_10_6_7  (
            .in0(N__25268),
            .in1(N__25251),
            .in2(N__27043),
            .in3(N__30528),
            .lcout(debug_CH3_20A_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47433),
            .ce(),
            .sr(N__43799));
    defparam \Commands_frame_decoder.source_data_valid_RNO_0_LC_10_7_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_data_valid_RNO_0_LC_10_7_6 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.source_data_valid_RNO_0_LC_10_7_6 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Commands_frame_decoder.source_data_valid_RNO_0_LC_10_7_6  (
            .in0(N__26654),
            .in1(N__26634),
            .in2(_gnd_net_),
            .in3(N__26482),
            .lcout(\Commands_frame_decoder.count_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNO_0_1_LC_10_8_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNO_0_1_LC_10_8_0 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNO_0_1_LC_10_8_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Commands_frame_decoder.state_RNO_0_1_LC_10_8_0  (
            .in0(N__26499),
            .in1(N__25242),
            .in2(N__44271),
            .in3(N__36839),
            .lcout(\Commands_frame_decoder.state_ns_0_a4_0_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNO_3_0_LC_10_8_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNO_3_0_LC_10_8_1 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNO_3_0_LC_10_8_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Commands_frame_decoder.state_RNO_3_0_LC_10_8_1  (
            .in0(N__25615),
            .in1(N__44254),
            .in2(N__36866),
            .in3(N__26498),
            .lcout(\Commands_frame_decoder.N_359 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_ns_i_a2_2_1_0_LC_10_8_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_ns_i_a2_2_1_0_LC_10_8_2 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_ns_i_a2_2_1_0_LC_10_8_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Commands_frame_decoder.state_ns_i_a2_2_1_0_LC_10_8_2  (
            .in0(_gnd_net_),
            .in1(N__45274),
            .in2(_gnd_net_),
            .in3(N__45176),
            .lcout(\Commands_frame_decoder.state_ns_i_a2_2_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNO_1_2_LC_10_8_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNO_1_2_LC_10_8_3 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNO_1_2_LC_10_8_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \Commands_frame_decoder.state_RNO_1_2_LC_10_8_3  (
            .in0(_gnd_net_),
            .in1(N__44954),
            .in2(_gnd_net_),
            .in3(N__27615),
            .lcout(),
            .ltout(\Commands_frame_decoder.state_ns_0_a4_0_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNO_0_2_LC_10_8_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNO_0_2_LC_10_8_4 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNO_0_2_LC_10_8_4 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \Commands_frame_decoder.state_RNO_0_2_LC_10_8_4  (
            .in0(N__44258),
            .in1(N__36838),
            .in2(N__25593),
            .in3(N__25583),
            .lcout(\Commands_frame_decoder.state_ns_0_a4_0_3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNO_4_0_LC_10_8_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNO_4_0_LC_10_8_6 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNO_4_0_LC_10_8_6 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \Commands_frame_decoder.state_RNO_4_0_LC_10_8_6  (
            .in0(N__27616),
            .in1(N__25866),
            .in2(N__36867),
            .in3(N__25582),
            .lcout(),
            .ltout(\Commands_frame_decoder.N_360_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNO_1_0_LC_10_8_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNO_1_0_LC_10_8_7 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNO_1_0_LC_10_8_7 .LUT_INIT=16'b0001000100010101;
    LogicCell40 \Commands_frame_decoder.state_RNO_1_0_LC_10_8_7  (
            .in0(N__26444),
            .in1(N__25561),
            .in2(N__25548),
            .in3(N__25545),
            .lcout(\Commands_frame_decoder.state_ns_i_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kp_4_LC_10_9_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kp_4_LC_10_9_0 .SEQ_MODE=4'b1001;
    defparam \Commands_frame_decoder.source_alt_kp_4_LC_10_9_0 .LUT_INIT=16'b1110101000101010;
    LogicCell40 \Commands_frame_decoder.source_alt_kp_4_LC_10_9_0  (
            .in0(N__25493),
            .in1(N__27022),
            .in2(N__25530),
            .in3(N__45296),
            .lcout(alt_kp_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47401),
            .ce(),
            .sr(N__43807));
    defparam \uart_pc.data_rdy_LC_10_9_1 .C_ON=1'b0;
    defparam \uart_pc.data_rdy_LC_10_9_1 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_rdy_LC_10_9_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uart_pc.data_rdy_LC_10_9_1  (
            .in0(N__26585),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31228),
            .lcout(uart_pc_data_rdy),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47401),
            .ce(),
            .sr(N__43807));
    defparam \Commands_frame_decoder.state_RNIGK1J_4_LC_10_9_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIGK1J_4_LC_10_9_4 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIGK1J_4_LC_10_9_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Commands_frame_decoder.state_RNIGK1J_4_LC_10_9_4  (
            .in0(_gnd_net_),
            .in1(N__25478),
            .in2(_gnd_net_),
            .in3(N__27020),
            .lcout(\Commands_frame_decoder.source_CH3data_1_sqmuxa ),
            .ltout(\Commands_frame_decoder.source_CH3data_1_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNID18S_4_LC_10_9_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNID18S_4_LC_10_9_5 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNID18S_4_LC_10_9_5 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \Commands_frame_decoder.state_RNID18S_4_LC_10_9_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__25731),
            .in3(N__44073),
            .lcout(\Commands_frame_decoder.source_CH3data_1_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNIHL1J_5_LC_10_9_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIHL1J_5_LC_10_9_6 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIHL1J_5_LC_10_9_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Commands_frame_decoder.state_RNIHL1J_5_LC_10_9_6  (
            .in0(_gnd_net_),
            .in1(N__25727),
            .in2(_gnd_net_),
            .in3(N__27021),
            .lcout(\Commands_frame_decoder.source_CH4data_1_sqmuxa ),
            .ltout(\Commands_frame_decoder.source_CH4data_1_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNIE28S_5_LC_10_9_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIE28S_5_LC_10_9_7 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIE28S_5_LC_10_9_7 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \Commands_frame_decoder.state_RNIE28S_5_LC_10_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__25707),
            .in3(N__44072),
            .lcout(\Commands_frame_decoder.source_CH4data_1_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.data_Aux_0_LC_10_10_0 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_0_LC_10_10_0 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_Aux_0_LC_10_10_0 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \uart_drone.data_Aux_0_LC_10_10_0  (
            .in0(N__26556),
            .in1(N__31382),
            .in2(N__25704),
            .in3(N__31430),
            .lcout(\uart_drone.data_AuxZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47386),
            .ce(),
            .sr(N__31869));
    defparam \uart_drone.data_Aux_1_LC_10_10_1 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_1_LC_10_10_1 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_Aux_1_LC_10_10_1 .LUT_INIT=16'b1111010010110000;
    LogicCell40 \uart_drone.data_Aux_1_LC_10_10_1  (
            .in0(N__31431),
            .in1(N__26550),
            .in2(N__25689),
            .in3(N__31389),
            .lcout(\uart_drone.data_AuxZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47386),
            .ce(),
            .sr(N__31869));
    defparam \uart_drone.data_Aux_2_LC_10_10_2 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_2_LC_10_10_2 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_Aux_2_LC_10_10_2 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \uart_drone.data_Aux_2_LC_10_10_2  (
            .in0(N__34089),
            .in1(N__31383),
            .in2(N__25674),
            .in3(N__31432),
            .lcout(\uart_drone.data_AuxZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47386),
            .ce(),
            .sr(N__31869));
    defparam \uart_drone.data_Aux_3_LC_10_10_3 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_3_LC_10_10_3 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_Aux_3_LC_10_10_3 .LUT_INIT=16'b1111010010110000;
    LogicCell40 \uart_drone.data_Aux_3_LC_10_10_3  (
            .in0(N__31433),
            .in1(N__27507),
            .in2(N__25659),
            .in3(N__31390),
            .lcout(\uart_drone.data_AuxZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47386),
            .ce(),
            .sr(N__31869));
    defparam \uart_drone.data_Aux_4_LC_10_10_4 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_4_LC_10_10_4 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_Aux_4_LC_10_10_4 .LUT_INIT=16'b1100110011100100;
    LogicCell40 \uart_drone.data_Aux_4_LC_10_10_4  (
            .in0(N__27519),
            .in1(N__25643),
            .in2(N__31397),
            .in3(N__31434),
            .lcout(\uart_drone.data_AuxZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47386),
            .ce(),
            .sr(N__31869));
    defparam \uart_drone.data_Aux_5_LC_10_10_5 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_5_LC_10_10_5 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_Aux_5_LC_10_10_5 .LUT_INIT=16'b1111010010110000;
    LogicCell40 \uart_drone.data_Aux_5_LC_10_10_5  (
            .in0(N__31435),
            .in1(N__27693),
            .in2(N__25632),
            .in3(N__31391),
            .lcout(\uart_drone.data_AuxZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47386),
            .ce(),
            .sr(N__31869));
    defparam \uart_drone.data_Aux_6_LC_10_10_6 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_6_LC_10_10_6 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_Aux_6_LC_10_10_6 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \uart_drone.data_Aux_6_LC_10_10_6  (
            .in0(N__34077),
            .in1(N__31384),
            .in2(N__25770),
            .in3(N__31436),
            .lcout(\uart_drone.data_AuxZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47386),
            .ce(),
            .sr(N__31869));
    defparam \uart_drone.data_Aux_7_LC_10_10_7 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_7_LC_10_10_7 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_Aux_7_LC_10_10_7 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \uart_drone.data_Aux_7_LC_10_10_7  (
            .in0(N__31437),
            .in1(N__31388),
            .in2(N__25755),
            .in3(N__44468),
            .lcout(\uart_drone.data_AuxZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47386),
            .ce(),
            .sr(N__31869));
    defparam \Commands_frame_decoder.source_CH3data_esr_0_LC_10_11_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH3data_esr_0_LC_10_11_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH3data_esr_0_LC_10_11_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH3data_esr_0_LC_10_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27652),
            .lcout(frame_decoder_CH3data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47374),
            .ce(N__25740),
            .sr(N__43813));
    defparam \Commands_frame_decoder.source_CH3data_esr_1_LC_10_11_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH3data_esr_1_LC_10_11_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH3data_esr_1_LC_10_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH3data_esr_1_LC_10_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45211),
            .lcout(frame_decoder_CH3data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47374),
            .ce(N__25740),
            .sr(N__43813));
    defparam \Commands_frame_decoder.source_CH3data_esr_2_LC_10_11_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH3data_esr_2_LC_10_11_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH3data_esr_2_LC_10_11_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Commands_frame_decoder.source_CH3data_esr_2_LC_10_11_2  (
            .in0(N__36864),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(frame_decoder_CH3data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47374),
            .ce(N__25740),
            .sr(N__43813));
    defparam \Commands_frame_decoder.source_CH3data_esr_3_LC_10_11_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH3data_esr_3_LC_10_11_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH3data_esr_3_LC_10_11_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH3data_esr_3_LC_10_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43339),
            .lcout(frame_decoder_CH3data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47374),
            .ce(N__25740),
            .sr(N__43813));
    defparam \Commands_frame_decoder.source_CH3data_esr_4_LC_10_11_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH3data_esr_4_LC_10_11_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH3data_esr_4_LC_10_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH3data_esr_4_LC_10_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45314),
            .lcout(frame_decoder_CH3data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47374),
            .ce(N__25740),
            .sr(N__43813));
    defparam \Commands_frame_decoder.source_CH3data_esr_5_LC_10_11_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH3data_esr_5_LC_10_11_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH3data_esr_5_LC_10_11_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH3data_esr_5_LC_10_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44262),
            .lcout(frame_decoder_CH3data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47374),
            .ce(N__25740),
            .sr(N__43813));
    defparam \Commands_frame_decoder.source_CH3data_esr_6_LC_10_11_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH3data_esr_6_LC_10_11_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH3data_esr_6_LC_10_11_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH3data_esr_6_LC_10_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33389),
            .lcout(frame_decoder_CH3data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47374),
            .ce(N__25740),
            .sr(N__43813));
    defparam \Commands_frame_decoder.source_CH3data_ess_7_LC_10_11_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH3data_ess_7_LC_10_11_7 .SEQ_MODE=4'b1001;
    defparam \Commands_frame_decoder.source_CH3data_ess_7_LC_10_11_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH3data_ess_7_LC_10_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44983),
            .lcout(frame_decoder_CH3data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47374),
            .ce(N__25740),
            .sr(N__43813));
    defparam \pid_alt.source_pid_1_esr_6_LC_10_12_7 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_esr_6_LC_10_12_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_esr_6_LC_10_12_7 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \pid_alt.source_pid_1_esr_6_LC_10_12_7  (
            .in0(N__28074),
            .in1(N__27980),
            .in2(_gnd_net_),
            .in3(N__26010),
            .lcout(throttle_command_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47361),
            .ce(N__27917),
            .sr(N__27862));
    defparam \pid_alt.source_pid_1_0_LC_10_13_0 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_0_LC_10_13_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_0_LC_10_13_0 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \pid_alt.source_pid_1_0_LC_10_13_0  (
            .in0(N__33163),
            .in1(N__25904),
            .in2(N__36992),
            .in3(N__25985),
            .lcout(throttle_command_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47346),
            .ce(),
            .sr(N__27864));
    defparam \pid_alt.source_pid_1_1_LC_10_13_1 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_1_LC_10_13_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_1_LC_10_13_1 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \pid_alt.source_pid_1_1_LC_10_13_1  (
            .in0(N__25905),
            .in1(N__33164),
            .in2(N__29300),
            .in3(N__25959),
            .lcout(throttle_command_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47346),
            .ce(),
            .sr(N__27864));
    defparam \pid_alt.source_pid_1_2_LC_10_13_2 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_2_LC_10_13_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_2_LC_10_13_2 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \pid_alt.source_pid_1_2_LC_10_13_2  (
            .in0(N__33165),
            .in1(N__25906),
            .in2(N__29345),
            .in3(N__25932),
            .lcout(throttle_command_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47346),
            .ce(),
            .sr(N__27864));
    defparam \pid_alt.source_pid_1_3_LC_10_13_3 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_3_LC_10_13_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_3_LC_10_13_3 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \pid_alt.source_pid_1_3_LC_10_13_3  (
            .in0(N__25907),
            .in1(N__33166),
            .in2(N__35477),
            .in3(N__25887),
            .lcout(throttle_command_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47346),
            .ce(),
            .sr(N__27864));
    defparam \scaler_3.un2_source_data_0_cry_1_c_RNO_LC_10_14_3 .C_ON=1'b0;
    defparam \scaler_3.un2_source_data_0_cry_1_c_RNO_LC_10_14_3 .SEQ_MODE=4'b0000;
    defparam \scaler_3.un2_source_data_0_cry_1_c_RNO_LC_10_14_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \scaler_3.un2_source_data_0_cry_1_c_RNO_LC_10_14_3  (
            .in0(N__29014),
            .in1(N__28981),
            .in2(_gnd_net_),
            .in3(N__28945),
            .lcout(\scaler_3.un2_source_data_0_cry_1_c_RNO_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_ns_i_a2_1_1_0_LC_10_14_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_ns_i_a2_1_1_0_LC_10_14_5 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_ns_i_a2_1_1_0_LC_10_14_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \Commands_frame_decoder.state_ns_i_a2_1_1_0_LC_10_14_5  (
            .in0(_gnd_net_),
            .in1(N__44263),
            .in2(_gnd_net_),
            .in3(N__45001),
            .lcout(\Commands_frame_decoder.state_ns_i_a2_1_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI9S511_5_LC_10_14_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI9S511_5_LC_10_14_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI9S511_5_LC_10_14_6 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI9S511_5_LC_10_14_6  (
            .in0(N__25847),
            .in1(N__25823),
            .in2(_gnd_net_),
            .in3(N__25802),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI9S511Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIRFO19_3_LC_10_15_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIRFO19_3_LC_10_15_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIRFO19_3_LC_10_15_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIRFO19_3_LC_10_15_0  (
            .in0(N__26075),
            .in1(N__29947),
            .in2(N__26118),
            .in3(N__26058),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIRFO19Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNICISB3_3_LC_10_15_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNICISB3_3_LC_10_15_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNICISB3_3_LC_10_15_2 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNICISB3_3_LC_10_15_2  (
            .in0(N__26076),
            .in1(N__26057),
            .in2(_gnd_net_),
            .in3(N__29948),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNICISB3Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_4_LC_10_15_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_4_LC_10_15_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_4_LC_10_15_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_4_LC_10_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45495),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47317),
            .ce(N__33598),
            .sr(N__43837));
    defparam \pid_alt.error_i_acumm_prereg_esr_4_LC_10_15_5 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_4_LC_10_15_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_4_LC_10_15_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_4_LC_10_15_5  (
            .in0(N__29949),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_i_acumm7lto4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47317),
            .ce(N__33598),
            .sr(N__43837));
    defparam \pid_alt.error_i_acumm_prereg_esr_5_LC_10_15_7 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_5_LC_10_15_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_5_LC_10_15_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_5_LC_10_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29910),
            .lcout(\pid_alt.error_i_acumm7lto5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47317),
            .ce(N__33598),
            .sr(N__43837));
    defparam \Commands_frame_decoder.source_CH4data_esr_1_LC_10_16_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH4data_esr_1_LC_10_16_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH4data_esr_1_LC_10_16_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH4data_esr_1_LC_10_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45214),
            .lcout(frame_decoder_CH4data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47306),
            .ce(N__26383),
            .sr(N__43845));
    defparam \Commands_frame_decoder.source_CH4data_esr_2_LC_10_16_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH4data_esr_2_LC_10_16_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH4data_esr_2_LC_10_16_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH4data_esr_2_LC_10_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36865),
            .lcout(frame_decoder_CH4data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47306),
            .ce(N__26383),
            .sr(N__43845));
    defparam \Commands_frame_decoder.source_CH4data_esr_3_LC_10_16_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH4data_esr_3_LC_10_16_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH4data_esr_3_LC_10_16_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH4data_esr_3_LC_10_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43349),
            .lcout(frame_decoder_CH4data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47306),
            .ce(N__26383),
            .sr(N__43845));
    defparam \Commands_frame_decoder.source_CH4data_esr_0_LC_10_16_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH4data_esr_0_LC_10_16_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH4data_esr_0_LC_10_16_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH4data_esr_0_LC_10_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27669),
            .lcout(frame_decoder_CH4data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47306),
            .ce(N__26383),
            .sr(N__43845));
    defparam \Commands_frame_decoder.source_CH4data_esr_6_LC_10_16_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH4data_esr_6_LC_10_16_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH4data_esr_6_LC_10_16_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH4data_esr_6_LC_10_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33409),
            .lcout(frame_decoder_CH4data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47306),
            .ce(N__26383),
            .sr(N__43845));
    defparam \Commands_frame_decoder.source_CH4data_ess_7_LC_10_16_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH4data_ess_7_LC_10_16_7 .SEQ_MODE=4'b1001;
    defparam \Commands_frame_decoder.source_CH4data_ess_7_LC_10_16_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH4data_ess_7_LC_10_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45005),
            .lcout(frame_decoder_CH4data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47306),
            .ce(N__26383),
            .sr(N__43845));
    defparam CONSTANT_ONE_LUT4_LC_10_17_2.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_10_17_2.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_10_17_2.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_10_17_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_CH1data8lto3_LC_10_17_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH1data8lto3_LC_10_17_3 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.source_CH1data8lto3_LC_10_17_3 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \Commands_frame_decoder.source_CH1data8lto3_LC_10_17_3  (
            .in0(N__43342),
            .in1(N__36857),
            .in2(_gnd_net_),
            .in3(N__45204),
            .lcout(\Commands_frame_decoder.source_CH1data8lt7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIUI2T2_6_LC_10_17_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIUI2T2_6_LC_10_17_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIUI2T2_6_LC_10_17_5 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIUI2T2_6_LC_10_17_5  (
            .in0(N__26352),
            .in1(N__26328),
            .in2(_gnd_net_),
            .in3(N__30479),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIUI2T2Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIGQS34_23_LC_10_18_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIGQS34_23_LC_10_18_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIGQS34_23_LC_10_18_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIGQS34_23_LC_10_18_6  (
            .in0(N__26286),
            .in1(N__26279),
            .in2(N__26250),
            .in3(N__30705),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIGQS34Z0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_11_LC_10_19_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_11_LC_10_19_1 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_11_LC_10_19_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_11_LC_10_19_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26205),
            .lcout(\dron_frame_decoder_1.drone_altitude_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47283),
            .ce(N__26147),
            .sr(N__43866));
    defparam \pid_alt.error_i_acumm_prereg_esr_7_LC_10_21_0 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_7_LC_10_21_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_7_LC_10_21_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_7_LC_10_21_0  (
            .in0(N__30475),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47270),
            .ce(N__33618),
            .sr(N__43880));
    defparam \pid_alt.error_i_acumm_prereg_esr_15_LC_10_21_5 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_15_LC_10_21_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_15_LC_10_21_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_15_LC_10_21_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30944),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47270),
            .ce(N__33618),
            .sr(N__43880));
    defparam \pid_alt.error_i_acumm_prereg_esr_6_LC_10_21_6 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_6_LC_10_21_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_6_LC_10_21_6 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_6_LC_10_21_6  (
            .in0(_gnd_net_),
            .in1(N__29870),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47270),
            .ce(N__33618),
            .sr(N__43880));
    defparam \uart_pc_sync.Q_0__0_LC_11_5_5 .C_ON=1'b0;
    defparam \uart_pc_sync.Q_0__0_LC_11_5_5 .SEQ_MODE=4'b1000;
    defparam \uart_pc_sync.Q_0__0_LC_11_5_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_pc_sync.Q_0__0_LC_11_5_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26421),
            .lcout(debug_CH2_18A_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47434),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNIRP8S_1_LC_11_6_0 .C_ON=1'b1;
    defparam \uart_pc.timer_Count_RNIRP8S_1_LC_11_6_0 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNIRP8S_1_LC_11_6_0 .LUT_INIT=16'b0001000100010001;
    LogicCell40 \uart_pc.timer_Count_RNIRP8S_1_LC_11_6_0  (
            .in0(N__26535),
            .in1(N__26510),
            .in2(N__26538),
            .in3(_gnd_net_),
            .lcout(\uart_pc.un1_state_2_0_a3_0 ),
            .ltout(),
            .carryin(bfn_11_6_0_),
            .carryout(\uart_pc.un4_timer_Count_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNO_0_2_LC_11_6_1 .C_ON=1'b1;
    defparam \uart_pc.timer_Count_RNO_0_2_LC_11_6_1 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNO_0_2_LC_11_6_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \uart_pc.timer_Count_RNO_0_2_LC_11_6_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__27495),
            .in3(N__26415),
            .lcout(\uart_pc.timer_Count_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(\uart_pc.un4_timer_Count_1_cry_1 ),
            .carryout(\uart_pc.un4_timer_Count_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNO_0_3_LC_11_6_2 .C_ON=1'b1;
    defparam \uart_pc.timer_Count_RNO_0_3_LC_11_6_2 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNO_0_3_LC_11_6_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \uart_pc.timer_Count_RNO_0_3_LC_11_6_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__31615),
            .in3(N__26412),
            .lcout(\uart_pc.timer_Count_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(\uart_pc.un4_timer_Count_1_cry_2 ),
            .carryout(\uart_pc.un4_timer_Count_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNO_0_4_LC_11_6_3 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_RNO_0_4_LC_11_6_3 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNO_0_4_LC_11_6_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uart_pc.timer_Count_RNO_0_4_LC_11_6_3  (
            .in0(_gnd_net_),
            .in1(N__31489),
            .in2(_gnd_net_),
            .in3(N__26409),
            .lcout(\uart_pc.timer_Count_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_2_LC_11_6_4 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_2_LC_11_6_4 .SEQ_MODE=4'b1000;
    defparam \uart_pc.timer_Count_2_LC_11_6_4 .LUT_INIT=16'b0101010000000000;
    LogicCell40 \uart_pc.timer_Count_2_LC_11_6_4  (
            .in0(N__44104),
            .in1(N__27462),
            .in2(N__27555),
            .in3(N__26406),
            .lcout(\uart_pc.timer_CountZ1Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47424),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_0_LC_11_6_5 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_0_LC_11_6_5 .SEQ_MODE=4'b1000;
    defparam \uart_pc.timer_Count_0_LC_11_6_5 .LUT_INIT=16'b0000000001010100;
    LogicCell40 \uart_pc.timer_Count_0_LC_11_6_5  (
            .in0(N__26537),
            .in1(N__27547),
            .in2(N__27467),
            .in3(N__44105),
            .lcout(\uart_pc.timer_CountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47424),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNIPD2K1_2_LC_11_6_6 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_RNIPD2K1_2_LC_11_6_6 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNIPD2K1_2_LC_11_6_6 .LUT_INIT=16'b1111100000000000;
    LogicCell40 \uart_pc.timer_Count_RNIPD2K1_2_LC_11_6_6  (
            .in0(N__31601),
            .in1(N__27490),
            .in2(N__31505),
            .in3(N__31546),
            .lcout(\uart_pc.data_rdyc_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_RNIMQ8T1_4_LC_11_6_7 .C_ON=1'b0;
    defparam \uart_pc.state_RNIMQ8T1_4_LC_11_6_7 .SEQ_MODE=4'b0000;
    defparam \uart_pc.state_RNIMQ8T1_4_LC_11_6_7 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \uart_pc.state_RNIMQ8T1_4_LC_11_6_7  (
            .in0(N__31547),
            .in1(N__31271),
            .in2(N__44135),
            .in3(N__31490),
            .lcout(\uart_pc.N_143 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNIMQ8T1_2_LC_11_7_1 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_RNIMQ8T1_2_LC_11_7_1 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNIMQ8T1_2_LC_11_7_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \uart_pc.timer_Count_RNIMQ8T1_2_LC_11_7_1  (
            .in0(_gnd_net_),
            .in1(N__26574),
            .in2(_gnd_net_),
            .in3(N__44079),
            .lcout(\uart_pc.timer_Count_RNIMQ8T1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_4_LC_11_7_3 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_4_LC_11_7_3 .SEQ_MODE=4'b1000;
    defparam \uart_pc.timer_Count_4_LC_11_7_3 .LUT_INIT=16'b0000000011001000;
    LogicCell40 \uart_pc.timer_Count_4_LC_11_7_3  (
            .in0(N__27553),
            .in1(N__26544),
            .in2(N__27468),
            .in3(N__44081),
            .lcout(\uart_pc.timer_CountZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47413),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNO_0_1_LC_11_7_5 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_RNO_0_1_LC_11_7_5 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNO_0_1_LC_11_7_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart_pc.timer_Count_RNO_0_1_LC_11_7_5  (
            .in0(_gnd_net_),
            .in1(N__26536),
            .in2(_gnd_net_),
            .in3(N__26511),
            .lcout(),
            .ltout(\uart_pc.timer_Count_RNO_0Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_1_LC_11_7_6 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_1_LC_11_7_6 .SEQ_MODE=4'b1000;
    defparam \uart_pc.timer_Count_1_LC_11_7_6 .LUT_INIT=16'b0101000001000000;
    LogicCell40 \uart_pc.timer_Count_1_LC_11_7_6  (
            .in0(N__44080),
            .in1(N__27463),
            .in2(N__26514),
            .in3(N__27552),
            .lcout(\uart_pc.timer_CountZ1Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47413),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_ns_0_a4_0_0_1_LC_11_8_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_ns_0_a4_0_0_1_LC_11_8_1 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_ns_0_a4_0_0_1_LC_11_8_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Commands_frame_decoder.state_ns_0_a4_0_0_1_LC_11_8_1  (
            .in0(_gnd_net_),
            .in1(N__44914),
            .in2(_gnd_net_),
            .in3(N__27613),
            .lcout(\Commands_frame_decoder.state_ns_0_a4_0_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNIVGCQ_12_LC_11_8_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIVGCQ_12_LC_11_8_2 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIVGCQ_12_LC_11_8_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \Commands_frame_decoder.state_RNIVGCQ_12_LC_11_8_2  (
            .in0(N__26953),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26484),
            .lcout(\Commands_frame_decoder.state_ns_i_a4_2_0_0 ),
            .ltout(\Commands_frame_decoder.state_ns_i_a4_2_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.count_0_LC_11_8_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.count_0_LC_11_8_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.count_0_LC_11_8_3 .LUT_INIT=16'b0000000000111100;
    LogicCell40 \Commands_frame_decoder.count_0_LC_11_8_3  (
            .in0(_gnd_net_),
            .in1(N__26650),
            .in2(N__26487),
            .in3(N__44107),
            .lcout(\Commands_frame_decoder.countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47402),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.count_RNI0V5H1_1_LC_11_8_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.count_RNI0V5H1_1_LC_11_8_4 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.count_RNI0V5H1_1_LC_11_8_4 .LUT_INIT=16'b0111000000000000;
    LogicCell40 \Commands_frame_decoder.count_RNI0V5H1_1_LC_11_8_4  (
            .in0(N__26649),
            .in1(N__26632),
            .in2(N__26999),
            .in3(N__26483),
            .lcout(\Commands_frame_decoder.N_330 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.reset_LC_11_8_5 .C_ON=1'b0;
    defparam \reset_module_System.reset_LC_11_8_5 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.reset_LC_11_8_5 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \reset_module_System.reset_LC_11_8_5  (
            .in0(N__33840),
            .in1(N__37320),
            .in2(_gnd_net_),
            .in3(N__33791),
            .lcout(reset_system),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47402),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.count_1_LC_11_8_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.count_1_LC_11_8_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.count_1_LC_11_8_6 .LUT_INIT=16'b0001010101000000;
    LogicCell40 \Commands_frame_decoder.count_1_LC_11_8_6  (
            .in0(N__44106),
            .in1(N__26430),
            .in2(N__26655),
            .in3(N__26633),
            .lcout(\Commands_frame_decoder.countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47402),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_0_LC_11_8_7 .C_ON=1'b0;
    defparam \uart_pc.data_0_LC_11_8_7 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_0_LC_11_8_7 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \uart_pc.data_0_LC_11_8_7  (
            .in0(N__31060),
            .in1(N__30992),
            .in2(N__28878),
            .in3(N__27614),
            .lcout(uart_pc_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47402),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_3.un3_source_data_un3_source_data_0_axb_7_LC_11_9_0 .C_ON=1'b0;
    defparam \scaler_3.un3_source_data_un3_source_data_0_axb_7_LC_11_9_0 .SEQ_MODE=4'b0000;
    defparam \scaler_3.un3_source_data_un3_source_data_0_axb_7_LC_11_9_0 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \scaler_3.un3_source_data_un3_source_data_0_axb_7_LC_11_9_0  (
            .in0(_gnd_net_),
            .in1(N__26708),
            .in2(_gnd_net_),
            .in3(N__26685),
            .lcout(\scaler_3.un3_source_data_0_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_0_LC_11_9_3 .C_ON=1'b0;
    defparam \reset_module_System.count_0_LC_11_9_3 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_0_LC_11_9_3 .LUT_INIT=16'b1000000011111111;
    LogicCell40 \reset_module_System.count_0_LC_11_9_3  (
            .in0(N__37319),
            .in1(N__33786),
            .in2(N__33849),
            .in3(N__34818),
            .lcout(\reset_module_System.countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47387),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_4_LC_11_9_4 .C_ON=1'b0;
    defparam \uart_pc.data_4_LC_11_9_4 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_4_LC_11_9_4 .LUT_INIT=16'b0011000100100000;
    LogicCell40 \uart_pc.data_4_LC_11_9_4  (
            .in0(N__26586),
            .in1(N__31043),
            .in2(N__28824),
            .in3(N__45297),
            .lcout(uart_pc_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47387),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_RNIES9Q1_2_LC_11_9_5 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_RNIES9Q1_2_LC_11_9_5 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNIES9Q1_2_LC_11_9_5 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \uart_drone.timer_Count_RNIES9Q1_2_LC_11_9_5  (
            .in0(N__31370),
            .in1(N__31642),
            .in2(_gnd_net_),
            .in3(N__44075),
            .lcout(\uart_drone.timer_Count_RNIES9Q1Z0Z_2 ),
            .ltout(\uart_drone.timer_Count_RNIES9Q1Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_RNIRC5U2_2_LC_11_9_6 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_RNIRC5U2_2_LC_11_9_6 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNIRC5U2_2_LC_11_9_6 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \uart_drone.timer_Count_RNIRC5U2_2_LC_11_9_6  (
            .in0(N__31643),
            .in1(_gnd_net_),
            .in2(N__26604),
            .in3(_gnd_net_),
            .lcout(\uart_drone.data_rdyc_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNILR1B2_2_LC_11_10_2 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_RNILR1B2_2_LC_11_10_2 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNILR1B2_2_LC_11_10_2 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \uart_pc.timer_Count_RNILR1B2_2_LC_11_10_2  (
            .in0(N__31178),
            .in1(N__26584),
            .in2(_gnd_net_),
            .in3(N__44078),
            .lcout(\uart_pc.timer_Count_RNILR1B2Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.data_Aux_RNO_0_0_LC_11_10_3 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_RNO_0_0_LC_11_10_3 .SEQ_MODE=4'b0000;
    defparam \uart_drone.data_Aux_RNO_0_0_LC_11_10_3 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \uart_drone.data_Aux_RNO_0_0_LC_11_10_3  (
            .in0(N__44423),
            .in1(N__36691),
            .in2(_gnd_net_),
            .in3(N__39516),
            .lcout(\uart_drone.data_Auxce_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.data_Aux_RNO_0_1_LC_11_10_4 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_RNO_0_1_LC_11_10_4 .SEQ_MODE=4'b0000;
    defparam \uart_drone.data_Aux_RNO_0_1_LC_11_10_4 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \uart_drone.data_Aux_RNO_0_1_LC_11_10_4  (
            .in0(N__39517),
            .in1(N__36692),
            .in2(_gnd_net_),
            .in3(N__44424),
            .lcout(\uart_drone.data_Auxce_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_3.N_1239_i_l_ofx_LC_11_10_6 .C_ON=1'b0;
    defparam \scaler_3.N_1239_i_l_ofx_LC_11_10_6 .SEQ_MODE=4'b0000;
    defparam \scaler_3.N_1239_i_l_ofx_LC_11_10_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \scaler_3.N_1239_i_l_ofx_LC_11_10_6  (
            .in0(_gnd_net_),
            .in1(N__26709),
            .in2(_gnd_net_),
            .in3(N__26684),
            .lcout(\scaler_3.N_1239_i_l_ofxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_2.un3_source_data_un3_source_data_0_axb_7_LC_11_10_7 .C_ON=1'b0;
    defparam \scaler_2.un3_source_data_un3_source_data_0_axb_7_LC_11_10_7 .SEQ_MODE=4'b0000;
    defparam \scaler_2.un3_source_data_un3_source_data_0_axb_7_LC_11_10_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \scaler_2.un3_source_data_un3_source_data_0_axb_7_LC_11_10_7  (
            .in0(_gnd_net_),
            .in1(N__28103),
            .in2(_gnd_net_),
            .in3(N__28091),
            .lcout(\scaler_2.un3_source_data_0_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_CH2data_esr_0_LC_11_11_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH2data_esr_0_LC_11_11_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH2data_esr_0_LC_11_11_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH2data_esr_0_LC_11_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27651),
            .lcout(frame_decoder_CH2data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47362),
            .ce(N__26670),
            .sr(N__43817));
    defparam \Commands_frame_decoder.source_CH2data_esr_1_LC_11_11_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH2data_esr_1_LC_11_11_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH2data_esr_1_LC_11_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH2data_esr_1_LC_11_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45190),
            .lcout(frame_decoder_CH2data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47362),
            .ce(N__26670),
            .sr(N__43817));
    defparam \Commands_frame_decoder.source_CH2data_esr_2_LC_11_11_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH2data_esr_2_LC_11_11_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH2data_esr_2_LC_11_11_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH2data_esr_2_LC_11_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36856),
            .lcout(frame_decoder_CH2data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47362),
            .ce(N__26670),
            .sr(N__43817));
    defparam \Commands_frame_decoder.source_CH2data_esr_3_LC_11_11_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH2data_esr_3_LC_11_11_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH2data_esr_3_LC_11_11_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Commands_frame_decoder.source_CH2data_esr_3_LC_11_11_3  (
            .in0(N__43312),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(frame_decoder_CH2data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47362),
            .ce(N__26670),
            .sr(N__43817));
    defparam \Commands_frame_decoder.source_CH2data_esr_4_LC_11_11_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH2data_esr_4_LC_11_11_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH2data_esr_4_LC_11_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH2data_esr_4_LC_11_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45313),
            .lcout(frame_decoder_CH2data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47362),
            .ce(N__26670),
            .sr(N__43817));
    defparam \Commands_frame_decoder.source_CH2data_esr_5_LC_11_11_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH2data_esr_5_LC_11_11_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH2data_esr_5_LC_11_11_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH2data_esr_5_LC_11_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44249),
            .lcout(frame_decoder_CH2data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47362),
            .ce(N__26670),
            .sr(N__43817));
    defparam \Commands_frame_decoder.source_CH2data_esr_6_LC_11_11_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH2data_esr_6_LC_11_11_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH2data_esr_6_LC_11_11_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Commands_frame_decoder.source_CH2data_esr_6_LC_11_11_6  (
            .in0(N__33393),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(frame_decoder_CH2data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47362),
            .ce(N__26670),
            .sr(N__43817));
    defparam \Commands_frame_decoder.source_CH2data_ess_7_LC_11_11_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH2data_ess_7_LC_11_11_7 .SEQ_MODE=4'b1001;
    defparam \Commands_frame_decoder.source_CH2data_ess_7_LC_11_11_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Commands_frame_decoder.source_CH2data_ess_7_LC_11_11_7  (
            .in0(N__44982),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(frame_decoder_CH2data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47362),
            .ce(N__26670),
            .sr(N__43817));
    defparam \Commands_frame_decoder.source_offset3data_esr_0_LC_11_12_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset3data_esr_0_LC_11_12_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset3data_esr_0_LC_11_12_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset3data_esr_0_LC_11_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27654),
            .lcout(frame_decoder_OFF3data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47347),
            .ce(N__26751),
            .sr(N__43822));
    defparam \Commands_frame_decoder.source_offset3data_esr_1_LC_11_12_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset3data_esr_1_LC_11_12_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset3data_esr_1_LC_11_12_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset3data_esr_1_LC_11_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45212),
            .lcout(frame_decoder_OFF3data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47347),
            .ce(N__26751),
            .sr(N__43822));
    defparam \Commands_frame_decoder.source_offset3data_esr_2_LC_11_12_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset3data_esr_2_LC_11_12_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset3data_esr_2_LC_11_12_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset3data_esr_2_LC_11_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36872),
            .lcout(frame_decoder_OFF3data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47347),
            .ce(N__26751),
            .sr(N__43822));
    defparam \Commands_frame_decoder.source_offset3data_esr_3_LC_11_12_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset3data_esr_3_LC_11_12_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset3data_esr_3_LC_11_12_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset3data_esr_3_LC_11_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43340),
            .lcout(frame_decoder_OFF3data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47347),
            .ce(N__26751),
            .sr(N__43822));
    defparam \Commands_frame_decoder.source_offset3data_esr_4_LC_11_12_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset3data_esr_4_LC_11_12_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset3data_esr_4_LC_11_12_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Commands_frame_decoder.source_offset3data_esr_4_LC_11_12_4  (
            .in0(N__45330),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(frame_decoder_OFF3data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47347),
            .ce(N__26751),
            .sr(N__43822));
    defparam \Commands_frame_decoder.source_offset3data_esr_5_LC_11_12_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset3data_esr_5_LC_11_12_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset3data_esr_5_LC_11_12_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset3data_esr_5_LC_11_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44250),
            .lcout(frame_decoder_OFF3data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47347),
            .ce(N__26751),
            .sr(N__43822));
    defparam \Commands_frame_decoder.source_offset3data_esr_6_LC_11_12_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset3data_esr_6_LC_11_12_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset3data_esr_6_LC_11_12_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset3data_esr_6_LC_11_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33394),
            .lcout(frame_decoder_OFF3data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47347),
            .ce(N__26751),
            .sr(N__43822));
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_0_c_LC_11_13_0 .C_ON=1'b1;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_0_c_LC_11_13_0 .SEQ_MODE=4'b0000;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_0_c_LC_11_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \scaler_3.un3_source_data_un3_source_data_0_cry_0_c_LC_11_13_0  (
            .in0(_gnd_net_),
            .in1(N__28944),
            .in2(N__28980),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_13_0_),
            .carryout(\scaler_3.un3_source_data_0_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_0_c_RNI10UK_LC_11_13_1 .C_ON=1'b1;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_0_c_RNI10UK_LC_11_13_1 .SEQ_MODE=4'b0000;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_0_c_RNI10UK_LC_11_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_3.un3_source_data_un3_source_data_0_cry_0_c_RNI10UK_LC_11_13_1  (
            .in0(_gnd_net_),
            .in1(N__26733),
            .in2(N__26727),
            .in3(N__26712),
            .lcout(\scaler_3.un2_source_data_0 ),
            .ltout(),
            .carryin(\scaler_3.un3_source_data_0_cry_0 ),
            .carryout(\scaler_3.un3_source_data_0_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_1_c_RNI44VK_LC_11_13_2 .C_ON=1'b1;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_1_c_RNI44VK_LC_11_13_2 .SEQ_MODE=4'b0000;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_1_c_RNI44VK_LC_11_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_3.un3_source_data_un3_source_data_0_cry_1_c_RNI44VK_LC_11_13_2  (
            .in0(_gnd_net_),
            .in1(N__26895),
            .in2(N__26886),
            .in3(N__26877),
            .lcout(\scaler_3.un3_source_data_0_cry_1_c_RNI44VK ),
            .ltout(),
            .carryin(\scaler_3.un3_source_data_0_cry_1 ),
            .carryout(\scaler_3.un3_source_data_0_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_2_c_RNI780L_LC_11_13_3 .C_ON=1'b1;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_2_c_RNI780L_LC_11_13_3 .SEQ_MODE=4'b0000;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_2_c_RNI780L_LC_11_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_3.un3_source_data_un3_source_data_0_cry_2_c_RNI780L_LC_11_13_3  (
            .in0(_gnd_net_),
            .in1(N__26874),
            .in2(N__26865),
            .in3(N__26856),
            .lcout(\scaler_3.un3_source_data_0_cry_2_c_RNI780L ),
            .ltout(),
            .carryin(\scaler_3.un3_source_data_0_cry_2 ),
            .carryout(\scaler_3.un3_source_data_0_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_3_c_RNIAC1L_LC_11_13_4 .C_ON=1'b1;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_3_c_RNIAC1L_LC_11_13_4 .SEQ_MODE=4'b0000;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_3_c_RNIAC1L_LC_11_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_3.un3_source_data_un3_source_data_0_cry_3_c_RNIAC1L_LC_11_13_4  (
            .in0(_gnd_net_),
            .in1(N__26853),
            .in2(N__26841),
            .in3(N__26832),
            .lcout(\scaler_3.un3_source_data_0_cry_3_c_RNIAC1L ),
            .ltout(),
            .carryin(\scaler_3.un3_source_data_0_cry_3 ),
            .carryout(\scaler_3.un3_source_data_0_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_4_c_RNIDG2L_LC_11_13_5 .C_ON=1'b1;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_4_c_RNIDG2L_LC_11_13_5 .SEQ_MODE=4'b0000;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_4_c_RNIDG2L_LC_11_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_3.un3_source_data_un3_source_data_0_cry_4_c_RNIDG2L_LC_11_13_5  (
            .in0(_gnd_net_),
            .in1(N__26829),
            .in2(N__26817),
            .in3(N__26805),
            .lcout(\scaler_3.un3_source_data_0_cry_4_c_RNIDG2L ),
            .ltout(),
            .carryin(\scaler_3.un3_source_data_0_cry_4 ),
            .carryout(\scaler_3.un3_source_data_0_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_5_c_RNIGK3L_LC_11_13_6 .C_ON=1'b1;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_5_c_RNIGK3L_LC_11_13_6 .SEQ_MODE=4'b0000;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_5_c_RNIGK3L_LC_11_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_3.un3_source_data_un3_source_data_0_cry_5_c_RNIGK3L_LC_11_13_6  (
            .in0(_gnd_net_),
            .in1(N__26802),
            .in2(N__26790),
            .in3(N__26781),
            .lcout(\scaler_3.un3_source_data_0_cry_5_c_RNIGK3L ),
            .ltout(),
            .carryin(\scaler_3.un3_source_data_0_cry_5 ),
            .carryout(\scaler_3.un3_source_data_0_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_6_c_RNILUAN_LC_11_13_7 .C_ON=1'b1;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_6_c_RNILUAN_LC_11_13_7 .SEQ_MODE=4'b0000;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_6_c_RNILUAN_LC_11_13_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \scaler_3.un3_source_data_un3_source_data_0_cry_6_c_RNILUAN_LC_11_13_7  (
            .in0(_gnd_net_),
            .in1(N__26778),
            .in2(_gnd_net_),
            .in3(N__26769),
            .lcout(\scaler_3.un3_source_data_0_cry_6_c_RNILUAN ),
            .ltout(),
            .carryin(\scaler_3.un3_source_data_0_cry_6 ),
            .carryout(\scaler_3.un3_source_data_0_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_7_c_RNIM0CN_LC_11_14_0 .C_ON=1'b1;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_7_c_RNIM0CN_LC_11_14_0 .SEQ_MODE=4'b0000;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_7_c_RNIM0CN_LC_11_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_3.un3_source_data_un3_source_data_0_cry_7_c_RNIM0CN_LC_11_14_0  (
            .in0(_gnd_net_),
            .in1(N__26766),
            .in2(N__42916),
            .in3(N__26757),
            .lcout(\scaler_3.un3_source_data_0_cry_7_c_RNIM0CN ),
            .ltout(),
            .carryin(bfn_11_14_0_),
            .carryout(\scaler_3.un3_source_data_0_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_8_c_RNIRV25_LC_11_14_1 .C_ON=1'b0;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_8_c_RNIRV25_LC_11_14_1 .SEQ_MODE=4'b0000;
    defparam \scaler_3.un3_source_data_un3_source_data_0_cry_8_c_RNIRV25_LC_11_14_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \scaler_3.un3_source_data_un3_source_data_0_cry_8_c_RNIRV25_LC_11_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26754),
            .lcout(\scaler_3.un3_source_data_0_cry_8_c_RNIRV25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNI7G141_10_LC_11_14_2 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNI7G141_10_LC_11_14_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNI7G141_10_LC_11_14_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \pid_alt.pid_prereg_esr_RNI7G141_10_LC_11_14_2  (
            .in0(N__27166),
            .in1(N__27947),
            .in2(N__27141),
            .in3(N__27104),
            .lcout(\pid_alt.source_pid_1_sqmuxa_0_a2_2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNILP1J_9_LC_11_14_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNILP1J_9_LC_11_14_5 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNILP1J_9_LC_11_14_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Commands_frame_decoder.state_RNILP1J_9_LC_11_14_5  (
            .in0(_gnd_net_),
            .in1(N__27066),
            .in2(_gnd_net_),
            .in3(N__27042),
            .lcout(\Commands_frame_decoder.source_offset4data_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_offset4data_esr_0_LC_11_15_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset4data_esr_0_LC_11_15_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset4data_esr_0_LC_11_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset4data_esr_0_LC_11_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27655),
            .lcout(frame_decoder_OFF4data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47307),
            .ce(N__27327),
            .sr(N__43846));
    defparam \Commands_frame_decoder.source_offset4data_esr_1_LC_11_15_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset4data_esr_1_LC_11_15_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset4data_esr_1_LC_11_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset4data_esr_1_LC_11_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45213),
            .lcout(frame_decoder_OFF4data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47307),
            .ce(N__27327),
            .sr(N__43846));
    defparam \Commands_frame_decoder.source_offset4data_esr_2_LC_11_15_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset4data_esr_2_LC_11_15_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset4data_esr_2_LC_11_15_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset4data_esr_2_LC_11_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36873),
            .lcout(frame_decoder_OFF4data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47307),
            .ce(N__27327),
            .sr(N__43846));
    defparam \Commands_frame_decoder.source_offset4data_esr_3_LC_11_15_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset4data_esr_3_LC_11_15_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset4data_esr_3_LC_11_15_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset4data_esr_3_LC_11_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43341),
            .lcout(frame_decoder_OFF4data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47307),
            .ce(N__27327),
            .sr(N__43846));
    defparam \Commands_frame_decoder.source_offset4data_esr_4_LC_11_15_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset4data_esr_4_LC_11_15_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset4data_esr_4_LC_11_15_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset4data_esr_4_LC_11_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45331),
            .lcout(frame_decoder_OFF4data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47307),
            .ce(N__27327),
            .sr(N__43846));
    defparam \Commands_frame_decoder.source_offset4data_esr_5_LC_11_15_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset4data_esr_5_LC_11_15_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset4data_esr_5_LC_11_15_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset4data_esr_5_LC_11_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44270),
            .lcout(frame_decoder_OFF4data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47307),
            .ce(N__27327),
            .sr(N__43846));
    defparam \Commands_frame_decoder.source_offset4data_esr_6_LC_11_15_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset4data_esr_6_LC_11_15_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset4data_esr_6_LC_11_15_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset4data_esr_6_LC_11_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33413),
            .lcout(frame_decoder_OFF4data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47307),
            .ce(N__27327),
            .sr(N__43846));
    defparam \Commands_frame_decoder.source_offset4data_ess_7_LC_11_15_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset4data_ess_7_LC_11_15_7 .SEQ_MODE=4'b1001;
    defparam \Commands_frame_decoder.source_offset4data_ess_7_LC_11_15_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset4data_ess_7_LC_11_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44988),
            .lcout(frame_decoder_OFF4data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47307),
            .ce(N__27327),
            .sr(N__43846));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_LC_11_16_0 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_LC_11_16_0 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_LC_11_16_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_LC_11_16_0  (
            .in0(_gnd_net_),
            .in1(N__29493),
            .in2(N__29550),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_16_0_),
            .carryout(\scaler_4.un3_source_data_0_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_RNI40BL_LC_11_16_1 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_RNI40BL_LC_11_16_1 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_RNI40BL_LC_11_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_RNI40BL_LC_11_16_1  (
            .in0(_gnd_net_),
            .in1(N__27309),
            .in2(N__27303),
            .in3(N__27294),
            .lcout(\scaler_4.un2_source_data_0 ),
            .ltout(),
            .carryin(\scaler_4.un3_source_data_0_cry_0 ),
            .carryout(\scaler_4.un3_source_data_0_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_1_c_RNI74CL_LC_11_16_2 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_1_c_RNI74CL_LC_11_16_2 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_1_c_RNI74CL_LC_11_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_1_c_RNI74CL_LC_11_16_2  (
            .in0(_gnd_net_),
            .in1(N__27291),
            .in2(N__27285),
            .in3(N__27273),
            .lcout(\scaler_4.un3_source_data_0_cry_1_c_RNI74CL ),
            .ltout(),
            .carryin(\scaler_4.un3_source_data_0_cry_1 ),
            .carryout(\scaler_4.un3_source_data_0_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_2_c_RNIA8DL_LC_11_16_3 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_2_c_RNIA8DL_LC_11_16_3 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_2_c_RNIA8DL_LC_11_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_2_c_RNIA8DL_LC_11_16_3  (
            .in0(_gnd_net_),
            .in1(N__27270),
            .in2(N__27264),
            .in3(N__27255),
            .lcout(\scaler_4.un3_source_data_0_cry_2_c_RNIA8DL ),
            .ltout(),
            .carryin(\scaler_4.un3_source_data_0_cry_2 ),
            .carryout(\scaler_4.un3_source_data_0_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_3_c_RNIDCEL_LC_11_16_4 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_3_c_RNIDCEL_LC_11_16_4 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_3_c_RNIDCEL_LC_11_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_3_c_RNIDCEL_LC_11_16_4  (
            .in0(_gnd_net_),
            .in1(N__27252),
            .in2(N__27237),
            .in3(N__27228),
            .lcout(\scaler_4.un3_source_data_0_cry_3_c_RNIDCEL ),
            .ltout(),
            .carryin(\scaler_4.un3_source_data_0_cry_3 ),
            .carryout(\scaler_4.un3_source_data_0_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_4_c_RNIGGFL_LC_11_16_5 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_4_c_RNIGGFL_LC_11_16_5 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_4_c_RNIGGFL_LC_11_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_4_c_RNIGGFL_LC_11_16_5  (
            .in0(_gnd_net_),
            .in1(N__27225),
            .in2(N__27219),
            .in3(N__27201),
            .lcout(\scaler_4.un3_source_data_0_cry_4_c_RNIGGFL ),
            .ltout(),
            .carryin(\scaler_4.un3_source_data_0_cry_4 ),
            .carryout(\scaler_4.un3_source_data_0_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_5_c_RNIJKGL_LC_11_16_6 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_5_c_RNIJKGL_LC_11_16_6 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_5_c_RNIJKGL_LC_11_16_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_5_c_RNIJKGL_LC_11_16_6  (
            .in0(_gnd_net_),
            .in1(N__27198),
            .in2(N__27192),
            .in3(N__27183),
            .lcout(\scaler_4.un3_source_data_0_cry_5_c_RNIJKGL ),
            .ltout(),
            .carryin(\scaler_4.un3_source_data_0_cry_5 ),
            .carryout(\scaler_4.un3_source_data_0_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_6_c_RNIOUNN_LC_11_16_7 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_6_c_RNIOUNN_LC_11_16_7 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_6_c_RNIOUNN_LC_11_16_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_6_c_RNIOUNN_LC_11_16_7  (
            .in0(_gnd_net_),
            .in1(N__27384),
            .in2(_gnd_net_),
            .in3(N__27180),
            .lcout(\scaler_4.un3_source_data_0_cry_6_c_RNIOUNN ),
            .ltout(),
            .carryin(\scaler_4.un3_source_data_0_cry_6 ),
            .carryout(\scaler_4.un3_source_data_0_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_7_c_RNIP0PN_LC_11_17_0 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_7_c_RNIP0PN_LC_11_17_0 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_7_c_RNIP0PN_LC_11_17_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_7_c_RNIP0PN_LC_11_17_0  (
            .in0(_gnd_net_),
            .in1(N__27354),
            .in2(N__42841),
            .in3(N__27390),
            .lcout(\scaler_4.un3_source_data_0_cry_7_c_RNIP0PN ),
            .ltout(),
            .carryin(bfn_11_17_0_),
            .carryout(\scaler_4.un3_source_data_0_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_8_c_RNIS918_LC_11_17_1 .C_ON=1'b0;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_8_c_RNIS918_LC_11_17_1 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_8_c_RNIS918_LC_11_17_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_8_c_RNIS918_LC_11_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27387),
            .lcout(\scaler_4.un3_source_data_0_cry_8_c_RNIS918 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_axb_7_LC_11_17_2 .C_ON=1'b0;
    defparam \scaler_4.un3_source_data_un3_source_data_0_axb_7_LC_11_17_2 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_axb_7_LC_11_17_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_axb_7_LC_11_17_2  (
            .in0(_gnd_net_),
            .in1(N__27365),
            .in2(_gnd_net_),
            .in3(N__27377),
            .lcout(\scaler_4.un3_source_data_0_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.N_1251_i_l_ofx_LC_11_17_3 .C_ON=1'b0;
    defparam \scaler_4.N_1251_i_l_ofx_LC_11_17_3 .SEQ_MODE=4'b0000;
    defparam \scaler_4.N_1251_i_l_ofx_LC_11_17_3 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \scaler_4.N_1251_i_l_ofx_LC_11_17_3  (
            .in0(N__27378),
            .in1(_gnd_net_),
            .in2(N__27369),
            .in3(_gnd_net_),
            .lcout(\scaler_4.N_1251_i_l_ofxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNII68S_9_LC_11_17_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNII68S_9_LC_11_17_7 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNII68S_9_LC_11_17_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \Commands_frame_decoder.state_RNII68S_9_LC_11_17_7  (
            .in0(_gnd_net_),
            .in1(N__27341),
            .in2(_gnd_net_),
            .in3(N__44091),
            .lcout(\Commands_frame_decoder.source_offset4data_1_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_1_LC_11_19_0 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_1_LC_11_19_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_1_LC_11_19_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_1_LC_11_19_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30085),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47275),
            .ce(N__33606),
            .sr(N__43875));
    defparam \pid_alt.error_i_acumm_prereg_esr_16_LC_11_19_6 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_16_LC_11_19_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_16_LC_11_19_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_16_LC_11_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30913),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47275),
            .ce(N__33606),
            .sr(N__43875));
    defparam \pid_alt.error_i_acumm_prereg_esr_11_LC_11_19_7 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_11_LC_11_19_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_11_LC_11_19_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_11_LC_11_19_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30298),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47275),
            .ce(N__33606),
            .sr(N__43875));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIIDE4_16_LC_11_20_0 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIIDE4_16_LC_11_20_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIIDE4_16_LC_11_20_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNIIDE4_16_LC_11_20_0  (
            .in0(N__27423),
            .in1(N__27402),
            .in2(N__27417),
            .in3(N__27315),
            .lcout(),
            .ltout(\pid_alt.m7_e_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIRRP7_14_LC_11_20_1 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIRRP7_14_LC_11_20_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIRRP7_14_LC_11_20_1 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNIRRP7_14_LC_11_20_1  (
            .in0(N__27396),
            .in1(N__27435),
            .in2(N__27429),
            .in3(N__27408),
            .lcout(\pid_alt.N_238 ),
            .ltout(\pid_alt.N_238_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI175B_12_LC_11_20_2 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI175B_12_LC_11_20_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI175B_12_LC_11_20_2 .LUT_INIT=16'b1011101011111010;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNI175B_12_LC_11_20_2  (
            .in0(N__32845),
            .in1(N__28595),
            .in2(N__27426),
            .in3(N__32822),
            .lcout(\pid_alt.N_128 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_18_LC_11_20_5 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_18_LC_11_20_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_18_LC_11_20_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_18_LC_11_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30839),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47271),
            .ce(N__33609),
            .sr(N__43881));
    defparam \pid_alt.error_i_acumm_prereg_esr_19_LC_11_20_6 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_19_LC_11_20_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_19_LC_11_20_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_19_LC_11_20_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30800),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47271),
            .ce(N__33609),
            .sr(N__43881));
    defparam \pid_alt.error_i_acumm_prereg_esr_14_LC_11_20_7 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_14_LC_11_20_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_14_LC_11_20_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_14_LC_11_20_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30179),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47271),
            .ce(N__33609),
            .sr(N__43881));
    defparam \pid_alt.error_i_acumm_prereg_esr_2_LC_11_21_1 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_2_LC_11_21_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_2_LC_11_21_1 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_2_LC_11_21_1  (
            .in0(_gnd_net_),
            .in1(N__30028),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47268),
            .ce(N__33614),
            .sr(N__43885));
    defparam \pid_alt.error_i_acumm_prereg_esr_17_LC_11_21_2 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_17_LC_11_21_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_17_LC_11_21_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_17_LC_11_21_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30875),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47268),
            .ce(N__33614),
            .sr(N__43885));
    defparam \pid_alt.error_i_acumm_prereg_esr_20_LC_11_21_3 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_20_LC_11_21_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_20_LC_11_21_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_20_LC_11_21_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30766),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47268),
            .ce(N__33614),
            .sr(N__43885));
    defparam \pid_alt.error_i_acumm_prereg_esr_12_LC_11_21_4 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_12_LC_11_21_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_12_LC_11_21_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_12_LC_11_21_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30254),
            .lcout(\pid_alt.error_i_acumm7lto12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47268),
            .ce(N__33614),
            .sr(N__43885));
    defparam \pid_alt.error_i_acumm_prereg_esr_10_LC_11_21_5 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_10_LC_11_21_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_10_LC_11_21_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_10_LC_11_21_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30334),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47268),
            .ce(N__33614),
            .sr(N__43885));
    defparam \pid_alt.error_i_acumm_prereg_esr_21_LC_11_21_6 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_21_LC_11_21_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_21_LC_11_21_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_21_LC_11_21_6  (
            .in0(N__30690),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47268),
            .ce(N__33614),
            .sr(N__43885));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIE3BQ1_0_6_LC_11_22_0 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIE3BQ1_0_6_LC_11_22_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIE3BQ1_0_6_LC_11_22_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNIE3BQ1_0_6_LC_11_22_0  (
            .in0(N__28732),
            .in1(N__28552),
            .in2(N__28718),
            .in3(N__33274),
            .lcout(\pid_alt.m21_e_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIE3BQ1_6_LC_11_22_2 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIE3BQ1_6_LC_11_22_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIE3BQ1_6_LC_11_22_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNIE3BQ1_6_LC_11_22_2  (
            .in0(N__28733),
            .in1(N__28553),
            .in2(N__28719),
            .in3(N__33275),
            .lcout(\pid_alt.m35_e_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_8_LC_11_22_4 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_8_LC_11_22_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_8_LC_11_22_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_8_LC_11_22_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30422),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47265),
            .ce(N__33619),
            .sr(N__43889));
    defparam \pid_alt.error_i_acumm_prereg_esr_9_LC_11_22_5 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_9_LC_11_22_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_9_LC_11_22_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_9_LC_11_22_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30376),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47265),
            .ce(N__33619),
            .sr(N__43889));
    defparam \uart_pc.timer_Count_RNIVT8S_2_LC_12_6_0 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_RNIVT8S_2_LC_12_6_0 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNIVT8S_2_LC_12_6_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uart_pc.timer_Count_RNIVT8S_2_LC_12_6_0  (
            .in0(_gnd_net_),
            .in1(N__31605),
            .in2(_gnd_net_),
            .in3(N__27494),
            .lcout(\uart_pc.N_126_li ),
            .ltout(\uart_pc.N_126_li_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_RNIBLRB2_4_LC_12_6_1 .C_ON=1'b0;
    defparam \uart_pc.state_RNIBLRB2_4_LC_12_6_1 .SEQ_MODE=4'b0000;
    defparam \uart_pc.state_RNIBLRB2_4_LC_12_6_1 .LUT_INIT=16'b1101111111001100;
    LogicCell40 \uart_pc.state_RNIBLRB2_4_LC_12_6_1  (
            .in0(N__27477),
            .in1(N__31554),
            .in2(N__27471),
            .in3(N__31709),
            .lcout(\uart_pc.un1_state_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_RNIGRIF1_2_LC_12_6_4 .C_ON=1'b0;
    defparam \uart_pc.state_RNIGRIF1_2_LC_12_6_4 .SEQ_MODE=4'b0000;
    defparam \uart_pc.state_RNIGRIF1_2_LC_12_6_4 .LUT_INIT=16'b0011001011111010;
    LogicCell40 \uart_pc.state_RNIGRIF1_2_LC_12_6_4  (
            .in0(N__31710),
            .in1(N__31503),
            .in2(N__31113),
            .in3(N__31606),
            .lcout(\uart_pc.timer_Count_0_sqmuxa ),
            .ltout(\uart_pc.timer_Count_0_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_3_LC_12_6_5 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_3_LC_12_6_5 .SEQ_MODE=4'b1000;
    defparam \uart_pc.timer_Count_3_LC_12_6_5 .LUT_INIT=16'b0000000010101000;
    LogicCell40 \uart_pc.timer_Count_3_LC_12_6_5  (
            .in0(N__27444),
            .in1(N__27554),
            .in2(N__27438),
            .in3(N__44125),
            .lcout(\uart_pc.timer_CountZ1Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47412),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_4_LC_12_7_3 .C_ON=1'b0;
    defparam \uart_pc.state_4_LC_12_7_3 .SEQ_MODE=4'b1000;
    defparam \uart_pc.state_4_LC_12_7_3 .LUT_INIT=16'b1111111101000000;
    LogicCell40 \uart_pc.state_4_LC_12_7_3  (
            .in0(N__44102),
            .in1(N__31722),
            .in2(N__28539),
            .in3(N__27551),
            .lcout(\uart_pc.stateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47400),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_RNO_0_3_LC_12_7_5 .C_ON=1'b0;
    defparam \uart_pc.state_RNO_0_3_LC_12_7_5 .SEQ_MODE=4'b0000;
    defparam \uart_pc.state_RNO_0_3_LC_12_7_5 .LUT_INIT=16'b0000000001111111;
    LogicCell40 \uart_pc.state_RNO_0_3_LC_12_7_5  (
            .in0(N__31504),
            .in1(N__31611),
            .in2(N__31112),
            .in3(N__31721),
            .lcout(),
            .ltout(\uart_pc.N_145_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_3_LC_12_7_6 .C_ON=1'b0;
    defparam \uart_pc.state_3_LC_12_7_6 .SEQ_MODE=4'b1000;
    defparam \uart_pc.state_3_LC_12_7_6 .LUT_INIT=16'b0000000000001011;
    LogicCell40 \uart_pc.state_3_LC_12_7_6  (
            .in0(N__31108),
            .in1(N__28535),
            .in2(N__27522),
            .in3(N__44103),
            .lcout(\uart_pc.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47400),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_5_LC_12_8_0 .C_ON=1'b0;
    defparam \uart_pc.data_5_LC_12_8_0 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_5_LC_12_8_0 .LUT_INIT=16'b0011101000001010;
    LogicCell40 \uart_pc.data_5_LC_12_8_0  (
            .in0(N__33345),
            .in1(N__31068),
            .in2(N__31001),
            .in3(N__28781),
            .lcout(uart_pc_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47385),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_RNIEAGS_4_LC_12_8_1 .C_ON=1'b0;
    defparam \uart_pc.state_RNIEAGS_4_LC_12_8_1 .SEQ_MODE=4'b0000;
    defparam \uart_pc.state_RNIEAGS_4_LC_12_8_1 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \uart_pc.state_RNIEAGS_4_LC_12_8_1  (
            .in0(N__31711),
            .in1(N__31555),
            .in2(_gnd_net_),
            .in3(N__44089),
            .lcout(\uart_pc.state_RNIEAGSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_6_LC_12_8_5 .C_ON=1'b0;
    defparam \uart_pc.data_6_LC_12_8_5 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_6_LC_12_8_5 .LUT_INIT=16'b0101110100001000;
    LogicCell40 \uart_pc.data_6_LC_12_8_5  (
            .in0(N__30990),
            .in1(N__29123),
            .in2(N__31074),
            .in3(N__44946),
            .lcout(uart_pc_data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47385),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_2_LC_12_8_6 .C_ON=1'b0;
    defparam \uart_pc.data_2_LC_12_8_6 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_2_LC_12_8_6 .LUT_INIT=16'b0011000010101010;
    LogicCell40 \uart_pc.data_2_LC_12_8_6  (
            .in0(N__36819),
            .in1(N__31067),
            .in2(N__28842),
            .in3(N__30991),
            .lcout(uart_pc_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47385),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.data_Aux_RNO_0_4_LC_12_8_7 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_RNO_0_4_LC_12_8_7 .SEQ_MODE=4'b0000;
    defparam \uart_drone.data_Aux_RNO_0_4_LC_12_8_7 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \uart_drone.data_Aux_RNO_0_4_LC_12_8_7  (
            .in0(N__39518),
            .in1(N__36679),
            .in2(_gnd_net_),
            .in3(N__44420),
            .lcout(\uart_drone.data_Auxce_0_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.data_Aux_RNO_0_3_LC_12_9_1 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_RNO_0_3_LC_12_9_1 .SEQ_MODE=4'b0000;
    defparam \uart_drone.data_Aux_RNO_0_3_LC_12_9_1 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \uart_drone.data_Aux_RNO_0_3_LC_12_9_1  (
            .in0(N__44421),
            .in1(N__36687),
            .in2(_gnd_net_),
            .in3(N__39502),
            .lcout(\uart_drone.data_Auxce_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.data_Aux_RNO_0_5_LC_12_9_6 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_RNO_0_5_LC_12_9_6 .SEQ_MODE=4'b0000;
    defparam \uart_drone.data_Aux_RNO_0_5_LC_12_9_6 .LUT_INIT=16'b0101000000000000;
    LogicCell40 \uart_drone.data_Aux_RNO_0_5_LC_12_9_6  (
            .in0(N__39503),
            .in1(_gnd_net_),
            .in2(N__36693),
            .in3(N__44422),
            .lcout(\uart_drone.data_Auxce_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_1_4_LC_12_9_7 .C_ON=1'b0;
    defparam \uart_pc.data_1_4_LC_12_9_7 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_1_4_LC_12_9_7 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \uart_pc.data_1_4_LC_12_9_7  (
            .in0(N__31052),
            .in1(N__31000),
            .in2(N__28800),
            .in3(N__44205),
            .lcout(uart_pc_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47373),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_offset2data_esr_0_LC_12_10_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset2data_esr_0_LC_12_10_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset2data_esr_0_LC_12_10_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset2data_esr_0_LC_12_10_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27653),
            .lcout(frame_decoder_OFF2data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47360),
            .ce(N__27567),
            .sr(N__43818));
    defparam \Commands_frame_decoder.source_offset2data_esr_1_LC_12_10_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset2data_esr_1_LC_12_10_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset2data_esr_1_LC_12_10_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset2data_esr_1_LC_12_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45161),
            .lcout(frame_decoder_OFF2data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47360),
            .ce(N__27567),
            .sr(N__43818));
    defparam \Commands_frame_decoder.source_offset2data_esr_2_LC_12_10_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset2data_esr_2_LC_12_10_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset2data_esr_2_LC_12_10_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset2data_esr_2_LC_12_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36855),
            .lcout(frame_decoder_OFF2data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47360),
            .ce(N__27567),
            .sr(N__43818));
    defparam \Commands_frame_decoder.source_offset2data_esr_3_LC_12_10_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset2data_esr_3_LC_12_10_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset2data_esr_3_LC_12_10_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset2data_esr_3_LC_12_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43308),
            .lcout(frame_decoder_OFF2data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47360),
            .ce(N__27567),
            .sr(N__43818));
    defparam \Commands_frame_decoder.source_offset2data_esr_4_LC_12_10_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset2data_esr_4_LC_12_10_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset2data_esr_4_LC_12_10_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset2data_esr_4_LC_12_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45298),
            .lcout(frame_decoder_OFF2data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47360),
            .ce(N__27567),
            .sr(N__43818));
    defparam \Commands_frame_decoder.source_offset2data_esr_5_LC_12_10_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset2data_esr_5_LC_12_10_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset2data_esr_5_LC_12_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset2data_esr_5_LC_12_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44206),
            .lcout(frame_decoder_OFF2data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47360),
            .ce(N__27567),
            .sr(N__43818));
    defparam \Commands_frame_decoder.source_offset2data_esr_6_LC_12_10_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset2data_esr_6_LC_12_10_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset2data_esr_6_LC_12_10_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Commands_frame_decoder.source_offset2data_esr_6_LC_12_10_6  (
            .in0(N__33362),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(frame_decoder_OFF2data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47360),
            .ce(N__27567),
            .sr(N__43818));
    defparam \Commands_frame_decoder.source_offset2data_ess_7_LC_12_10_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset2data_ess_7_LC_12_10_7 .SEQ_MODE=4'b1001;
    defparam \Commands_frame_decoder.source_offset2data_ess_7_LC_12_10_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset2data_ess_7_LC_12_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44953),
            .lcout(frame_decoder_OFF2data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47360),
            .ce(N__27567),
            .sr(N__43818));
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_0_c_LC_12_11_0 .C_ON=1'b1;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_0_c_LC_12_11_0 .SEQ_MODE=4'b0000;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_0_c_LC_12_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \scaler_2.un3_source_data_un3_source_data_0_cry_0_c_LC_12_11_0  (
            .in0(_gnd_net_),
            .in1(N__29035),
            .in2(N__29081),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_11_0_),
            .carryout(\scaler_2.un3_source_data_0_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_0_c_RNIUVGK_LC_12_11_1 .C_ON=1'b1;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_0_c_RNIUVGK_LC_12_11_1 .SEQ_MODE=4'b0000;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_0_c_RNIUVGK_LC_12_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_2.un3_source_data_un3_source_data_0_cry_0_c_RNIUVGK_LC_12_11_1  (
            .in0(_gnd_net_),
            .in1(N__27810),
            .in2(N__27804),
            .in3(N__27795),
            .lcout(\scaler_2.un2_source_data_0 ),
            .ltout(),
            .carryin(\scaler_2.un3_source_data_0_cry_0 ),
            .carryout(\scaler_2.un3_source_data_0_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_1_c_RNI14IK_LC_12_11_2 .C_ON=1'b1;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_1_c_RNI14IK_LC_12_11_2 .SEQ_MODE=4'b0000;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_1_c_RNI14IK_LC_12_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_2.un3_source_data_un3_source_data_0_cry_1_c_RNI14IK_LC_12_11_2  (
            .in0(_gnd_net_),
            .in1(N__27792),
            .in2(N__27786),
            .in3(N__27777),
            .lcout(\scaler_2.un3_source_data_0_cry_1_c_RNI14IK ),
            .ltout(),
            .carryin(\scaler_2.un3_source_data_0_cry_1 ),
            .carryout(\scaler_2.un3_source_data_0_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_2_c_RNI48JK_LC_12_11_3 .C_ON=1'b1;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_2_c_RNI48JK_LC_12_11_3 .SEQ_MODE=4'b0000;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_2_c_RNI48JK_LC_12_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_2.un3_source_data_un3_source_data_0_cry_2_c_RNI48JK_LC_12_11_3  (
            .in0(_gnd_net_),
            .in1(N__27774),
            .in2(N__27768),
            .in3(N__27759),
            .lcout(\scaler_2.un3_source_data_0_cry_2_c_RNI48JK ),
            .ltout(),
            .carryin(\scaler_2.un3_source_data_0_cry_2 ),
            .carryout(\scaler_2.un3_source_data_0_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_3_c_RNI7CKK_LC_12_11_4 .C_ON=1'b1;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_3_c_RNI7CKK_LC_12_11_4 .SEQ_MODE=4'b0000;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_3_c_RNI7CKK_LC_12_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_2.un3_source_data_un3_source_data_0_cry_3_c_RNI7CKK_LC_12_11_4  (
            .in0(_gnd_net_),
            .in1(N__27756),
            .in2(N__27750),
            .in3(N__27741),
            .lcout(\scaler_2.un3_source_data_0_cry_3_c_RNI7CKK ),
            .ltout(),
            .carryin(\scaler_2.un3_source_data_0_cry_3 ),
            .carryout(\scaler_2.un3_source_data_0_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_4_c_RNIAGLK_LC_12_11_5 .C_ON=1'b1;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_4_c_RNIAGLK_LC_12_11_5 .SEQ_MODE=4'b0000;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_4_c_RNIAGLK_LC_12_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_2.un3_source_data_un3_source_data_0_cry_4_c_RNIAGLK_LC_12_11_5  (
            .in0(_gnd_net_),
            .in1(N__27738),
            .in2(N__27732),
            .in3(N__27723),
            .lcout(\scaler_2.un3_source_data_0_cry_4_c_RNIAGLK ),
            .ltout(),
            .carryin(\scaler_2.un3_source_data_0_cry_4 ),
            .carryout(\scaler_2.un3_source_data_0_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_5_c_RNIDKMK_LC_12_11_6 .C_ON=1'b1;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_5_c_RNIDKMK_LC_12_11_6 .SEQ_MODE=4'b0000;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_5_c_RNIDKMK_LC_12_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_2.un3_source_data_un3_source_data_0_cry_5_c_RNIDKMK_LC_12_11_6  (
            .in0(_gnd_net_),
            .in1(N__27720),
            .in2(N__27714),
            .in3(N__27705),
            .lcout(\scaler_2.un3_source_data_0_cry_5_c_RNIDKMK ),
            .ltout(),
            .carryin(\scaler_2.un3_source_data_0_cry_5 ),
            .carryout(\scaler_2.un3_source_data_0_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_6_c_RNIIUTM_LC_12_11_7 .C_ON=1'b1;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_6_c_RNIIUTM_LC_12_11_7 .SEQ_MODE=4'b0000;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_6_c_RNIIUTM_LC_12_11_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \scaler_2.un3_source_data_un3_source_data_0_cry_6_c_RNIIUTM_LC_12_11_7  (
            .in0(_gnd_net_),
            .in1(N__27702),
            .in2(_gnd_net_),
            .in3(N__27696),
            .lcout(\scaler_2.un3_source_data_0_cry_6_c_RNIIUTM ),
            .ltout(),
            .carryin(\scaler_2.un3_source_data_0_cry_6 ),
            .carryout(\scaler_2.un3_source_data_0_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_7_c_RNIJ0VM_LC_12_12_0 .C_ON=1'b1;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_7_c_RNIJ0VM_LC_12_12_0 .SEQ_MODE=4'b0000;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_7_c_RNIJ0VM_LC_12_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_2.un3_source_data_un3_source_data_0_cry_7_c_RNIJ0VM_LC_12_12_0  (
            .in0(_gnd_net_),
            .in1(N__28080),
            .in2(N__43123),
            .in3(N__28113),
            .lcout(\scaler_2.un3_source_data_0_cry_7_c_RNIJ0VM ),
            .ltout(),
            .carryin(bfn_12_12_0_),
            .carryout(\scaler_2.un3_source_data_0_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_8_c_RNIQL42_LC_12_12_1 .C_ON=1'b0;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_8_c_RNIQL42_LC_12_12_1 .SEQ_MODE=4'b0000;
    defparam \scaler_2.un3_source_data_un3_source_data_0_cry_8_c_RNIQL42_LC_12_12_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \scaler_2.un3_source_data_un3_source_data_0_cry_8_c_RNIQL42_LC_12_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28110),
            .lcout(\scaler_2.un3_source_data_0_cry_8_c_RNIQL42 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI7O1N_2_LC_12_12_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI7O1N_2_LC_12_12_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI7O1N_2_LC_12_12_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI7O1N_2_LC_12_12_2  (
            .in0(_gnd_net_),
            .in1(N__42274),
            .in2(_gnd_net_),
            .in3(N__42010),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI7O1NZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_2.N_1227_i_l_ofx_LC_12_12_7 .C_ON=1'b0;
    defparam \scaler_2.N_1227_i_l_ofx_LC_12_12_7 .SEQ_MODE=4'b0000;
    defparam \scaler_2.N_1227_i_l_ofx_LC_12_12_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \scaler_2.N_1227_i_l_ofx_LC_12_12_7  (
            .in0(_gnd_net_),
            .in1(N__28107),
            .in2(_gnd_net_),
            .in3(N__28092),
            .lcout(\scaler_2.N_1227_i_l_ofxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.source_pid_1_esr_9_LC_12_13_0 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_esr_9_LC_12_13_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_esr_9_LC_12_13_0 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \pid_alt.source_pid_1_esr_9_LC_12_13_0  (
            .in0(N__28066),
            .in1(N__27987),
            .in2(_gnd_net_),
            .in3(N__27951),
            .lcout(throttle_command_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47316),
            .ce(N__27918),
            .sr(N__27876));
    defparam \scaler_2.un2_source_data_0_cry_1_c_RNO_LC_12_13_2 .C_ON=1'b0;
    defparam \scaler_2.un2_source_data_0_cry_1_c_RNO_LC_12_13_2 .SEQ_MODE=4'b0000;
    defparam \scaler_2.un2_source_data_0_cry_1_c_RNO_LC_12_13_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \scaler_2.un2_source_data_0_cry_1_c_RNO_LC_12_13_2  (
            .in0(N__32284),
            .in1(N__29044),
            .in2(_gnd_net_),
            .in3(N__29082),
            .lcout(\scaler_2.un2_source_data_0_cry_1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un2_source_data_0_cry_1_c_RNO_LC_12_13_4 .C_ON=1'b0;
    defparam \scaler_4.un2_source_data_0_cry_1_c_RNO_LC_12_13_4 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un2_source_data_0_cry_1_c_RNO_LC_12_13_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \scaler_4.un2_source_data_0_cry_1_c_RNO_LC_12_13_4  (
            .in0(N__28913),
            .in1(N__29551),
            .in2(_gnd_net_),
            .in3(N__29512),
            .lcout(\scaler_4.un2_source_data_0_cry_1_c_RNO_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_3.un2_source_data_0_cry_1_c_LC_12_14_0 .C_ON=1'b1;
    defparam \scaler_3.un2_source_data_0_cry_1_c_LC_12_14_0 .SEQ_MODE=4'b0000;
    defparam \scaler_3.un2_source_data_0_cry_1_c_LC_12_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \scaler_3.un2_source_data_0_cry_1_c_LC_12_14_0  (
            .in0(_gnd_net_),
            .in1(N__29007),
            .in2(N__27825),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_14_0_),
            .carryout(\scaler_3.un2_source_data_0_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_3.source_data_1_esr_6_LC_12_14_1 .C_ON=1'b1;
    defparam \scaler_3.source_data_1_esr_6_LC_12_14_1 .SEQ_MODE=4'b1000;
    defparam \scaler_3.source_data_1_esr_6_LC_12_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_3.source_data_1_esr_6_LC_12_14_1  (
            .in0(_gnd_net_),
            .in1(N__28226),
            .in2(N__29015),
            .in3(N__27813),
            .lcout(scaler_3_data_6),
            .ltout(),
            .carryin(\scaler_3.un2_source_data_0_cry_1 ),
            .carryout(\scaler_3.un2_source_data_0_cry_2 ),
            .clk(N__47305),
            .ce(N__32403),
            .sr(N__43847));
    defparam \scaler_3.source_data_1_esr_7_LC_12_14_2 .C_ON=1'b1;
    defparam \scaler_3.source_data_1_esr_7_LC_12_14_2 .SEQ_MODE=4'b1000;
    defparam \scaler_3.source_data_1_esr_7_LC_12_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_3.source_data_1_esr_7_LC_12_14_2  (
            .in0(_gnd_net_),
            .in1(N__28211),
            .in2(N__28230),
            .in3(N__28218),
            .lcout(scaler_3_data_7),
            .ltout(),
            .carryin(\scaler_3.un2_source_data_0_cry_2 ),
            .carryout(\scaler_3.un2_source_data_0_cry_3 ),
            .clk(N__47305),
            .ce(N__32403),
            .sr(N__43847));
    defparam \scaler_3.source_data_1_esr_8_LC_12_14_3 .C_ON=1'b1;
    defparam \scaler_3.source_data_1_esr_8_LC_12_14_3 .SEQ_MODE=4'b1000;
    defparam \scaler_3.source_data_1_esr_8_LC_12_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_3.source_data_1_esr_8_LC_12_14_3  (
            .in0(_gnd_net_),
            .in1(N__28196),
            .in2(N__28215),
            .in3(N__28203),
            .lcout(scaler_3_data_8),
            .ltout(),
            .carryin(\scaler_3.un2_source_data_0_cry_3 ),
            .carryout(\scaler_3.un2_source_data_0_cry_4 ),
            .clk(N__47305),
            .ce(N__32403),
            .sr(N__43847));
    defparam \scaler_3.source_data_1_esr_9_LC_12_14_4 .C_ON=1'b1;
    defparam \scaler_3.source_data_1_esr_9_LC_12_14_4 .SEQ_MODE=4'b1000;
    defparam \scaler_3.source_data_1_esr_9_LC_12_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_3.source_data_1_esr_9_LC_12_14_4  (
            .in0(_gnd_net_),
            .in1(N__28181),
            .in2(N__28200),
            .in3(N__28188),
            .lcout(scaler_3_data_9),
            .ltout(),
            .carryin(\scaler_3.un2_source_data_0_cry_4 ),
            .carryout(\scaler_3.un2_source_data_0_cry_5 ),
            .clk(N__47305),
            .ce(N__32403),
            .sr(N__43847));
    defparam \scaler_3.source_data_1_esr_10_LC_12_14_5 .C_ON=1'b1;
    defparam \scaler_3.source_data_1_esr_10_LC_12_14_5 .SEQ_MODE=4'b1000;
    defparam \scaler_3.source_data_1_esr_10_LC_12_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_3.source_data_1_esr_10_LC_12_14_5  (
            .in0(_gnd_net_),
            .in1(N__28166),
            .in2(N__28185),
            .in3(N__28173),
            .lcout(scaler_3_data_10),
            .ltout(),
            .carryin(\scaler_3.un2_source_data_0_cry_5 ),
            .carryout(\scaler_3.un2_source_data_0_cry_6 ),
            .clk(N__47305),
            .ce(N__32403),
            .sr(N__43847));
    defparam \scaler_3.source_data_1_esr_11_LC_12_14_6 .C_ON=1'b1;
    defparam \scaler_3.source_data_1_esr_11_LC_12_14_6 .SEQ_MODE=4'b1000;
    defparam \scaler_3.source_data_1_esr_11_LC_12_14_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_3.source_data_1_esr_11_LC_12_14_6  (
            .in0(_gnd_net_),
            .in1(N__28151),
            .in2(N__28170),
            .in3(N__28158),
            .lcout(scaler_3_data_11),
            .ltout(),
            .carryin(\scaler_3.un2_source_data_0_cry_6 ),
            .carryout(\scaler_3.un2_source_data_0_cry_7 ),
            .clk(N__47305),
            .ce(N__32403),
            .sr(N__43847));
    defparam \scaler_3.source_data_1_esr_12_LC_12_14_7 .C_ON=1'b1;
    defparam \scaler_3.source_data_1_esr_12_LC_12_14_7 .SEQ_MODE=4'b1000;
    defparam \scaler_3.source_data_1_esr_12_LC_12_14_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_3.source_data_1_esr_12_LC_12_14_7  (
            .in0(_gnd_net_),
            .in1(N__28139),
            .in2(N__28155),
            .in3(N__28143),
            .lcout(scaler_3_data_12),
            .ltout(),
            .carryin(\scaler_3.un2_source_data_0_cry_7 ),
            .carryout(\scaler_3.un2_source_data_0_cry_8 ),
            .clk(N__47305),
            .ce(N__32403),
            .sr(N__43847));
    defparam \scaler_3.source_data_1_esr_13_LC_12_15_0 .C_ON=1'b1;
    defparam \scaler_3.source_data_1_esr_13_LC_12_15_0 .SEQ_MODE=4'b1000;
    defparam \scaler_3.source_data_1_esr_13_LC_12_15_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_3.source_data_1_esr_13_LC_12_15_0  (
            .in0(_gnd_net_),
            .in1(N__28140),
            .in2(N__28128),
            .in3(N__28119),
            .lcout(scaler_3_data_13),
            .ltout(),
            .carryin(bfn_12_15_0_),
            .carryout(\scaler_3.un2_source_data_0_cry_9 ),
            .clk(N__47297),
            .ce(N__32402),
            .sr(N__43852));
    defparam \scaler_3.source_data_1_esr_14_LC_12_15_1 .C_ON=1'b0;
    defparam \scaler_3.source_data_1_esr_14_LC_12_15_1 .SEQ_MODE=4'b1000;
    defparam \scaler_3.source_data_1_esr_14_LC_12_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \scaler_3.source_data_1_esr_14_LC_12_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28116),
            .lcout(scaler_3_data_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47297),
            .ce(N__32402),
            .sr(N__43852));
    defparam \scaler_4.un2_source_data_0_cry_1_c_LC_12_16_0 .C_ON=1'b1;
    defparam \scaler_4.un2_source_data_0_cry_1_c_LC_12_16_0 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un2_source_data_0_cry_1_c_LC_12_16_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \scaler_4.un2_source_data_0_cry_1_c_LC_12_16_0  (
            .in0(_gnd_net_),
            .in1(N__28899),
            .in2(N__28359),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_16_0_),
            .carryout(\scaler_4.un2_source_data_0_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.source_data_1_esr_6_LC_12_16_1 .C_ON=1'b1;
    defparam \scaler_4.source_data_1_esr_6_LC_12_16_1 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_6_LC_12_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.source_data_1_esr_6_LC_12_16_1  (
            .in0(_gnd_net_),
            .in1(N__28340),
            .in2(N__28909),
            .in3(N__28347),
            .lcout(scaler_4_data_6),
            .ltout(),
            .carryin(\scaler_4.un2_source_data_0_cry_1 ),
            .carryout(\scaler_4.un2_source_data_0_cry_2 ),
            .clk(N__47290),
            .ce(N__32401),
            .sr(N__43858));
    defparam \scaler_4.source_data_1_esr_7_LC_12_16_2 .C_ON=1'b1;
    defparam \scaler_4.source_data_1_esr_7_LC_12_16_2 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_7_LC_12_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.source_data_1_esr_7_LC_12_16_2  (
            .in0(_gnd_net_),
            .in1(N__28325),
            .in2(N__28344),
            .in3(N__28332),
            .lcout(scaler_4_data_7),
            .ltout(),
            .carryin(\scaler_4.un2_source_data_0_cry_2 ),
            .carryout(\scaler_4.un2_source_data_0_cry_3 ),
            .clk(N__47290),
            .ce(N__32401),
            .sr(N__43858));
    defparam \scaler_4.source_data_1_esr_8_LC_12_16_3 .C_ON=1'b1;
    defparam \scaler_4.source_data_1_esr_8_LC_12_16_3 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_8_LC_12_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.source_data_1_esr_8_LC_12_16_3  (
            .in0(_gnd_net_),
            .in1(N__28310),
            .in2(N__28329),
            .in3(N__28317),
            .lcout(scaler_4_data_8),
            .ltout(),
            .carryin(\scaler_4.un2_source_data_0_cry_3 ),
            .carryout(\scaler_4.un2_source_data_0_cry_4 ),
            .clk(N__47290),
            .ce(N__32401),
            .sr(N__43858));
    defparam \scaler_4.source_data_1_esr_9_LC_12_16_4 .C_ON=1'b1;
    defparam \scaler_4.source_data_1_esr_9_LC_12_16_4 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_9_LC_12_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.source_data_1_esr_9_LC_12_16_4  (
            .in0(_gnd_net_),
            .in1(N__28295),
            .in2(N__28314),
            .in3(N__28302),
            .lcout(scaler_4_data_9),
            .ltout(),
            .carryin(\scaler_4.un2_source_data_0_cry_4 ),
            .carryout(\scaler_4.un2_source_data_0_cry_5 ),
            .clk(N__47290),
            .ce(N__32401),
            .sr(N__43858));
    defparam \scaler_4.source_data_1_esr_10_LC_12_16_5 .C_ON=1'b1;
    defparam \scaler_4.source_data_1_esr_10_LC_12_16_5 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_10_LC_12_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.source_data_1_esr_10_LC_12_16_5  (
            .in0(_gnd_net_),
            .in1(N__28280),
            .in2(N__28299),
            .in3(N__28287),
            .lcout(scaler_4_data_10),
            .ltout(),
            .carryin(\scaler_4.un2_source_data_0_cry_5 ),
            .carryout(\scaler_4.un2_source_data_0_cry_6 ),
            .clk(N__47290),
            .ce(N__32401),
            .sr(N__43858));
    defparam \scaler_4.source_data_1_esr_11_LC_12_16_6 .C_ON=1'b1;
    defparam \scaler_4.source_data_1_esr_11_LC_12_16_6 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_11_LC_12_16_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.source_data_1_esr_11_LC_12_16_6  (
            .in0(_gnd_net_),
            .in1(N__28265),
            .in2(N__28284),
            .in3(N__28272),
            .lcout(scaler_4_data_11),
            .ltout(),
            .carryin(\scaler_4.un2_source_data_0_cry_6 ),
            .carryout(\scaler_4.un2_source_data_0_cry_7 ),
            .clk(N__47290),
            .ce(N__32401),
            .sr(N__43858));
    defparam \scaler_4.source_data_1_esr_12_LC_12_16_7 .C_ON=1'b1;
    defparam \scaler_4.source_data_1_esr_12_LC_12_16_7 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_12_LC_12_16_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.source_data_1_esr_12_LC_12_16_7  (
            .in0(_gnd_net_),
            .in1(N__28253),
            .in2(N__28269),
            .in3(N__28257),
            .lcout(scaler_4_data_12),
            .ltout(),
            .carryin(\scaler_4.un2_source_data_0_cry_7 ),
            .carryout(\scaler_4.un2_source_data_0_cry_8 ),
            .clk(N__47290),
            .ce(N__32401),
            .sr(N__43858));
    defparam \scaler_4.source_data_1_esr_13_LC_12_17_0 .C_ON=1'b1;
    defparam \scaler_4.source_data_1_esr_13_LC_12_17_0 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_13_LC_12_17_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.source_data_1_esr_13_LC_12_17_0  (
            .in0(_gnd_net_),
            .in1(N__28254),
            .in2(N__28242),
            .in3(N__28233),
            .lcout(scaler_4_data_13),
            .ltout(),
            .carryin(bfn_12_17_0_),
            .carryout(\scaler_4.un2_source_data_0_cry_9 ),
            .clk(N__47282),
            .ce(N__32400),
            .sr(N__43867));
    defparam \scaler_4.source_data_1_esr_14_LC_12_17_1 .C_ON=1'b0;
    defparam \scaler_4.source_data_1_esr_14_LC_12_17_1 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_14_LC_12_17_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \scaler_4.source_data_1_esr_14_LC_12_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28365),
            .lcout(scaler_4_data_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47282),
            .ce(N__32400),
            .sr(N__43867));
    defparam \ppm_encoder_1.init_pulses_RNI0KRP_0_17_LC_12_18_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI0KRP_0_17_LC_12_18_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI0KRP_0_17_LC_12_18_7 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI0KRP_0_17_LC_12_18_7  (
            .in0(N__41922),
            .in1(N__40755),
            .in2(_gnd_net_),
            .in3(N__42275),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_axb_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIHB5T_5_LC_12_19_3 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIHB5T_5_LC_12_19_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIHB5T_5_LC_12_19_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNIHB5T_5_LC_12_19_3  (
            .in0(_gnd_net_),
            .in1(N__28626),
            .in2(_gnd_net_),
            .in3(N__28507),
            .lcout(\pid_alt.m21_e_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.state_RNIAAPN5_1_LC_12_19_5 .C_ON=1'b0;
    defparam \pid_alt.state_RNIAAPN5_1_LC_12_19_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.state_RNIAAPN5_1_LC_12_19_5 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \pid_alt.state_RNIAAPN5_1_LC_12_19_5  (
            .in0(N__33208),
            .in1(N__32942),
            .in2(_gnd_net_),
            .in3(N__28425),
            .lcout(\pid_alt.un1_reset_1_0_i ),
            .ltout(\pid_alt.un1_reset_1_0_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.state_RNIVV066_1_LC_12_19_6 .C_ON=1'b0;
    defparam \pid_alt.state_RNIVV066_1_LC_12_19_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.state_RNIVV066_1_LC_12_19_6 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \pid_alt.state_RNIVV066_1_LC_12_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__28362),
            .in3(N__33209),
            .lcout(\pid_alt.N_96_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_esr_0_LC_12_20_0 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_esr_0_LC_12_20_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_esr_0_LC_12_20_0 .LUT_INIT=16'b1100010010000000;
    LogicCell40 \pid_alt.error_i_acumm_esr_0_LC_12_20_0  (
            .in0(N__28520),
            .in1(N__33654),
            .in2(N__28672),
            .in3(N__28401),
            .lcout(\pid_alt.error_i_acummZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47267),
            .ce(N__32771),
            .sr(N__33693));
    defparam \pid_alt.error_i_acumm_esr_1_LC_12_20_2 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_esr_1_LC_12_20_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_esr_1_LC_12_20_2 .LUT_INIT=16'b1100010010000000;
    LogicCell40 \pid_alt.error_i_acumm_esr_1_LC_12_20_2  (
            .in0(N__28521),
            .in1(N__28388),
            .in2(N__28673),
            .in3(N__28402),
            .lcout(\pid_alt.error_i_acummZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47267),
            .ce(N__32771),
            .sr(N__33693));
    defparam \pid_alt.error_i_acumm_esr_2_LC_12_20_3 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_esr_2_LC_12_20_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_esr_2_LC_12_20_3 .LUT_INIT=16'b1100101000000000;
    LogicCell40 \pid_alt.error_i_acumm_esr_2_LC_12_20_3  (
            .in0(N__28403),
            .in1(N__28667),
            .in2(N__28527),
            .in3(N__28487),
            .lcout(\pid_alt.error_i_acummZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47267),
            .ce(N__32771),
            .sr(N__33693));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIAP1A_13_LC_12_20_4 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIAP1A_13_LC_12_20_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIAP1A_13_LC_12_20_4 .LUT_INIT=16'b1010101011101110;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNIAP1A_13_LC_12_20_4  (
            .in0(N__32844),
            .in1(N__32795),
            .in2(_gnd_net_),
            .in3(N__32821),
            .lcout(\pid_alt.N_9_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_esr_4_LC_12_20_6 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_esr_4_LC_12_20_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_esr_4_LC_12_20_6 .LUT_INIT=16'b1010111010111111;
    LogicCell40 \pid_alt.error_i_acumm_esr_4_LC_12_20_6  (
            .in0(N__28522),
            .in1(N__28637),
            .in2(N__28674),
            .in3(N__33076),
            .lcout(\pid_alt.error_i_acummZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47267),
            .ce(N__32771),
            .sr(N__33693));
    defparam \pid_alt.error_i_acumm_esr_3_LC_12_20_7 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_esr_3_LC_12_20_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_esr_3_LC_12_20_7 .LUT_INIT=16'b1100000010100000;
    LogicCell40 \pid_alt.error_i_acumm_esr_3_LC_12_20_7  (
            .in0(N__28404),
            .in1(N__28668),
            .in2(N__28467),
            .in3(N__28523),
            .lcout(\pid_alt.error_i_acummZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47267),
            .ce(N__32771),
            .sr(N__33693));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNICMLK3_2_LC_12_21_0 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNICMLK3_2_LC_12_21_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNICMLK3_2_LC_12_21_0 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNICMLK3_2_LC_12_21_0  (
            .in0(N__28488),
            .in1(N__28473),
            .in2(N__28466),
            .in3(N__28437),
            .lcout(),
            .ltout(\pid_alt.m21_e_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIO7B05_21_LC_12_21_1 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIO7B05_21_LC_12_21_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIO7B05_21_LC_12_21_1 .LUT_INIT=16'b1110101000101010;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNIO7B05_21_LC_12_21_1  (
            .in0(N__32852),
            .in1(N__28371),
            .in2(N__28428),
            .in3(N__28573),
            .lcout(\pid_alt.N_138 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI4SOH2_10_LC_12_21_2 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI4SOH2_10_LC_12_21_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI4SOH2_10_LC_12_21_2 .LUT_INIT=16'b1011111110000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNI4SOH2_10_LC_12_21_2  (
            .in0(N__28574),
            .in1(N__28416),
            .in2(N__28683),
            .in3(N__33049),
            .lcout(\pid_alt.N_62_mux ),
            .ltout(\pid_alt.N_62_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIEPGB3_5_LC_12_21_3 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIEPGB3_5_LC_12_21_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIEPGB3_5_LC_12_21_3 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNIEPGB3_5_LC_12_21_3  (
            .in0(N__33050),
            .in1(_gnd_net_),
            .in2(N__28407),
            .in3(N__28636),
            .lcout(\pid_alt.N_129 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI935T_0_LC_12_21_5 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI935T_0_LC_12_21_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI935T_0_LC_12_21_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNI935T_0_LC_12_21_5  (
            .in0(_gnd_net_),
            .in1(N__28389),
            .in2(_gnd_net_),
            .in3(N__33653),
            .lcout(),
            .ltout(\pid_alt.m21_e_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIB9F01_10_LC_12_21_6 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIB9F01_10_LC_12_21_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIB9F01_10_LC_12_21_6 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNIB9F01_10_LC_12_21_6  (
            .in0(N__33097),
            .in1(N__28696),
            .in2(N__28374),
            .in3(N__28594),
            .lcout(\pid_alt.m21_e_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_10_LC_12_22_0 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_10_LC_12_22_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_10_LC_12_22_0 .LUT_INIT=16'b1101100011111010;
    LogicCell40 \pid_alt.error_i_acumm_10_LC_12_22_0  (
            .in0(N__33230),
            .in1(N__28698),
            .in2(N__30354),
            .in3(N__33067),
            .lcout(\pid_alt.error_i_acummZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47264),
            .ce(),
            .sr(N__33703));
    defparam \pid_alt.error_i_acumm_8_LC_12_22_4 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_8_LC_12_22_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_8_LC_12_22_4 .LUT_INIT=16'b1100101011111010;
    LogicCell40 \pid_alt.error_i_acumm_8_LC_12_22_4  (
            .in0(N__30444),
            .in1(N__28734),
            .in2(N__33244),
            .in3(N__33068),
            .lcout(\pid_alt.error_i_acummZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47264),
            .ce(),
            .sr(N__33703));
    defparam \pid_alt.error_i_acumm_9_LC_12_22_5 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_9_LC_12_22_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_9_LC_12_22_5 .LUT_INIT=16'b1111110001110100;
    LogicCell40 \pid_alt.error_i_acumm_9_LC_12_22_5  (
            .in0(N__33069),
            .in1(N__33235),
            .in2(N__30399),
            .in3(N__28717),
            .lcout(\pid_alt.error_i_acummZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47264),
            .ce(),
            .sr(N__33703));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIBO62_10_LC_12_22_6 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIBO62_10_LC_12_22_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIBO62_10_LC_12_22_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNIBO62_10_LC_12_22_6  (
            .in0(N__33098),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28697),
            .lcout(\pid_alt.m35_e_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_5_LC_12_22_7 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_5_LC_12_22_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_5_LC_12_22_7 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \pid_alt.error_i_acumm_5_LC_12_22_7  (
            .in0(N__28660),
            .in1(N__29924),
            .in2(N__28641),
            .in3(N__33231),
            .lcout(\pid_alt.error_i_acummZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47264),
            .ce(),
            .sr(N__33703));
    defparam \pid_alt.error_i_acumm_12_LC_12_23_1 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_12_LC_12_23_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_12_LC_12_23_1 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \pid_alt.error_i_acumm_12_LC_12_23_1  (
            .in0(N__33236),
            .in1(N__30267),
            .in2(N__28602),
            .in3(N__28578),
            .lcout(\pid_alt.error_i_acummZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47263),
            .ce(),
            .sr(N__33718));
    defparam \pid_alt.error_i_acumm_7_LC_12_23_7 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_7_LC_12_23_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_7_LC_12_23_7 .LUT_INIT=16'b1111101000111010;
    LogicCell40 \pid_alt.error_i_acumm_7_LC_12_23_7  (
            .in0(N__30494),
            .in1(N__33070),
            .in2(N__33245),
            .in3(N__28560),
            .lcout(\pid_alt.error_i_acummZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47263),
            .ce(),
            .sr(N__33718));
    defparam \uart_drone.state_RNO_0_0_LC_13_6_6 .C_ON=1'b0;
    defparam \uart_drone.state_RNO_0_0_LC_13_6_6 .SEQ_MODE=4'b0000;
    defparam \uart_drone.state_RNO_0_0_LC_13_6_6 .LUT_INIT=16'b0000000011011101;
    LogicCell40 \uart_drone.state_RNO_0_0_LC_13_6_6  (
            .in0(N__31658),
            .in1(N__31372),
            .in2(_gnd_net_),
            .in3(N__44090),
            .lcout(\uart_drone.state_srsts_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNI5UFA2_3_LC_13_7_2 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_RNI5UFA2_3_LC_13_7_2 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNI5UFA2_3_LC_13_7_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uart_pc.timer_Count_RNI5UFA2_3_LC_13_7_2  (
            .in0(N__31509),
            .in1(N__31773),
            .in2(_gnd_net_),
            .in3(N__31607),
            .lcout(\uart_pc.N_144_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_1_LC_13_7_3 .C_ON=1'b0;
    defparam \uart_pc.data_1_LC_13_7_3 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_1_LC_13_7_3 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \uart_pc.data_1_LC_13_7_3  (
            .in0(N__30999),
            .in1(N__31072),
            .in2(N__28857),
            .in3(N__45130),
            .lcout(uart_pc_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47414),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNO_0_1_LC_13_7_6 .C_ON=1'b0;
    defparam \reset_module_System.count_RNO_0_1_LC_13_7_6 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNO_0_1_LC_13_7_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \reset_module_System.count_RNO_0_1_LC_13_7_6  (
            .in0(_gnd_net_),
            .in1(N__34832),
            .in2(_gnd_net_),
            .in3(N__34853),
            .lcout(),
            .ltout(\reset_module_System.count_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_1_LC_13_7_7 .C_ON=1'b0;
    defparam \reset_module_System.count_1_LC_13_7_7 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_1_LC_13_7_7 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \reset_module_System.count_1_LC_13_7_7  (
            .in0(N__33842),
            .in1(N__37318),
            .in2(N__28881),
            .in3(N__33792),
            .lcout(\reset_module_System.countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47414),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_Aux_0_LC_13_8_0 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_0_LC_13_8_0 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_Aux_0_LC_13_8_0 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \uart_pc.data_Aux_0_LC_13_8_0  (
            .in0(N__29214),
            .in1(N__31220),
            .in2(N__28874),
            .in3(N__28760),
            .lcout(\uart_pc.data_AuxZ1Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47403),
            .ce(),
            .sr(N__29109));
    defparam \uart_pc.data_Aux_1_LC_13_8_1 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_1_LC_13_8_1 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_Aux_1_LC_13_8_1 .LUT_INIT=16'b1101110010001100;
    LogicCell40 \uart_pc.data_Aux_1_LC_13_8_1  (
            .in0(N__28761),
            .in1(N__28853),
            .in2(N__29205),
            .in3(N__31224),
            .lcout(\uart_pc.data_AuxZ1Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47403),
            .ce(),
            .sr(N__29109));
    defparam \uart_pc.data_Aux_2_LC_13_8_2 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_2_LC_13_8_2 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_Aux_2_LC_13_8_2 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \uart_pc.data_Aux_2_LC_13_8_2  (
            .in0(N__29094),
            .in1(N__31221),
            .in2(N__28841),
            .in3(N__28762),
            .lcout(\uart_pc.data_AuxZ1Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47403),
            .ce(),
            .sr(N__29109));
    defparam \uart_pc.data_Aux_3_LC_13_8_3 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_3_LC_13_8_3 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_Aux_3_LC_13_8_3 .LUT_INIT=16'b1111010010110000;
    LogicCell40 \uart_pc.data_Aux_3_LC_13_8_3  (
            .in0(N__28763),
            .in1(N__29100),
            .in2(N__31019),
            .in3(N__31225),
            .lcout(\uart_pc.data_AuxZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47403),
            .ce(),
            .sr(N__29109));
    defparam \uart_pc.data_Aux_4_LC_13_8_4 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_4_LC_13_8_4 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_Aux_4_LC_13_8_4 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \uart_pc.data_Aux_4_LC_13_8_4  (
            .in0(N__29193),
            .in1(N__31222),
            .in2(N__28817),
            .in3(N__28764),
            .lcout(\uart_pc.data_AuxZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47403),
            .ce(),
            .sr(N__29109));
    defparam \uart_pc.data_Aux_5_LC_13_8_5 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_5_LC_13_8_5 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_Aux_5_LC_13_8_5 .LUT_INIT=16'b1111010010110000;
    LogicCell40 \uart_pc.data_Aux_5_LC_13_8_5  (
            .in0(N__28765),
            .in1(N__29088),
            .in2(N__28799),
            .in3(N__31226),
            .lcout(\uart_pc.data_AuxZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47403),
            .ce(),
            .sr(N__29109));
    defparam \uart_pc.data_Aux_6_LC_13_8_6 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_6_LC_13_8_6 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_Aux_6_LC_13_8_6 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \uart_pc.data_Aux_6_LC_13_8_6  (
            .in0(N__31992),
            .in1(N__31223),
            .in2(N__28782),
            .in3(N__28766),
            .lcout(\uart_pc.data_AuxZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47403),
            .ce(),
            .sr(N__29109));
    defparam \uart_pc.data_Aux_7_LC_13_8_7 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_7_LC_13_8_7 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_Aux_7_LC_13_8_7 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \uart_pc.data_Aux_7_LC_13_8_7  (
            .in0(N__28767),
            .in1(N__31227),
            .in2(N__29127),
            .in3(N__31772),
            .lcout(\uart_pc.data_AuxZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47403),
            .ce(),
            .sr(N__29109));
    defparam \uart_pc.data_Aux_RNO_0_3_LC_13_9_1 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_RNO_0_3_LC_13_9_1 .SEQ_MODE=4'b0000;
    defparam \uart_pc.data_Aux_RNO_0_3_LC_13_9_1 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \uart_pc.data_Aux_RNO_0_3_LC_13_9_1  (
            .in0(N__32031),
            .in1(N__32075),
            .in2(_gnd_net_),
            .in3(N__32123),
            .lcout(\uart_pc.data_Auxce_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_Aux_RNO_0_2_LC_13_9_3 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_RNO_0_2_LC_13_9_3 .SEQ_MODE=4'b0000;
    defparam \uart_pc.data_Aux_RNO_0_2_LC_13_9_3 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \uart_pc.data_Aux_RNO_0_2_LC_13_9_3  (
            .in0(N__32030),
            .in1(N__32074),
            .in2(_gnd_net_),
            .in3(N__32122),
            .lcout(\uart_pc.data_Auxce_0_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_Aux_RNO_0_5_LC_13_9_7 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_RNO_0_5_LC_13_9_7 .SEQ_MODE=4'b0000;
    defparam \uart_pc.data_Aux_RNO_0_5_LC_13_9_7 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \uart_pc.data_Aux_RNO_0_5_LC_13_9_7  (
            .in0(N__32032),
            .in1(N__32076),
            .in2(_gnd_net_),
            .in3(N__32124),
            .lcout(\uart_pc.data_Auxce_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_5_LC_13_10_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_5_LC_13_10_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_5_LC_13_10_0 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.throttle_5_LC_13_10_0  (
            .in0(N__29235),
            .in1(N__29259),
            .in2(N__37261),
            .in3(N__35218),
            .lcout(\ppm_encoder_1.throttleZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47375),
            .ce(),
            .sr(N__43823));
    defparam \scaler_2.source_data_1_4_LC_13_10_1 .C_ON=1'b0;
    defparam \scaler_2.source_data_1_4_LC_13_10_1 .SEQ_MODE=4'b1000;
    defparam \scaler_2.source_data_1_4_LC_13_10_1 .LUT_INIT=16'b0111001011011000;
    LogicCell40 \scaler_2.source_data_1_4_LC_13_10_1  (
            .in0(N__30566),
            .in1(N__29079),
            .in2(N__29180),
            .in3(N__29051),
            .lcout(scaler_2_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47375),
            .ce(),
            .sr(N__43823));
    defparam \scaler_3.source_data_1_4_LC_13_10_3 .C_ON=1'b0;
    defparam \scaler_3.source_data_1_4_LC_13_10_3 .SEQ_MODE=4'b1000;
    defparam \scaler_3.source_data_1_4_LC_13_10_3 .LUT_INIT=16'b0111001011011000;
    LogicCell40 \scaler_3.source_data_1_4_LC_13_10_3  (
            .in0(N__30567),
            .in1(N__28989),
            .in2(N__29156),
            .in3(N__28952),
            .lcout(scaler_3_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47375),
            .ce(),
            .sr(N__43823));
    defparam \scaler_2.source_data_1_esr_5_LC_13_11_0 .C_ON=1'b0;
    defparam \scaler_2.source_data_1_esr_5_LC_13_11_0 .SEQ_MODE=4'b1000;
    defparam \scaler_2.source_data_1_esr_5_LC_13_11_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \scaler_2.source_data_1_esr_5_LC_13_11_0  (
            .in0(N__32278),
            .in1(N__29080),
            .in2(_gnd_net_),
            .in3(N__29052),
            .lcout(scaler_2_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47363),
            .ce(N__32406),
            .sr(N__43829));
    defparam \scaler_3.source_data_1_esr_5_LC_13_11_1 .C_ON=1'b0;
    defparam \scaler_3.source_data_1_esr_5_LC_13_11_1 .SEQ_MODE=4'b1000;
    defparam \scaler_3.source_data_1_esr_5_LC_13_11_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \scaler_3.source_data_1_esr_5_LC_13_11_1  (
            .in0(N__29019),
            .in1(N__28988),
            .in2(_gnd_net_),
            .in3(N__28953),
            .lcout(scaler_3_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47363),
            .ce(N__32406),
            .sr(N__43829));
    defparam \scaler_4.source_data_1_esr_5_LC_13_11_2 .C_ON=1'b0;
    defparam \scaler_4.source_data_1_esr_5_LC_13_11_2 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_5_LC_13_11_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \scaler_4.source_data_1_esr_5_LC_13_11_2  (
            .in0(N__28917),
            .in1(N__29556),
            .in2(_gnd_net_),
            .in3(N__29517),
            .lcout(scaler_4_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47363),
            .ce(N__32406),
            .sr(N__43829));
    defparam \uart_pc.data_Aux_RNO_0_0_LC_13_11_3 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_RNO_0_0_LC_13_11_3 .SEQ_MODE=4'b0000;
    defparam \uart_pc.data_Aux_RNO_0_0_LC_13_11_3 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \uart_pc.data_Aux_RNO_0_0_LC_13_11_3  (
            .in0(N__32071),
            .in1(N__32119),
            .in2(_gnd_net_),
            .in3(N__32025),
            .lcout(\uart_pc.data_Auxce_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_Aux_RNO_0_1_LC_13_11_4 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_RNO_0_1_LC_13_11_4 .SEQ_MODE=4'b0000;
    defparam \uart_pc.data_Aux_RNO_0_1_LC_13_11_4 .LUT_INIT=16'b0000000000001010;
    LogicCell40 \uart_pc.data_Aux_RNO_0_1_LC_13_11_4  (
            .in0(N__32120),
            .in1(_gnd_net_),
            .in2(N__32034),
            .in3(N__32072),
            .lcout(\uart_pc.data_Auxce_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_Aux_RNO_0_4_LC_13_11_7 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_RNO_0_4_LC_13_11_7 .SEQ_MODE=4'b0000;
    defparam \uart_pc.data_Aux_RNO_0_4_LC_13_11_7 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \uart_pc.data_Aux_RNO_0_4_LC_13_11_7  (
            .in0(N__32073),
            .in1(N__32121),
            .in2(_gnd_net_),
            .in3(N__32029),
            .lcout(\uart_pc.data_Auxce_0_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_esr_4_LC_13_12_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_esr_4_LC_13_12_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.aileron_esr_4_LC_13_12_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.aileron_esr_4_LC_13_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29181),
            .lcout(\ppm_encoder_1.aileronZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47348),
            .ce(N__36267),
            .sr(N__43838));
    defparam \ppm_encoder_1.aileron_esr_5_LC_13_12_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_esr_5_LC_13_12_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.aileron_esr_5_LC_13_12_1 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \ppm_encoder_1.aileron_esr_5_LC_13_12_1  (
            .in0(_gnd_net_),
            .in1(N__29163),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\ppm_encoder_1.aileronZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47348),
            .ce(N__36267),
            .sr(N__43838));
    defparam \ppm_encoder_1.elevator_esr_4_LC_13_12_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_esr_4_LC_13_12_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.elevator_esr_4_LC_13_12_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.elevator_esr_4_LC_13_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29157),
            .lcout(\ppm_encoder_1.elevatorZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47348),
            .ce(N__36267),
            .sr(N__43838));
    defparam \ppm_encoder_1.elevator_esr_5_LC_13_12_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_esr_5_LC_13_12_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.elevator_esr_5_LC_13_12_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.elevator_esr_5_LC_13_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29139),
            .lcout(\ppm_encoder_1.elevatorZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47348),
            .ce(N__36267),
            .sr(N__43838));
    defparam \ppm_encoder_1.rudder_esr_4_LC_13_12_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_esr_4_LC_13_12_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.rudder_esr_4_LC_13_12_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.rudder_esr_4_LC_13_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29475),
            .lcout(\ppm_encoder_1.rudderZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47348),
            .ce(N__36267),
            .sr(N__43838));
    defparam \ppm_encoder_1.rudder_esr_5_LC_13_12_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_esr_5_LC_13_12_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.rudder_esr_5_LC_13_12_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.rudder_esr_5_LC_13_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29133),
            .lcout(\ppm_encoder_1.rudderZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47348),
            .ce(N__36267),
            .sr(N__43838));
    defparam \ppm_encoder_1.un1_throttle_cry_0_c_LC_13_13_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_0_c_LC_13_13_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_0_c_LC_13_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_0_c_LC_13_13_0  (
            .in0(_gnd_net_),
            .in1(N__36988),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_13_13_0_),
            .carryout(\ppm_encoder_1.un1_throttle_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_0_THRU_LUT4_0_LC_13_13_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_0_THRU_LUT4_0_LC_13_13_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_0_THRU_LUT4_0_LC_13_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_0_THRU_LUT4_0_LC_13_13_1  (
            .in0(_gnd_net_),
            .in1(N__29296),
            .in2(N__42994),
            .in3(N__29271),
            .lcout(\ppm_encoder_1.un1_throttle_cry_0_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_0 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_1_THRU_LUT4_0_LC_13_13_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_1_THRU_LUT4_0_LC_13_13_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_1_THRU_LUT4_0_LC_13_13_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_1_THRU_LUT4_0_LC_13_13_2  (
            .in0(_gnd_net_),
            .in1(N__29341),
            .in2(_gnd_net_),
            .in3(N__29268),
            .lcout(\ppm_encoder_1.un1_throttle_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_1 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_2_THRU_LUT4_0_LC_13_13_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_2_THRU_LUT4_0_LC_13_13_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_2_THRU_LUT4_0_LC_13_13_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_2_THRU_LUT4_0_LC_13_13_3  (
            .in0(_gnd_net_),
            .in1(N__35473),
            .in2(N__42995),
            .in3(N__29265),
            .lcout(\ppm_encoder_1.un1_throttle_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_2 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_3_THRU_LUT4_0_LC_13_13_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_3_THRU_LUT4_0_LC_13_13_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_3_THRU_LUT4_0_LC_13_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_3_THRU_LUT4_0_LC_13_13_4  (
            .in0(_gnd_net_),
            .in1(N__29392),
            .in2(_gnd_net_),
            .in3(N__29262),
            .lcout(\ppm_encoder_1.un1_throttle_cry_3_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_3 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_4_THRU_LUT4_0_LC_13_13_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_4_THRU_LUT4_0_LC_13_13_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_4_THRU_LUT4_0_LC_13_13_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_4_THRU_LUT4_0_LC_13_13_5  (
            .in0(_gnd_net_),
            .in1(N__29258),
            .in2(_gnd_net_),
            .in3(N__29226),
            .lcout(\ppm_encoder_1.un1_throttle_cry_4_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_4 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_5_THRU_LUT4_0_LC_13_13_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_5_THRU_LUT4_0_LC_13_13_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_5_THRU_LUT4_0_LC_13_13_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_5_THRU_LUT4_0_LC_13_13_6  (
            .in0(_gnd_net_),
            .in1(N__42923),
            .in2(N__34307),
            .in3(N__29223),
            .lcout(\ppm_encoder_1.un1_throttle_cry_5_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_5 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_6_THRU_LUT4_0_LC_13_13_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_6_THRU_LUT4_0_LC_13_13_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_6_THRU_LUT4_0_LC_13_13_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_6_THRU_LUT4_0_LC_13_13_7  (
            .in0(_gnd_net_),
            .in1(N__31892),
            .in2(_gnd_net_),
            .in3(N__29220),
            .lcout(\ppm_encoder_1.un1_throttle_cry_6_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_6 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_7_THRU_LUT4_0_LC_13_14_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_7_THRU_LUT4_0_LC_13_14_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_7_THRU_LUT4_0_LC_13_14_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_7_THRU_LUT4_0_LC_13_14_0  (
            .in0(_gnd_net_),
            .in1(N__34223),
            .in2(_gnd_net_),
            .in3(N__29217),
            .lcout(\ppm_encoder_1.un1_throttle_cry_7_THRU_CO ),
            .ltout(),
            .carryin(bfn_13_14_0_),
            .carryout(\ppm_encoder_1.un1_throttle_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_8_THRU_LUT4_0_LC_13_14_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_8_THRU_LUT4_0_LC_13_14_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_8_THRU_LUT4_0_LC_13_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_8_THRU_LUT4_0_LC_13_14_1  (
            .in0(_gnd_net_),
            .in1(N__32588),
            .in2(_gnd_net_),
            .in3(N__29367),
            .lcout(\ppm_encoder_1.un1_throttle_cry_8_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_8 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_9_THRU_LUT4_0_LC_13_14_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_9_THRU_LUT4_0_LC_13_14_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_9_THRU_LUT4_0_LC_13_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_9_THRU_LUT4_0_LC_13_14_2  (
            .in0(_gnd_net_),
            .in1(N__29435),
            .in2(_gnd_net_),
            .in3(N__29364),
            .lcout(\ppm_encoder_1.un1_throttle_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_9 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_10_THRU_LUT4_0_LC_13_14_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_10_THRU_LUT4_0_LC_13_14_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_10_THRU_LUT4_0_LC_13_14_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_10_THRU_LUT4_0_LC_13_14_3  (
            .in0(_gnd_net_),
            .in1(N__32723),
            .in2(_gnd_net_),
            .in3(N__29361),
            .lcout(\ppm_encoder_1.un1_throttle_cry_10_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_10 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_11_THRU_LUT4_0_LC_13_14_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_11_THRU_LUT4_0_LC_13_14_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_11_THRU_LUT4_0_LC_13_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_11_THRU_LUT4_0_LC_13_14_4  (
            .in0(_gnd_net_),
            .in1(N__32492),
            .in2(_gnd_net_),
            .in3(N__29358),
            .lcout(\ppm_encoder_1.un1_throttle_cry_11_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_11 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_12_THRU_LUT4_0_LC_13_14_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_12_THRU_LUT4_0_LC_13_14_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_12_THRU_LUT4_0_LC_13_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_12_THRU_LUT4_0_LC_13_14_5  (
            .in0(_gnd_net_),
            .in1(N__34460),
            .in2(N__43081),
            .in3(N__29355),
            .lcout(\ppm_encoder_1.un1_throttle_cry_12_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_12 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_esr_14_LC_13_14_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_esr_14_LC_13_14_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_esr_14_LC_13_14_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.throttle_esr_14_LC_13_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29352),
            .lcout(\ppm_encoder_1.throttleZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47318),
            .ce(N__36262),
            .sr(N__43853));
    defparam \ppm_encoder_1.throttle_2_LC_13_15_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_2_LC_13_15_0 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.throttle_2_LC_13_15_0 .LUT_INIT=16'b0111001011011000;
    LogicCell40 \ppm_encoder_1.throttle_2_LC_13_15_0  (
            .in0(N__37091),
            .in1(N__29349),
            .in2(N__37631),
            .in3(N__29319),
            .lcout(\ppm_encoder_1.throttleZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47308),
            .ce(),
            .sr(N__43859));
    defparam \ppm_encoder_1.pulses2count_16_LC_13_15_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_16_LC_13_15_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_16_LC_13_15_1 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \ppm_encoder_1.pulses2count_16_LC_13_15_1  (
            .in0(N__40809),
            .in1(N__39773),
            .in2(N__39738),
            .in3(N__41892),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47308),
            .ce(),
            .sr(N__43859));
    defparam \ppm_encoder_1.throttle_1_LC_13_15_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_1_LC_13_15_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_1_LC_13_15_2 .LUT_INIT=16'b1001111110010000;
    LogicCell40 \ppm_encoder_1.throttle_1_LC_13_15_2  (
            .in0(N__29310),
            .in1(N__29301),
            .in2(N__37148),
            .in3(N__34570),
            .lcout(\ppm_encoder_1.throttleZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47308),
            .ce(),
            .sr(N__43859));
    defparam \ppm_encoder_1.rudder_6_LC_13_15_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_6_LC_13_15_3 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.rudder_6_LC_13_15_3 .LUT_INIT=16'b0111011101000100;
    LogicCell40 \ppm_encoder_1.rudder_6_LC_13_15_3  (
            .in0(N__29790),
            .in1(N__37092),
            .in2(_gnd_net_),
            .in3(N__36205),
            .lcout(\ppm_encoder_1.rudderZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47308),
            .ce(),
            .sr(N__43859));
    defparam \dron_frame_decoder_1.source_data_valid_LC_13_15_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_data_valid_LC_13_15_4 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_data_valid_LC_13_15_4 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \dron_frame_decoder_1.source_data_valid_LC_13_15_4  (
            .in0(N__29721),
            .in1(N__29676),
            .in2(_gnd_net_),
            .in3(N__29577),
            .lcout(debug_CH1_0A_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47308),
            .ce(),
            .sr(N__43859));
    defparam \scaler_4.source_data_1_4_LC_13_15_7 .C_ON=1'b0;
    defparam \scaler_4.source_data_1_4_LC_13_15_7 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_4_LC_13_15_7 .LUT_INIT=16'b0111001011011000;
    LogicCell40 \scaler_4.source_data_1_4_LC_13_15_7  (
            .in0(N__30577),
            .in1(N__29552),
            .in2(N__29474),
            .in3(N__29513),
            .lcout(scaler_4_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47308),
            .ce(),
            .sr(N__43859));
    defparam \ppm_encoder_1.ppm_output_reg_LC_13_16_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.ppm_output_reg_LC_13_16_0 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.ppm_output_reg_LC_13_16_0 .LUT_INIT=16'b1111001111010000;
    LogicCell40 \ppm_encoder_1.ppm_output_reg_LC_13_16_0  (
            .in0(N__34680),
            .in1(N__32868),
            .in2(N__29453),
            .in3(N__39042),
            .lcout(ppm_output_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47298),
            .ce(),
            .sr(N__43868));
    defparam \ppm_encoder_1.rudder_7_LC_13_16_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_7_LC_13_16_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.rudder_7_LC_13_16_2 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \ppm_encoder_1.rudder_7_LC_13_16_2  (
            .in0(N__29766),
            .in1(N__29778),
            .in2(N__40690),
            .in3(N__37102),
            .lcout(\ppm_encoder_1.rudderZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47298),
            .ce(),
            .sr(N__43868));
    defparam \ppm_encoder_1.rudder_9_LC_13_16_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_9_LC_13_16_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.rudder_9_LC_13_16_3 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.rudder_9_LC_13_16_3  (
            .in0(N__29742),
            .in1(N__29754),
            .in2(N__37150),
            .in3(N__40535),
            .lcout(\ppm_encoder_1.rudderZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47298),
            .ce(),
            .sr(N__43868));
    defparam \ppm_encoder_1.throttle_10_LC_13_16_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_10_LC_13_16_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_10_LC_13_16_4 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \ppm_encoder_1.throttle_10_LC_13_16_4  (
            .in0(N__29436),
            .in1(N__29418),
            .in2(N__32618),
            .in3(N__37103),
            .lcout(\ppm_encoder_1.throttleZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47298),
            .ce(),
            .sr(N__43868));
    defparam \ppm_encoder_1.elevator_8_LC_13_16_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_8_LC_13_16_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.elevator_8_LC_13_16_5 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.elevator_8_LC_13_16_5  (
            .in0(N__29817),
            .in1(N__29834),
            .in2(N__37149),
            .in3(N__34241),
            .lcout(\ppm_encoder_1.elevatorZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47298),
            .ce(),
            .sr(N__43868));
    defparam \ppm_encoder_1.throttle_4_LC_13_16_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_4_LC_13_16_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_4_LC_13_16_6 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \ppm_encoder_1.throttle_4_LC_13_16_6  (
            .in0(N__29409),
            .in1(N__29400),
            .in2(N__35374),
            .in3(N__37104),
            .lcout(\ppm_encoder_1.throttleZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47298),
            .ce(),
            .sr(N__43868));
    defparam \ppm_encoder_1.un1_rudder_cry_6_c_LC_13_17_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_rudder_cry_6_c_LC_13_17_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_rudder_cry_6_c_LC_13_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.un1_rudder_cry_6_c_LC_13_17_0  (
            .in0(_gnd_net_),
            .in1(N__29789),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_13_17_0_),
            .carryout(\ppm_encoder_1.un1_rudder_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_rudder_cry_6_THRU_LUT4_0_LC_13_17_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_rudder_cry_6_THRU_LUT4_0_LC_13_17_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_rudder_cry_6_THRU_LUT4_0_LC_13_17_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_rudder_cry_6_THRU_LUT4_0_LC_13_17_1  (
            .in0(_gnd_net_),
            .in1(N__29777),
            .in2(_gnd_net_),
            .in3(N__29760),
            .lcout(\ppm_encoder_1.un1_rudder_cry_6_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_rudder_cry_6 ),
            .carryout(\ppm_encoder_1.un1_rudder_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_rudder_cry_7_THRU_LUT4_0_LC_13_17_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_rudder_cry_7_THRU_LUT4_0_LC_13_17_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_rudder_cry_7_THRU_LUT4_0_LC_13_17_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_rudder_cry_7_THRU_LUT4_0_LC_13_17_2  (
            .in0(_gnd_net_),
            .in1(N__34520),
            .in2(_gnd_net_),
            .in3(N__29757),
            .lcout(\ppm_encoder_1.un1_rudder_cry_7_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_rudder_cry_7 ),
            .carryout(\ppm_encoder_1.un1_rudder_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_rudder_cry_8_THRU_LUT4_0_LC_13_17_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_rudder_cry_8_THRU_LUT4_0_LC_13_17_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_rudder_cry_8_THRU_LUT4_0_LC_13_17_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_rudder_cry_8_THRU_LUT4_0_LC_13_17_3  (
            .in0(_gnd_net_),
            .in1(N__29753),
            .in2(_gnd_net_),
            .in3(N__29736),
            .lcout(\ppm_encoder_1.un1_rudder_cry_8_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_rudder_cry_8 ),
            .carryout(\ppm_encoder_1.un1_rudder_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_rudder_cry_9_THRU_LUT4_0_LC_13_17_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_rudder_cry_9_THRU_LUT4_0_LC_13_17_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_rudder_cry_9_THRU_LUT4_0_LC_13_17_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_rudder_cry_9_THRU_LUT4_0_LC_13_17_4  (
            .in0(_gnd_net_),
            .in1(N__32960),
            .in2(_gnd_net_),
            .in3(N__29733),
            .lcout(\ppm_encoder_1.un1_rudder_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_rudder_cry_9 ),
            .carryout(\ppm_encoder_1.un1_rudder_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_rudder_cry_10_THRU_LUT4_0_LC_13_17_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_rudder_cry_10_THRU_LUT4_0_LC_13_17_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_rudder_cry_10_THRU_LUT4_0_LC_13_17_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_rudder_cry_10_THRU_LUT4_0_LC_13_17_5  (
            .in0(_gnd_net_),
            .in1(N__32741),
            .in2(_gnd_net_),
            .in3(N__29730),
            .lcout(\ppm_encoder_1.un1_rudder_cry_10_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_rudder_cry_10 ),
            .carryout(\ppm_encoder_1.un1_rudder_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_rudder_cry_11_THRU_LUT4_0_LC_13_17_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_rudder_cry_11_THRU_LUT4_0_LC_13_17_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_rudder_cry_11_THRU_LUT4_0_LC_13_17_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_rudder_cry_11_THRU_LUT4_0_LC_13_17_6  (
            .in0(_gnd_net_),
            .in1(N__32654),
            .in2(_gnd_net_),
            .in3(N__29727),
            .lcout(\ppm_encoder_1.un1_rudder_cry_11_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_rudder_cry_11 ),
            .carryout(\ppm_encoder_1.un1_rudder_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_rudder_cry_12_THRU_LUT4_0_LC_13_17_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_rudder_cry_12_THRU_LUT4_0_LC_13_17_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_rudder_cry_12_THRU_LUT4_0_LC_13_17_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_rudder_cry_12_THRU_LUT4_0_LC_13_17_7  (
            .in0(_gnd_net_),
            .in1(N__36290),
            .in2(N__42885),
            .in3(N__29724),
            .lcout(\ppm_encoder_1.un1_rudder_cry_12_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_rudder_cry_12 ),
            .carryout(\ppm_encoder_1.un1_rudder_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.rudder_esr_14_LC_13_18_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_esr_14_LC_13_18_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.rudder_esr_14_LC_13_18_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ppm_encoder_1.rudder_esr_14_LC_13_18_0  (
            .in0(_gnd_net_),
            .in1(N__29847),
            .in2(_gnd_net_),
            .in3(N__29841),
            .lcout(\ppm_encoder_1.rudderZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47284),
            .ce(N__36244),
            .sr(N__43882));
    defparam \ppm_encoder_1.un1_elevator_cry_6_c_LC_13_19_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_6_c_LC_13_19_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_6_c_LC_13_19_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_6_c_LC_13_19_0  (
            .in0(_gnd_net_),
            .in1(N__34356),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_13_19_0_),
            .carryout(\ppm_encoder_1.un1_elevator_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_6_THRU_LUT4_0_LC_13_19_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_6_THRU_LUT4_0_LC_13_19_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_6_THRU_LUT4_0_LC_13_19_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_6_THRU_LUT4_0_LC_13_19_1  (
            .in0(_gnd_net_),
            .in1(N__31943),
            .in2(_gnd_net_),
            .in3(N__29838),
            .lcout(\ppm_encoder_1.un1_elevator_cry_6_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_6 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_7_THRU_LUT4_0_LC_13_19_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_7_THRU_LUT4_0_LC_13_19_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_7_THRU_LUT4_0_LC_13_19_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_7_THRU_LUT4_0_LC_13_19_2  (
            .in0(_gnd_net_),
            .in1(N__29835),
            .in2(_gnd_net_),
            .in3(N__29808),
            .lcout(\ppm_encoder_1.un1_elevator_cry_7_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_7 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_8_THRU_LUT4_0_LC_13_19_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_8_THRU_LUT4_0_LC_13_19_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_8_THRU_LUT4_0_LC_13_19_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_8_THRU_LUT4_0_LC_13_19_3  (
            .in0(_gnd_net_),
            .in1(N__32351),
            .in2(_gnd_net_),
            .in3(N__29805),
            .lcout(\ppm_encoder_1.un1_elevator_cry_8_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_8 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_9_THRU_LUT4_0_LC_13_19_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_9_THRU_LUT4_0_LC_13_19_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_9_THRU_LUT4_0_LC_13_19_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_9_THRU_LUT4_0_LC_13_19_4  (
            .in0(_gnd_net_),
            .in1(N__33011),
            .in2(_gnd_net_),
            .in3(N__29802),
            .lcout(\ppm_encoder_1.un1_elevator_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_9 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_10_THRU_LUT4_0_LC_13_19_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_10_THRU_LUT4_0_LC_13_19_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_10_THRU_LUT4_0_LC_13_19_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_10_THRU_LUT4_0_LC_13_19_5  (
            .in0(_gnd_net_),
            .in1(N__32696),
            .in2(_gnd_net_),
            .in3(N__29799),
            .lcout(\ppm_encoder_1.un1_elevator_cry_10_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_10 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_11_THRU_LUT4_0_LC_13_19_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_11_THRU_LUT4_0_LC_13_19_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_11_THRU_LUT4_0_LC_13_19_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_11_THRU_LUT4_0_LC_13_19_6  (
            .in0(_gnd_net_),
            .in1(N__32528),
            .in2(_gnd_net_),
            .in3(N__29796),
            .lcout(\ppm_encoder_1.un1_elevator_cry_11_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_11 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_12_THRU_LUT4_0_LC_13_19_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_12_THRU_LUT4_0_LC_13_19_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_12_THRU_LUT4_0_LC_13_19_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_12_THRU_LUT4_0_LC_13_19_7  (
            .in0(_gnd_net_),
            .in1(N__34499),
            .in2(N__43020),
            .in3(N__29793),
            .lcout(\ppm_encoder_1.un1_elevator_cry_12_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_12 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_esr_14_LC_13_20_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_esr_14_LC_13_20_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.elevator_esr_14_LC_13_20_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ppm_encoder_1.elevator_esr_14_LC_13_20_0  (
            .in0(_gnd_net_),
            .in1(N__30153),
            .in2(_gnd_net_),
            .in3(N__30141),
            .lcout(\ppm_encoder_1.elevatorZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47272),
            .ce(N__36266),
            .sr(N__43890));
    defparam \pid_alt.error_i_acumm_esr_RNIB9IP_0_LC_13_21_0 .C_ON=1'b1;
    defparam \pid_alt.error_i_acumm_esr_RNIB9IP_0_LC_13_21_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_esr_RNIB9IP_0_LC_13_21_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \pid_alt.error_i_acumm_esr_RNIB9IP_0_LC_13_21_0  (
            .in0(_gnd_net_),
            .in1(N__33665),
            .in2(N__39585),
            .in3(_gnd_net_),
            .lcout(\pid_alt.un1_pid_prereg_0 ),
            .ltout(),
            .carryin(bfn_13_21_0_),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_esr_RNIQMD91_1_LC_13_21_1 .C_ON=1'b1;
    defparam \pid_alt.error_i_acumm_esr_RNIQMD91_1_LC_13_21_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_esr_RNIQMD91_1_LC_13_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_i_acumm_esr_RNIQMD91_1_LC_13_21_1  (
            .in0(_gnd_net_),
            .in1(N__30108),
            .in2(N__34866),
            .in3(N__30048),
            .lcout(\pid_alt.error_i_acumm_esr_RNIQMD91Z0Z_1 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_0 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_esr_RNITQE91_2_LC_13_21_2 .C_ON=1'b1;
    defparam \pid_alt.error_i_acumm_esr_RNITQE91_2_LC_13_21_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_esr_RNITQE91_2_LC_13_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_i_acumm_esr_RNITQE91_2_LC_13_21_2  (
            .in0(_gnd_net_),
            .in1(N__30045),
            .in2(N__36729),
            .in3(N__30006),
            .lcout(\pid_alt.error_i_acumm_esr_RNITQE91Z0Z_2 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_1 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_esr_RNI0VF91_3_LC_13_21_3 .C_ON=1'b1;
    defparam \pid_alt.error_i_acumm_esr_RNI0VF91_3_LC_13_21_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_esr_RNI0VF91_3_LC_13_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_i_acumm_esr_RNI0VF91_3_LC_13_21_3  (
            .in0(_gnd_net_),
            .in1(N__30003),
            .in2(N__39552),
            .in3(N__29958),
            .lcout(\pid_alt.error_i_acumm_esr_RNI0VF91Z0Z_3 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_2 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_esr_RNI33H91_4_LC_13_21_4 .C_ON=1'b1;
    defparam \pid_alt.error_i_acumm_esr_RNI33H91_4_LC_13_21_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_esr_RNI33H91_4_LC_13_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_i_acumm_esr_RNI33H91_4_LC_13_21_4  (
            .in0(_gnd_net_),
            .in1(N__29955),
            .in2(N__43206),
            .in3(N__29928),
            .lcout(\pid_alt.error_i_acumm_esr_RNI33H91Z0Z_4 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_3 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_reg_esr_RNIT8KA1_5_LC_13_21_5 .C_ON=1'b1;
    defparam \pid_alt.error_i_reg_esr_RNIT8KA1_5_LC_13_21_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_reg_esr_RNIT8KA1_5_LC_13_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_i_reg_esr_RNIT8KA1_5_LC_13_21_5  (
            .in0(_gnd_net_),
            .in1(N__45408),
            .in2(N__29925),
            .in3(N__29883),
            .lcout(\pid_alt.error_i_reg_esr_RNIT8KA1Z0Z_5 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_4 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_5_c_RNI0DLQ_LC_13_21_6 .C_ON=1'b1;
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_5_c_RNI0DLQ_LC_13_21_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_5_c_RNI0DLQ_LC_13_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_5_c_RNI0DLQ_LC_13_21_6  (
            .in0(_gnd_net_),
            .in1(N__46215),
            .in2(N__33261),
            .in3(N__29850),
            .lcout(\pid_alt.un1_error_i_acumm_prereg_cry_5_c_RNI0DLQ ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_5 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_6_c_RNI3HMQ_LC_13_21_7 .C_ON=1'b1;
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_6_c_RNI3HMQ_LC_13_21_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_6_c_RNI3HMQ_LC_13_21_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_6_c_RNI3HMQ_LC_13_21_7  (
            .in0(_gnd_net_),
            .in1(N__30498),
            .in2(N__46239),
            .in3(N__30447),
            .lcout(\pid_alt.un1_error_i_acumm_prereg_cry_6_c_RNI3HMQ ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_6 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_7_c_RNI6LNQ_LC_13_22_0 .C_ON=1'b1;
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_7_c_RNI6LNQ_LC_13_22_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_7_c_RNI6LNQ_LC_13_22_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_7_c_RNI6LNQ_LC_13_22_0  (
            .in0(_gnd_net_),
            .in1(N__30443),
            .in2(N__45384),
            .in3(N__30402),
            .lcout(\pid_alt.un1_error_i_acumm_prereg_cry_7_c_RNI6LNQ ),
            .ltout(),
            .carryin(bfn_13_22_0_),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_8_c_RNI9POQ_LC_13_22_1 .C_ON=1'b1;
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_8_c_RNI9POQ_LC_13_22_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_8_c_RNI9POQ_LC_13_22_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_8_c_RNI9POQ_LC_13_22_1  (
            .in0(_gnd_net_),
            .in1(N__47616),
            .in2(N__30395),
            .in3(N__30357),
            .lcout(\pid_alt.un1_error_i_acumm_prereg_cry_8_c_RNI9POQ ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_8 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_9_c_RNIQN3F_LC_13_22_2 .C_ON=1'b1;
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_9_c_RNIQN3F_LC_13_22_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_9_c_RNIQN3F_LC_13_22_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_9_c_RNIQN3F_LC_13_22_2  (
            .in0(_gnd_net_),
            .in1(N__30350),
            .in2(N__44760),
            .in3(N__30303),
            .lcout(\pid_alt.un1_error_i_acumm_prereg_cry_9_c_RNIQN3F ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_9 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_reg_esr_RNI4NMP_11_LC_13_22_3 .C_ON=1'b1;
    defparam \pid_alt.error_i_reg_esr_RNI4NMP_11_LC_13_22_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_reg_esr_RNI4NMP_11_LC_13_22_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_i_reg_esr_RNI4NMP_11_LC_13_22_3  (
            .in0(_gnd_net_),
            .in1(N__33026),
            .in2(N__44727),
            .in3(N__30270),
            .lcout(\pid_alt.error_i_reg_esr_RNI4NMPZ0Z_11 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_10 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_reg_esr_RNI7RNP_12_LC_13_22_4 .C_ON=1'b1;
    defparam \pid_alt.error_i_reg_esr_RNI7RNP_12_LC_13_22_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_reg_esr_RNI7RNP_12_LC_13_22_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_i_reg_esr_RNI7RNP_12_LC_13_22_4  (
            .in0(_gnd_net_),
            .in1(N__30266),
            .in2(N__44694),
            .in3(N__30222),
            .lcout(\pid_alt.error_i_reg_esr_RNI7RNPZ0Z_12 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_11 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_esr_RNIJ6LM_13_LC_13_22_5 .C_ON=1'b1;
    defparam \pid_alt.error_i_acumm_esr_RNIJ6LM_13_LC_13_22_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_esr_RNIJ6LM_13_LC_13_22_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_i_acumm_esr_RNIJ6LM_13_LC_13_22_5  (
            .in0(_gnd_net_),
            .in1(N__32784),
            .in2(N__45819),
            .in3(N__30189),
            .lcout(\pid_alt.error_i_acumm_esr_RNIJ6LMZ0Z_13 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_12 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_reg_esr_RNI15KJ_14_LC_13_22_6 .C_ON=1'b1;
    defparam \pid_alt.error_i_reg_esr_RNI15KJ_14_LC_13_22_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_reg_esr_RNI15KJ_14_LC_13_22_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_i_reg_esr_RNI15KJ_14_LC_13_22_6  (
            .in0(_gnd_net_),
            .in1(N__47595),
            .in2(_gnd_net_),
            .in3(N__30156),
            .lcout(\pid_alt.error_i_reg_esr_RNI15KJZ0Z_14 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_13 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_reg_esr_RNI38LJ_15_LC_13_22_7 .C_ON=1'b1;
    defparam \pid_alt.error_i_reg_esr_RNI38LJ_15_LC_13_22_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_reg_esr_RNI38LJ_15_LC_13_22_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_i_reg_esr_RNI38LJ_15_LC_13_22_7  (
            .in0(_gnd_net_),
            .in1(N__46194),
            .in2(_gnd_net_),
            .in3(N__30918),
            .lcout(\pid_alt.error_i_reg_esr_RNI38LJZ0Z_15 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_14 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_reg_esr_RNI5BMJ_16_LC_13_23_0 .C_ON=1'b1;
    defparam \pid_alt.error_i_reg_esr_RNI5BMJ_16_LC_13_23_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_reg_esr_RNI5BMJ_16_LC_13_23_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_i_reg_esr_RNI5BMJ_16_LC_13_23_0  (
            .in0(_gnd_net_),
            .in1(N__47511),
            .in2(_gnd_net_),
            .in3(N__30885),
            .lcout(\pid_alt.error_i_reg_esr_RNI5BMJZ0Z_16 ),
            .ltout(),
            .carryin(bfn_13_23_0_),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_reg_esr_RNI7ENJ_17_LC_13_23_1 .C_ON=1'b1;
    defparam \pid_alt.error_i_reg_esr_RNI7ENJ_17_LC_13_23_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_reg_esr_RNI7ENJ_17_LC_13_23_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_i_reg_esr_RNI7ENJ_17_LC_13_23_1  (
            .in0(_gnd_net_),
            .in1(N__47553),
            .in2(_gnd_net_),
            .in3(N__30849),
            .lcout(\pid_alt.error_i_reg_esr_RNI7ENJZ0Z_17 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_16 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_reg_esr_RNI9HOJ_18_LC_13_23_2 .C_ON=1'b1;
    defparam \pid_alt.error_i_reg_esr_RNI9HOJ_18_LC_13_23_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_reg_esr_RNI9HOJ_18_LC_13_23_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_i_reg_esr_RNI9HOJ_18_LC_13_23_2  (
            .in0(_gnd_net_),
            .in1(N__47532),
            .in2(_gnd_net_),
            .in3(N__30813),
            .lcout(\pid_alt.error_i_reg_esr_RNI9HOJZ0Z_18 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_17 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_reg_esr_RNIBKPJ_19_LC_13_23_3 .C_ON=1'b1;
    defparam \pid_alt.error_i_reg_esr_RNIBKPJ_19_LC_13_23_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_reg_esr_RNIBKPJ_19_LC_13_23_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_i_reg_esr_RNIBKPJ_19_LC_13_23_3  (
            .in0(_gnd_net_),
            .in1(N__47496),
            .in2(_gnd_net_),
            .in3(N__30774),
            .lcout(\pid_alt.error_i_reg_esr_RNIBKPJZ0Z_19 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_18 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_19_c_RNI4FRJ_LC_13_23_4 .C_ON=1'b1;
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_19_c_RNI4FRJ_LC_13_23_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_19_c_RNI4FRJ_LC_13_23_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_19_c_RNI4FRJ_LC_13_23_4  (
            .in0(_gnd_net_),
            .in1(N__47576),
            .in2(_gnd_net_),
            .in3(N__30726),
            .lcout(\pid_alt.un1_error_i_acumm_prereg_cry_19_c_RNI4FRJ ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_19 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_20_c_RNISVKK_LC_13_23_5 .C_ON=1'b0;
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_20_c_RNISVKK_LC_13_23_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_20_c_RNISVKK_LC_13_23_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_20_c_RNISVKK_LC_13_23_5  (
            .in0(N__47577),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30723),
            .lcout(\pid_alt.un1_error_i_acumm_prereg_cry_20_c_RNISVKK ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_2.source_data_1_esr_ctle_14_LC_13_29_7 .C_ON=1'b0;
    defparam \scaler_2.source_data_1_esr_ctle_14_LC_13_29_7 .SEQ_MODE=4'b0000;
    defparam \scaler_2.source_data_1_esr_ctle_14_LC_13_29_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \scaler_2.source_data_1_esr_ctle_14_LC_13_29_7  (
            .in0(_gnd_net_),
            .in1(N__30579),
            .in2(_gnd_net_),
            .in3(N__44071),
            .lcout(debug_CH3_20A_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_RNO_0_0_LC_14_4_6 .C_ON=1'b0;
    defparam \uart_pc.state_RNO_0_0_LC_14_4_6 .SEQ_MODE=4'b0000;
    defparam \uart_pc.state_RNO_0_0_LC_14_4_6 .LUT_INIT=16'b0000000011011101;
    LogicCell40 \uart_pc.state_RNO_0_0_LC_14_4_6  (
            .in0(N__31244),
            .in1(N__31216),
            .in2(_gnd_net_),
            .in3(N__44101),
            .lcout(),
            .ltout(\uart_pc.state_srsts_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_0_LC_14_4_7 .C_ON=1'b0;
    defparam \uart_pc.state_0_LC_14_4_7 .SEQ_MODE=4'b1000;
    defparam \uart_pc.state_0_LC_14_4_7 .LUT_INIT=16'b1110111100001111;
    LogicCell40 \uart_pc.state_0_LC_14_4_7  (
            .in0(N__31520),
            .in1(N__31278),
            .in2(N__31260),
            .in3(N__31563),
            .lcout(\uart_pc.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47451),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_2_LC_14_6_1 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_2_LC_14_6_1 .SEQ_MODE=4'b1000;
    defparam \uart_drone.timer_Count_2_LC_14_6_1 .LUT_INIT=16'b0000000010101000;
    LogicCell40 \uart_drone.timer_Count_2_LC_14_6_1  (
            .in0(N__33489),
            .in1(N__33916),
            .in2(N__33885),
            .in3(N__44126),
            .lcout(\uart_drone.timer_CountZ1Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47435),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_0_LC_14_6_4 .C_ON=1'b0;
    defparam \uart_drone.state_0_LC_14_6_4 .SEQ_MODE=4'b1000;
    defparam \uart_drone.state_0_LC_14_6_4 .LUT_INIT=16'b1111110101010101;
    LogicCell40 \uart_drone.state_0_LC_14_6_4  (
            .in0(N__31257),
            .in1(N__36616),
            .in2(N__31452),
            .in3(N__36488),
            .lcout(\uart_drone.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47435),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_1_LC_14_6_5 .C_ON=1'b0;
    defparam \uart_pc.state_1_LC_14_6_5 .SEQ_MODE=4'b1000;
    defparam \uart_pc.state_1_LC_14_6_5 .LUT_INIT=16'b0000000011001000;
    LogicCell40 \uart_pc.state_1_LC_14_6_5  (
            .in0(N__31130),
            .in1(N__31230),
            .in2(N__31251),
            .in3(N__44127),
            .lcout(\uart_pc.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47435),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_RNI9E9J_2_LC_14_7_0 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_RNI9E9J_2_LC_14_7_0 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNI9E9J_2_LC_14_7_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uart_drone.timer_Count_RNI9E9J_2_LC_14_7_0  (
            .in0(_gnd_net_),
            .in1(N__33508),
            .in2(_gnd_net_),
            .in3(N__36531),
            .lcout(\uart_drone.N_126_li ),
            .ltout(\uart_drone.N_126_li_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_RNIAT1D1_4_LC_14_7_1 .C_ON=1'b0;
    defparam \uart_drone.state_RNIAT1D1_4_LC_14_7_1 .SEQ_MODE=4'b0000;
    defparam \uart_drone.state_RNIAT1D1_4_LC_14_7_1 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \uart_drone.state_RNIAT1D1_4_LC_14_7_1  (
            .in0(N__36605),
            .in1(N__36483),
            .in2(N__31233),
            .in3(N__44096),
            .lcout(\uart_drone.N_143 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_RNO_0_2_LC_14_7_2 .C_ON=1'b0;
    defparam \uart_pc.state_RNO_0_2_LC_14_7_2 .SEQ_MODE=4'b0000;
    defparam \uart_pc.state_RNO_0_2_LC_14_7_2 .LUT_INIT=16'b0000010001010100;
    LogicCell40 \uart_pc.state_RNO_0_2_LC_14_7_2  (
            .in0(N__44097),
            .in1(N__31101),
            .in2(N__31131),
            .in3(N__31212),
            .lcout(),
            .ltout(\uart_pc.state_srsts_i_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_2_LC_14_7_3 .C_ON=1'b0;
    defparam \uart_pc.state_2_LC_14_7_3 .SEQ_MODE=4'b1000;
    defparam \uart_pc.state_2_LC_14_7_3 .LUT_INIT=16'b1111000001110000;
    LogicCell40 \uart_pc.state_2_LC_14_7_3  (
            .in0(N__31620),
            .in1(N__31519),
            .in2(N__31134),
            .in3(N__31129),
            .lcout(\uart_pc.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47425),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_3_LC_14_7_4 .C_ON=1'b0;
    defparam \uart_pc.data_3_LC_14_7_4 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_3_LC_14_7_4 .LUT_INIT=16'b0011000010101010;
    LogicCell40 \uart_pc.data_3_LC_14_7_4  (
            .in0(N__43266),
            .in1(N__31073),
            .in2(N__31020),
            .in3(N__31002),
            .lcout(uart_pc_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47425),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNIR9N6_1_LC_14_7_5 .C_ON=1'b0;
    defparam \reset_module_System.count_RNIR9N6_1_LC_14_7_5 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNIR9N6_1_LC_14_7_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \reset_module_System.count_RNIR9N6_1_LC_14_7_5  (
            .in0(_gnd_net_),
            .in1(N__34755),
            .in2(_gnd_net_),
            .in3(N__34849),
            .lcout(\reset_module_System.reset6_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_1_LC_14_7_6 .C_ON=1'b0;
    defparam \uart_drone.state_1_LC_14_7_6 .SEQ_MODE=4'b1000;
    defparam \uart_drone.state_1_LC_14_7_6 .LUT_INIT=16'b0101010000000000;
    LogicCell40 \uart_drone.state_1_LC_14_7_6  (
            .in0(N__44098),
            .in1(N__31659),
            .in2(N__31301),
            .in3(N__31393),
            .lcout(\uart_drone.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47425),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_3_LC_14_8_3 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_3_LC_14_8_3 .SEQ_MODE=4'b1000;
    defparam \uart_drone.timer_Count_3_LC_14_8_3 .LUT_INIT=16'b0000101000001000;
    LogicCell40 \uart_drone.timer_Count_3_LC_14_8_3  (
            .in0(N__33480),
            .in1(N__33917),
            .in2(N__44138),
            .in3(N__33870),
            .lcout(\uart_drone.timer_CountZ1Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47415),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_RNIDGR31_2_LC_14_8_4 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_RNIDGR31_2_LC_14_8_4 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNIDGR31_2_LC_14_8_4 .LUT_INIT=16'b1111100000000000;
    LogicCell40 \uart_drone.timer_Count_RNIDGR31_2_LC_14_8_4  (
            .in0(N__36525),
            .in1(N__33510),
            .in2(N__36608),
            .in3(N__36475),
            .lcout(\uart_drone.data_rdyc_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_4_LC_14_8_5 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_4_LC_14_8_5 .SEQ_MODE=4'b1000;
    defparam \uart_drone.timer_Count_4_LC_14_8_5 .LUT_INIT=16'b0000101000001000;
    LogicCell40 \uart_drone.timer_Count_4_LC_14_8_5  (
            .in0(N__33462),
            .in1(N__33918),
            .in2(N__44139),
            .in3(N__33871),
            .lcout(\uart_drone.timer_CountZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47415),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_RNIITIF1_4_LC_14_8_6 .C_ON=1'b0;
    defparam \uart_pc.state_RNIITIF1_4_LC_14_8_6 .SEQ_MODE=4'b0000;
    defparam \uart_pc.state_RNIITIF1_4_LC_14_8_6 .LUT_INIT=16'b0010000000110011;
    LogicCell40 \uart_pc.state_RNIITIF1_4_LC_14_8_6  (
            .in0(N__31619),
            .in1(N__31562),
            .in2(N__31521),
            .in3(N__31723),
            .lcout(\uart_pc.un1_state_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_RNI9ADK1_4_LC_14_8_7 .C_ON=1'b0;
    defparam \uart_drone.state_RNI9ADK1_4_LC_14_8_7 .SEQ_MODE=4'b0000;
    defparam \uart_drone.state_RNI9ADK1_4_LC_14_8_7 .LUT_INIT=16'b1011111110101010;
    LogicCell40 \uart_drone.state_RNI9ADK1_4_LC_14_8_7  (
            .in0(N__36476),
            .in1(N__31448),
            .in2(N__33525),
            .in3(N__44539),
            .lcout(\uart_drone.un1_state_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_RNO_0_2_LC_14_9_1 .C_ON=1'b0;
    defparam \uart_drone.state_RNO_0_2_LC_14_9_1 .SEQ_MODE=4'b0000;
    defparam \uart_drone.state_RNO_0_2_LC_14_9_1 .LUT_INIT=16'b0000000000111010;
    LogicCell40 \uart_drone.state_RNO_0_2_LC_14_9_1  (
            .in0(N__33750),
            .in1(N__31392),
            .in2(N__31302),
            .in3(N__44077),
            .lcout(),
            .ltout(\uart_drone.state_srsts_i_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_2_LC_14_9_2 .C_ON=1'b0;
    defparam \uart_drone.state_2_LC_14_9_2 .SEQ_MODE=4'b1000;
    defparam \uart_drone.state_2_LC_14_9_2 .LUT_INIT=16'b1111000001110000;
    LogicCell40 \uart_drone.state_2_LC_14_9_2  (
            .in0(N__36537),
            .in1(N__36607),
            .in2(N__31305),
            .in3(N__31300),
            .lcout(\uart_drone.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47404),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_RNIOU0N_4_LC_14_9_4 .C_ON=1'b0;
    defparam \uart_drone.state_RNIOU0N_4_LC_14_9_4 .SEQ_MODE=4'b0000;
    defparam \uart_drone.state_RNIOU0N_4_LC_14_9_4 .LUT_INIT=16'b1010101010111011;
    LogicCell40 \uart_drone.state_RNIOU0N_4_LC_14_9_4  (
            .in0(N__44076),
            .in1(N__36484),
            .in2(_gnd_net_),
            .in3(N__44541),
            .lcout(\uart_drone.state_RNIOU0NZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.bit_Count_0_LC_14_10_0 .C_ON=1'b0;
    defparam \uart_pc.bit_Count_0_LC_14_10_0 .SEQ_MODE=4'b1000;
    defparam \uart_pc.bit_Count_0_LC_14_10_0 .LUT_INIT=16'b0000001011110000;
    LogicCell40 \uart_pc.bit_Count_0_LC_14_10_0  (
            .in0(N__31725),
            .in1(N__31768),
            .in2(N__32130),
            .in3(N__31748),
            .lcout(\uart_pc.bit_CountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47388),
            .ce(),
            .sr(N__43830));
    defparam \uart_pc.bit_Count_RNO_0_2_LC_14_10_1 .C_ON=1'b0;
    defparam \uart_pc.bit_Count_RNO_0_2_LC_14_10_1 .SEQ_MODE=4'b0000;
    defparam \uart_pc.bit_Count_RNO_0_2_LC_14_10_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uart_pc.bit_Count_RNO_0_2_LC_14_10_1  (
            .in0(N__31747),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32125),
            .lcout(),
            .ltout(\uart_pc.CO0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.bit_Count_2_LC_14_10_2 .C_ON=1'b0;
    defparam \uart_pc.bit_Count_2_LC_14_10_2 .SEQ_MODE=4'b1000;
    defparam \uart_pc.bit_Count_2_LC_14_10_2 .LUT_INIT=16'b0001010001000100;
    LogicCell40 \uart_pc.bit_Count_2_LC_14_10_2  (
            .in0(N__31671),
            .in1(N__32033),
            .in2(N__31854),
            .in3(N__32080),
            .lcout(\uart_pc.bit_CountZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47388),
            .ce(),
            .sr(N__43830));
    defparam \uart_pc.bit_Count_1_LC_14_10_3 .C_ON=1'b0;
    defparam \uart_pc.bit_Count_1_LC_14_10_3 .SEQ_MODE=4'b1000;
    defparam \uart_pc.bit_Count_1_LC_14_10_3 .LUT_INIT=16'b0000000001111000;
    LogicCell40 \uart_pc.bit_Count_1_LC_14_10_3  (
            .in0(N__31749),
            .in1(N__32129),
            .in2(N__32082),
            .in3(N__31670),
            .lcout(\uart_pc.bit_CountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47388),
            .ce(),
            .sr(N__43830));
    defparam \Commands_frame_decoder.state_RNIBV7S_2_LC_14_10_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIBV7S_2_LC_14_10_7 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIBV7S_2_LC_14_10_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \Commands_frame_decoder.state_RNIBV7S_2_LC_14_10_7  (
            .in0(_gnd_net_),
            .in1(N__31828),
            .in2(_gnd_net_),
            .in3(N__44070),
            .lcout(\Commands_frame_decoder.un1_sink_data_valid_2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI5QE01_0_LC_14_11_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI5QE01_0_LC_14_11_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI5QE01_0_LC_14_11_2 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI5QE01_0_LC_14_11_2  (
            .in0(N__33998),
            .in1(N__40408),
            .in2(N__33981),
            .in3(N__41815),
            .lcout(\ppm_encoder_1.init_pulses_1_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.bit_Count_RNI4U6E1_2_LC_14_11_3 .C_ON=1'b0;
    defparam \uart_pc.bit_Count_RNI4U6E1_2_LC_14_11_3 .SEQ_MODE=4'b0000;
    defparam \uart_pc.bit_Count_RNI4U6E1_2_LC_14_11_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uart_pc.bit_Count_RNI4U6E1_2_LC_14_11_3  (
            .in0(N__32023),
            .in1(N__32117),
            .in2(_gnd_net_),
            .in3(N__32067),
            .lcout(\uart_pc.N_152 ),
            .ltout(\uart_pc.N_152_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_RNIUPE73_3_LC_14_11_4 .C_ON=1'b0;
    defparam \uart_pc.state_RNIUPE73_3_LC_14_11_4 .SEQ_MODE=4'b0000;
    defparam \uart_pc.state_RNIUPE73_3_LC_14_11_4 .LUT_INIT=16'b1100000011001100;
    LogicCell40 \uart_pc.state_RNIUPE73_3_LC_14_11_4  (
            .in0(_gnd_net_),
            .in1(N__31746),
            .in2(N__31728),
            .in3(N__31724),
            .lcout(\uart_pc.un1_state_7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.PPM_STATE_RNI2APU1_2_1_LC_14_11_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_RNI2APU1_2_1_LC_14_11_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.PPM_STATE_RNI2APU1_2_1_LC_14_11_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ppm_encoder_1.PPM_STATE_RNI2APU1_2_1_LC_14_11_5  (
            .in0(N__41816),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37686),
            .lcout(\ppm_encoder_1.PPM_STATE_RNI2APU1_2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_Aux_RNO_0_6_LC_14_11_6 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_RNO_0_6_LC_14_11_6 .SEQ_MODE=4'b0000;
    defparam \uart_pc.data_Aux_RNO_0_6_LC_14_11_6 .LUT_INIT=16'b0101000000000000;
    LogicCell40 \uart_pc.data_Aux_RNO_0_6_LC_14_11_6  (
            .in0(N__32118),
            .in1(_gnd_net_),
            .in2(N__32081),
            .in3(N__32024),
            .lcout(\uart_pc.data_Auxce_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNIAIVN2_7_LC_14_12_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNIAIVN2_7_LC_14_12_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNIAIVN2_7_LC_14_12_0 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \ppm_encoder_1.elevator_RNIAIVN2_7_LC_14_12_0  (
            .in0(N__31969),
            .in1(N__35784),
            .in2(N__31920),
            .in3(N__35697),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_1_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIJII96_7_LC_14_12_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIJII96_7_LC_14_12_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIJII96_7_LC_14_12_1 .LUT_INIT=16'b0011111100111111;
    LogicCell40 \ppm_encoder_1.throttle_RNIJII96_7_LC_14_12_1  (
            .in0(_gnd_net_),
            .in1(N__35319),
            .in2(N__31980),
            .in3(N__40251),
            .lcout(\ppm_encoder_1.throttle_RNIJII96Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_7_LC_14_12_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_7_LC_14_12_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_7_LC_14_12_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_7_LC_14_12_3  (
            .in0(N__40135),
            .in1(N__35338),
            .in2(_gnd_net_),
            .in3(N__31918),
            .lcout(),
            .ltout(\ppm_encoder_1.N_299_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_7_LC_14_12_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_7_LC_14_12_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_7_LC_14_12_4 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_7_LC_14_12_4  (
            .in0(N__31970),
            .in1(_gnd_net_),
            .in2(N__31977),
            .in3(N__38925),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_7_LC_14_12_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_7_LC_14_12_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.aileron_7_LC_14_12_5 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \ppm_encoder_1.aileron_7_LC_14_12_5  (
            .in0(N__35568),
            .in1(N__35582),
            .in2(N__31974),
            .in3(N__37089),
            .lcout(\ppm_encoder_1.aileronZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47364),
            .ce(),
            .sr(N__43848));
    defparam \ppm_encoder_1.elevator_7_LC_14_12_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_7_LC_14_12_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.elevator_7_LC_14_12_6 .LUT_INIT=16'b0011101011001010;
    LogicCell40 \ppm_encoder_1.elevator_7_LC_14_12_6  (
            .in0(N__31919),
            .in1(N__31956),
            .in2(N__37147),
            .in3(N__31944),
            .lcout(\ppm_encoder_1.elevatorZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47364),
            .ce(),
            .sr(N__43848));
    defparam \ppm_encoder_1.throttle_7_LC_14_12_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_7_LC_14_12_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_7_LC_14_12_7 .LUT_INIT=16'b0101101011001100;
    LogicCell40 \ppm_encoder_1.throttle_7_LC_14_12_7  (
            .in0(N__31905),
            .in1(N__35339),
            .in2(N__31899),
            .in3(N__37090),
            .lcout(\ppm_encoder_1.throttleZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47364),
            .ce(),
            .sr(N__43848));
    defparam \scaler_2.un2_source_data_0_cry_1_c_LC_14_13_0 .C_ON=1'b1;
    defparam \scaler_2.un2_source_data_0_cry_1_c_LC_14_13_0 .SEQ_MODE=4'b0000;
    defparam \scaler_2.un2_source_data_0_cry_1_c_LC_14_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \scaler_2.un2_source_data_0_cry_1_c_LC_14_13_0  (
            .in0(_gnd_net_),
            .in1(N__32285),
            .in2(N__32301),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_13_0_),
            .carryout(\scaler_2.un2_source_data_0_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_2.source_data_1_esr_6_LC_14_13_1 .C_ON=1'b1;
    defparam \scaler_2.source_data_1_esr_6_LC_14_13_1 .SEQ_MODE=4'b1000;
    defparam \scaler_2.source_data_1_esr_6_LC_14_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_2.source_data_1_esr_6_LC_14_13_1  (
            .in0(_gnd_net_),
            .in1(N__32252),
            .in2(N__32289),
            .in3(N__32259),
            .lcout(scaler_2_data_6),
            .ltout(),
            .carryin(\scaler_2.un2_source_data_0_cry_1 ),
            .carryout(\scaler_2.un2_source_data_0_cry_2 ),
            .clk(N__47349),
            .ce(N__32405),
            .sr(N__43854));
    defparam \scaler_2.source_data_1_esr_7_LC_14_13_2 .C_ON=1'b1;
    defparam \scaler_2.source_data_1_esr_7_LC_14_13_2 .SEQ_MODE=4'b1000;
    defparam \scaler_2.source_data_1_esr_7_LC_14_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_2.source_data_1_esr_7_LC_14_13_2  (
            .in0(_gnd_net_),
            .in1(N__32231),
            .in2(N__32256),
            .in3(N__32238),
            .lcout(scaler_2_data_7),
            .ltout(),
            .carryin(\scaler_2.un2_source_data_0_cry_2 ),
            .carryout(\scaler_2.un2_source_data_0_cry_3 ),
            .clk(N__47349),
            .ce(N__32405),
            .sr(N__43854));
    defparam \scaler_2.source_data_1_esr_8_LC_14_13_3 .C_ON=1'b1;
    defparam \scaler_2.source_data_1_esr_8_LC_14_13_3 .SEQ_MODE=4'b1000;
    defparam \scaler_2.source_data_1_esr_8_LC_14_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_2.source_data_1_esr_8_LC_14_13_3  (
            .in0(_gnd_net_),
            .in1(N__32210),
            .in2(N__32235),
            .in3(N__32217),
            .lcout(scaler_2_data_8),
            .ltout(),
            .carryin(\scaler_2.un2_source_data_0_cry_3 ),
            .carryout(\scaler_2.un2_source_data_0_cry_4 ),
            .clk(N__47349),
            .ce(N__32405),
            .sr(N__43854));
    defparam \scaler_2.source_data_1_esr_9_LC_14_13_4 .C_ON=1'b1;
    defparam \scaler_2.source_data_1_esr_9_LC_14_13_4 .SEQ_MODE=4'b1000;
    defparam \scaler_2.source_data_1_esr_9_LC_14_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_2.source_data_1_esr_9_LC_14_13_4  (
            .in0(_gnd_net_),
            .in1(N__32189),
            .in2(N__32214),
            .in3(N__32196),
            .lcout(scaler_2_data_9),
            .ltout(),
            .carryin(\scaler_2.un2_source_data_0_cry_4 ),
            .carryout(\scaler_2.un2_source_data_0_cry_5 ),
            .clk(N__47349),
            .ce(N__32405),
            .sr(N__43854));
    defparam \scaler_2.source_data_1_esr_10_LC_14_13_5 .C_ON=1'b1;
    defparam \scaler_2.source_data_1_esr_10_LC_14_13_5 .SEQ_MODE=4'b1000;
    defparam \scaler_2.source_data_1_esr_10_LC_14_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_2.source_data_1_esr_10_LC_14_13_5  (
            .in0(_gnd_net_),
            .in1(N__32168),
            .in2(N__32193),
            .in3(N__32175),
            .lcout(scaler_2_data_10),
            .ltout(),
            .carryin(\scaler_2.un2_source_data_0_cry_5 ),
            .carryout(\scaler_2.un2_source_data_0_cry_6 ),
            .clk(N__47349),
            .ce(N__32405),
            .sr(N__43854));
    defparam \scaler_2.source_data_1_esr_11_LC_14_13_6 .C_ON=1'b1;
    defparam \scaler_2.source_data_1_esr_11_LC_14_13_6 .SEQ_MODE=4'b1000;
    defparam \scaler_2.source_data_1_esr_11_LC_14_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_2.source_data_1_esr_11_LC_14_13_6  (
            .in0(_gnd_net_),
            .in1(N__32147),
            .in2(N__32172),
            .in3(N__32154),
            .lcout(scaler_2_data_11),
            .ltout(),
            .carryin(\scaler_2.un2_source_data_0_cry_6 ),
            .carryout(\scaler_2.un2_source_data_0_cry_7 ),
            .clk(N__47349),
            .ce(N__32405),
            .sr(N__43854));
    defparam \scaler_2.source_data_1_esr_12_LC_14_13_7 .C_ON=1'b1;
    defparam \scaler_2.source_data_1_esr_12_LC_14_13_7 .SEQ_MODE=4'b1000;
    defparam \scaler_2.source_data_1_esr_12_LC_14_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_2.source_data_1_esr_12_LC_14_13_7  (
            .in0(_gnd_net_),
            .in1(N__32450),
            .in2(N__32151),
            .in3(N__32133),
            .lcout(scaler_2_data_12),
            .ltout(),
            .carryin(\scaler_2.un2_source_data_0_cry_7 ),
            .carryout(\scaler_2.un2_source_data_0_cry_8 ),
            .clk(N__47349),
            .ce(N__32405),
            .sr(N__43854));
    defparam \scaler_2.source_data_1_esr_13_LC_14_14_0 .C_ON=1'b1;
    defparam \scaler_2.source_data_1_esr_13_LC_14_14_0 .SEQ_MODE=4'b1000;
    defparam \scaler_2.source_data_1_esr_13_LC_14_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_2.source_data_1_esr_13_LC_14_14_0  (
            .in0(_gnd_net_),
            .in1(N__32451),
            .in2(N__32427),
            .in3(N__32412),
            .lcout(scaler_2_data_13),
            .ltout(),
            .carryin(bfn_14_14_0_),
            .carryout(\scaler_2.un2_source_data_0_cry_9 ),
            .clk(N__47332),
            .ce(N__32404),
            .sr(N__43860));
    defparam \scaler_2.source_data_1_esr_14_LC_14_14_1 .C_ON=1'b0;
    defparam \scaler_2.source_data_1_esr_14_LC_14_14_1 .SEQ_MODE=4'b1000;
    defparam \scaler_2.source_data_1_esr_14_LC_14_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \scaler_2.source_data_1_esr_14_LC_14_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32409),
            .lcout(scaler_2_data_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47332),
            .ce(N__32404),
            .sr(N__43860));
    defparam \ppm_encoder_1.throttle_RNIU7KK2_9_LC_14_15_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIU7KK2_9_LC_14_15_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIU7KK2_9_LC_14_15_0 .LUT_INIT=16'b1011000010111011;
    LogicCell40 \ppm_encoder_1.throttle_RNIU7KK2_9_LC_14_15_0  (
            .in0(N__40531),
            .in1(N__35286),
            .in2(N__32571),
            .in3(N__37581),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNITSI96_9_LC_14_15_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNITSI96_9_LC_14_15_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNITSI96_9_LC_14_15_1 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ppm_encoder_1.throttle_RNITSI96_9_LC_14_15_1  (
            .in0(N__40574),
            .in1(_gnd_net_),
            .in2(N__32379),
            .in3(N__32376),
            .lcout(\ppm_encoder_1.throttle_RNITSI96Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNIEMVN2_9_LC_14_15_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNIEMVN2_9_LC_14_15_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNIEMVN2_9_LC_14_15_2 .LUT_INIT=16'b1100010011110101;
    LogicCell40 \ppm_encoder_1.elevator_RNIEMVN2_9_LC_14_15_2  (
            .in0(N__35801),
            .in1(N__32365),
            .in2(N__32316),
            .in3(N__35731),
            .lcout(\ppm_encoder_1.un2_throttle_iv_1_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_9_LC_14_15_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_9_LC_14_15_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_9_LC_14_15_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_9_LC_14_15_3  (
            .in0(N__40127),
            .in1(N__32569),
            .in2(_gnd_net_),
            .in3(N__32314),
            .lcout(),
            .ltout(\ppm_encoder_1.N_301_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_9_LC_14_15_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_9_LC_14_15_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_9_LC_14_15_4 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_9_LC_14_15_4  (
            .in0(N__38945),
            .in1(_gnd_net_),
            .in2(N__32370),
            .in3(N__32366),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_9_LC_14_15_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_9_LC_14_15_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.aileron_9_LC_14_15_5 .LUT_INIT=16'b0011101011001010;
    LogicCell40 \ppm_encoder_1.aileron_9_LC_14_15_5  (
            .in0(N__32367),
            .in1(N__36014),
            .in2(N__37242),
            .in3(N__35997),
            .lcout(\ppm_encoder_1.aileronZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47319),
            .ce(),
            .sr(N__43869));
    defparam \ppm_encoder_1.elevator_9_LC_14_15_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_9_LC_14_15_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.elevator_9_LC_14_15_6 .LUT_INIT=16'b0010111011100010;
    LogicCell40 \ppm_encoder_1.elevator_9_LC_14_15_6  (
            .in0(N__32315),
            .in1(N__37193),
            .in2(N__32355),
            .in3(N__32328),
            .lcout(\ppm_encoder_1.elevatorZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47319),
            .ce(),
            .sr(N__43869));
    defparam \ppm_encoder_1.throttle_9_LC_14_15_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_9_LC_14_15_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_9_LC_14_15_7 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.throttle_9_LC_14_15_7  (
            .in0(N__32595),
            .in1(N__32577),
            .in2(N__37243),
            .in3(N__32570),
            .lcout(\ppm_encoder_1.throttleZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47319),
            .ce(),
            .sr(N__43869));
    defparam \ppm_encoder_1.throttle_RNII6JI2_12_LC_14_16_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNII6JI2_12_LC_14_16_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNII6JI2_12_LC_14_16_0 .LUT_INIT=16'b0001001101011111;
    LogicCell40 \ppm_encoder_1.throttle_RNII6JI2_12_LC_14_16_0  (
            .in0(N__37582),
            .in1(N__32635),
            .in2(N__34064),
            .in3(N__35288),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNIFQRT5_12_LC_14_16_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNIFQRT5_12_LC_14_16_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNIFQRT5_12_LC_14_16_1 .LUT_INIT=16'b0000111111111111;
    LogicCell40 \ppm_encoder_1.elevator_RNIFQRT5_12_LC_14_16_1  (
            .in0(N__38096),
            .in1(_gnd_net_),
            .in2(N__32556),
            .in3(N__32553),
            .lcout(\ppm_encoder_1.elevator_RNIFQRT5Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNI25DH2_12_LC_14_16_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNI25DH2_12_LC_14_16_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNI25DH2_12_LC_14_16_2 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \ppm_encoder_1.elevator_RNI25DH2_12_LC_14_16_2  (
            .in0(N__32542),
            .in1(N__35818),
            .in2(N__34040),
            .in3(N__35733),
            .lcout(\ppm_encoder_1.un2_throttle_iv_1_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_12_LC_14_16_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_12_LC_14_16_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_12_LC_14_16_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_12_LC_14_16_4  (
            .in0(N__32543),
            .in1(N__38983),
            .in2(_gnd_net_),
            .in3(N__34020),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_12_LC_14_16_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_12_LC_14_16_5 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.aileron_12_LC_14_16_5 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \ppm_encoder_1.aileron_12_LC_14_16_5  (
            .in0(N__35946),
            .in1(N__35922),
            .in2(N__32547),
            .in3(N__37191),
            .lcout(\ppm_encoder_1.aileronZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47309),
            .ce(),
            .sr(N__43876));
    defparam \ppm_encoder_1.elevator_12_LC_14_16_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_12_LC_14_16_6 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.elevator_12_LC_14_16_6 .LUT_INIT=16'b0011101011001010;
    LogicCell40 \ppm_encoder_1.elevator_12_LC_14_16_6  (
            .in0(N__34036),
            .in1(N__32529),
            .in2(N__37241),
            .in3(N__32505),
            .lcout(\ppm_encoder_1.elevatorZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47309),
            .ce(),
            .sr(N__43876));
    defparam \ppm_encoder_1.throttle_12_LC_14_16_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_12_LC_14_16_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_12_LC_14_16_7 .LUT_INIT=16'b0111101101001000;
    LogicCell40 \ppm_encoder_1.throttle_12_LC_14_16_7  (
            .in0(N__32493),
            .in1(N__37192),
            .in2(N__32463),
            .in3(N__34060),
            .lcout(\ppm_encoder_1.throttleZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47309),
            .ce(),
            .sr(N__43876));
    defparam \ppm_encoder_1.throttle_RNIG4JI2_11_LC_14_17_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIG4JI2_11_LC_14_17_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIG4JI2_11_LC_14_17_0 .LUT_INIT=16'b0000011101110111;
    LogicCell40 \ppm_encoder_1.throttle_RNIG4JI2_11_LC_14_17_0  (
            .in0(N__34600),
            .in1(N__35287),
            .in2(N__34632),
            .in3(N__37591),
            .lcout(\ppm_encoder_1.un2_throttle_iv_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.rudder_11_LC_14_17_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_11_LC_14_17_1 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.rudder_11_LC_14_17_1 .LUT_INIT=16'b0111001011011000;
    LogicCell40 \ppm_encoder_1.rudder_11_LC_14_17_1  (
            .in0(N__37233),
            .in1(N__32754),
            .in2(N__34605),
            .in3(N__32748),
            .lcout(\ppm_encoder_1.rudderZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47299),
            .ce(),
            .sr(N__43883));
    defparam \ppm_encoder_1.throttle_11_LC_14_17_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_11_LC_14_17_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_11_LC_14_17_2 .LUT_INIT=16'b0010111011100010;
    LogicCell40 \ppm_encoder_1.throttle_11_LC_14_17_2  (
            .in0(N__34630),
            .in1(N__37232),
            .in2(N__32730),
            .in3(N__32706),
            .lcout(\ppm_encoder_1.throttleZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47299),
            .ce(),
            .sr(N__43883));
    defparam \ppm_encoder_1.elevator_11_LC_14_17_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_11_LC_14_17_4 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.elevator_11_LC_14_17_4 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \ppm_encoder_1.elevator_11_LC_14_17_4  (
            .in0(N__32697),
            .in1(N__32673),
            .in2(N__34928),
            .in3(N__37231),
            .lcout(\ppm_encoder_1.elevatorZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47299),
            .ce(),
            .sr(N__43883));
    defparam \ppm_encoder_1.rudder_12_LC_14_17_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_12_LC_14_17_5 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.rudder_12_LC_14_17_5 .LUT_INIT=16'b0011101011001010;
    LogicCell40 \ppm_encoder_1.rudder_12_LC_14_17_5  (
            .in0(N__32637),
            .in1(N__32661),
            .in2(N__37258),
            .in3(N__32643),
            .lcout(\ppm_encoder_1.rudderZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47299),
            .ce(),
            .sr(N__43883));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_12_LC_14_17_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_12_LC_14_17_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_12_LC_14_17_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_12_LC_14_17_6  (
            .in0(N__40928),
            .in1(N__37740),
            .in2(_gnd_net_),
            .in3(N__32636),
            .lcout(),
            .ltout(\ppm_encoder_1.N_320_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_12_LC_14_17_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_12_LC_14_17_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_12_LC_14_17_7 .LUT_INIT=16'b1010000011110101;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_12_LC_14_17_7  (
            .in0(N__41141),
            .in1(_gnd_net_),
            .in2(N__32622),
            .in3(N__35532),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNIU0DH2_10_LC_14_18_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNIU0DH2_10_LC_14_18_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNIU0DH2_10_LC_14_18_0 .LUT_INIT=16'b1010001011110011;
    LogicCell40 \ppm_encoder_1.elevator_RNIU0DH2_10_LC_14_18_0  (
            .in0(N__34735),
            .in1(N__35814),
            .in2(N__32982),
            .in3(N__35732),
            .lcout(\ppm_encoder_1.un2_throttle_iv_1_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIE2JI2_10_LC_14_18_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIE2JI2_10_LC_14_18_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIE2JI2_10_LC_14_18_2 .LUT_INIT=16'b1011000010111011;
    LogicCell40 \ppm_encoder_1.throttle_RNIE2JI2_10_LC_14_18_2  (
            .in0(N__35848),
            .in1(N__35285),
            .in2(N__32619),
            .in3(N__37590),
            .lcout(\ppm_encoder_1.un2_throttle_iv_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_10_LC_14_18_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_10_LC_14_18_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_10_LC_14_18_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_10_LC_14_18_3  (
            .in0(N__40128),
            .in1(N__32617),
            .in2(_gnd_net_),
            .in3(N__32980),
            .lcout(\ppm_encoder_1.N_302 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_10_LC_14_18_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_10_LC_14_18_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.elevator_10_LC_14_18_4 .LUT_INIT=16'b0011101011001010;
    LogicCell40 \ppm_encoder_1.elevator_10_LC_14_18_4  (
            .in0(N__32981),
            .in1(N__33015),
            .in2(N__37260),
            .in3(N__32988),
            .lcout(\ppm_encoder_1.elevatorZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47291),
            .ce(),
            .sr(N__43886));
    defparam \ppm_encoder_1.aileron_10_LC_14_18_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_10_LC_14_18_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.aileron_10_LC_14_18_6 .LUT_INIT=16'b0011101011001010;
    LogicCell40 \ppm_encoder_1.aileron_10_LC_14_18_6  (
            .in0(N__34736),
            .in1(N__35985),
            .in2(N__37259),
            .in3(N__35964),
            .lcout(\ppm_encoder_1.aileronZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47291),
            .ce(),
            .sr(N__43886));
    defparam \ppm_encoder_1.rudder_10_LC_14_18_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_10_LC_14_18_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.rudder_10_LC_14_18_7 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \ppm_encoder_1.rudder_10_LC_14_18_7  (
            .in0(N__32967),
            .in1(N__32949),
            .in2(N__35858),
            .in3(N__37240),
            .lcout(\ppm_encoder_1.rudderZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47291),
            .ce(),
            .sr(N__43886));
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNIGCO83_LC_14_19_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNIGCO83_LC_14_19_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNIGCO83_LC_14_19_0 .LUT_INIT=16'b1111110011111110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_57_c_RNIGCO83_LC_14_19_0  (
            .in0(N__40300),
            .in1(N__34711),
            .in2(N__32943),
            .in3(N__44665),
            .lcout(\ppm_encoder_1.counter24_0_I_57_c_RNIGCOZ0Z83 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.PPM_STATE_RNIV4V5_1_LC_14_19_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_RNIV4V5_1_LC_14_19_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.PPM_STATE_RNIV4V5_1_LC_14_19_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \ppm_encoder_1.PPM_STATE_RNIV4V5_1_LC_14_19_1  (
            .in0(_gnd_net_),
            .in1(N__34671),
            .in2(_gnd_net_),
            .in3(N__40299),
            .lcout(\ppm_encoder_1.PPM_STATE_59_d ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.PPM_STATE_0_LC_14_19_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_0_LC_14_19_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.PPM_STATE_0_LC_14_19_2 .LUT_INIT=16'b1100111011001100;
    LogicCell40 \ppm_encoder_1.PPM_STATE_0_LC_14_19_2  (
            .in0(N__40301),
            .in1(N__34712),
            .in2(N__34679),
            .in3(N__44666),
            .lcout(\ppm_encoder_1.PPM_STATEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47285),
            .ce(),
            .sr(N__43891));
    defparam \ppm_encoder_1.PPM_STATE_1_LC_14_19_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_1_LC_14_19_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.PPM_STATE_1_LC_14_19_4 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \ppm_encoder_1.PPM_STATE_1_LC_14_19_4  (
            .in0(N__40302),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34713),
            .lcout(\ppm_encoder_1.PPM_STATEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47285),
            .ce(),
            .sr(N__43891));
    defparam \ppm_encoder_1.ppm_output_reg_RNO_1_LC_14_19_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.ppm_output_reg_RNO_1_LC_14_19_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.ppm_output_reg_RNO_1_LC_14_19_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \ppm_encoder_1.ppm_output_reg_RNO_1_LC_14_19_7  (
            .in0(N__34893),
            .in1(N__34722),
            .in2(N__34701),
            .in3(N__39642),
            .lcout(\ppm_encoder_1.N_145 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_esr_13_LC_14_20_0 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_esr_13_LC_14_20_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_esr_13_LC_14_20_0 .LUT_INIT=16'b1100110011011101;
    LogicCell40 \pid_alt.error_i_acumm_esr_13_LC_14_20_0  (
            .in0(N__32856),
            .in1(N__32826),
            .in2(_gnd_net_),
            .in3(N__32799),
            .lcout(\pid_alt.error_i_acummZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47276),
            .ce(N__32775),
            .sr(N__33719));
    defparam \ppm_encoder_1.init_pulses_RNIQDRP_0_11_LC_14_20_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIQDRP_0_11_LC_14_20_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIQDRP_0_11_LC_14_20_2 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIQDRP_0_11_LC_14_20_2  (
            .in0(N__41771),
            .in1(N__42276),
            .in2(_gnd_net_),
            .in3(N__37764),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIQDRP_11_LC_14_20_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIQDRP_11_LC_14_20_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIQDRP_11_LC_14_20_3 .LUT_INIT=16'b0101101010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIQDRP_11_LC_14_20_3  (
            .in0(N__37763),
            .in1(_gnd_net_),
            .in2(N__42291),
            .in3(N__41775),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIRERP_0_12_LC_14_20_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIRERP_0_12_LC_14_20_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIRERP_0_12_LC_14_20_4 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIRERP_0_12_LC_14_20_4  (
            .in0(N__41772),
            .in1(N__42277),
            .in2(_gnd_net_),
            .in3(N__37739),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIRERP_12_LC_14_20_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIRERP_12_LC_14_20_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIRERP_12_LC_14_20_5 .LUT_INIT=16'b0101101010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIRERP_12_LC_14_20_5  (
            .in0(N__37738),
            .in1(_gnd_net_),
            .in2(N__42290),
            .in3(N__41774),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.PPM_STATE_RNIV4V5_0_1_LC_14_20_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_RNIV4V5_0_1_LC_14_20_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.PPM_STATE_RNIV4V5_0_1_LC_14_20_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \ppm_encoder_1.PPM_STATE_RNIV4V5_0_1_LC_14_20_6  (
            .in0(N__41773),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\ppm_encoder_1.N_1330_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.PPM_STATE_RNI2APU1_0_1_LC_14_20_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_RNI2APU1_0_1_LC_14_20_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.PPM_STATE_RNI2APU1_0_1_LC_14_20_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ppm_encoder_1.PPM_STATE_RNI2APU1_0_1_LC_14_20_7  (
            .in0(_gnd_net_),
            .in1(N__37712),
            .in2(_gnd_net_),
            .in3(N__41770),
            .lcout(\ppm_encoder_1.PPM_STATE_RNI2APU1_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_ki_6_LC_14_21_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_ki_6_LC_14_21_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_ki_6_LC_14_21_5 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_ki_6_LC_14_21_5  (
            .in0(_gnd_net_),
            .in1(N__33440),
            .in2(_gnd_net_),
            .in3(N__46681),
            .lcout(alt_ki_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47273),
            .ce(N__44828),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_6_LC_14_22_3 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_6_LC_14_22_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_6_LC_14_22_3 .LUT_INIT=16'b1100101011111010;
    LogicCell40 \pid_alt.error_i_acumm_6_LC_14_22_3  (
            .in0(N__33260),
            .in1(N__33282),
            .in2(N__33246),
            .in3(N__33078),
            .lcout(\pid_alt.error_i_acummZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47269),
            .ce(),
            .sr(N__33720));
    defparam \pid_alt.error_i_acumm_11_LC_14_22_7 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_11_LC_14_22_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_11_LC_14_22_7 .LUT_INIT=16'b1110010011101110;
    LogicCell40 \pid_alt.error_i_acumm_11_LC_14_22_7  (
            .in0(N__33240),
            .in1(N__33027),
            .in2(N__33105),
            .in3(N__33077),
            .lcout(\pid_alt.error_i_acummZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47269),
            .ce(),
            .sr(N__33720));
    defparam \pid_alt.error_i_acumm_prereg_esr_0_LC_14_23_5 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_0_LC_14_23_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_0_LC_14_23_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_0_LC_14_23_5  (
            .in0(_gnd_net_),
            .in1(N__39581),
            .in2(_gnd_net_),
            .in3(N__33672),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47266),
            .ce(N__33627),
            .sr(N__43899));
    defparam \uart_drone.timer_Count_RNI5A9J_1_LC_15_6_0 .C_ON=1'b1;
    defparam \uart_drone.timer_Count_RNI5A9J_1_LC_15_6_0 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNI5A9J_1_LC_15_6_0 .LUT_INIT=16'b0001000100010001;
    LogicCell40 \uart_drone.timer_Count_RNI5A9J_1_LC_15_6_0  (
            .in0(N__33954),
            .in1(N__33929),
            .in2(N__33957),
            .in3(_gnd_net_),
            .lcout(\uart_drone.un1_state_2_0_a3_0 ),
            .ltout(),
            .carryin(bfn_15_6_0_),
            .carryout(\uart_drone.un4_timer_Count_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_RNO_0_2_LC_15_6_1 .C_ON=1'b1;
    defparam \uart_drone.timer_Count_RNO_0_2_LC_15_6_1 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNO_0_2_LC_15_6_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_drone.timer_Count_RNO_0_2_LC_15_6_1  (
            .in0(_gnd_net_),
            .in1(N__33509),
            .in2(_gnd_net_),
            .in3(N__33483),
            .lcout(\uart_drone.timer_Count_RNO_0_0_2 ),
            .ltout(),
            .carryin(\uart_drone.un4_timer_Count_1_cry_1 ),
            .carryout(\uart_drone.un4_timer_Count_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_RNO_0_3_LC_15_6_2 .C_ON=1'b1;
    defparam \uart_drone.timer_Count_RNO_0_3_LC_15_6_2 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNO_0_3_LC_15_6_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_drone.timer_Count_RNO_0_3_LC_15_6_2  (
            .in0(_gnd_net_),
            .in1(N__36544),
            .in2(_gnd_net_),
            .in3(N__33468),
            .lcout(\uart_drone.timer_Count_RNO_0_0_3 ),
            .ltout(),
            .carryin(\uart_drone.un4_timer_Count_1_cry_2 ),
            .carryout(\uart_drone.un4_timer_Count_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_RNO_0_4_LC_15_6_3 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_RNO_0_4_LC_15_6_3 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNO_0_4_LC_15_6_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uart_drone.timer_Count_RNO_0_4_LC_15_6_3  (
            .in0(_gnd_net_),
            .in1(N__36615),
            .in2(_gnd_net_),
            .in3(N__33465),
            .lcout(\uart_drone.timer_Count_RNO_0_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_0_LC_15_6_7 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_0_LC_15_6_7 .SEQ_MODE=4'b1000;
    defparam \uart_drone.timer_Count_0_LC_15_6_7 .LUT_INIT=16'b0000000001010100;
    LogicCell40 \uart_drone.timer_Count_0_LC_15_6_7  (
            .in0(N__33956),
            .in1(N__33914),
            .in2(N__33884),
            .in3(N__44122),
            .lcout(\uart_drone.timer_CountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47442),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_2_LC_15_7_1 .C_ON=1'b0;
    defparam \reset_module_System.count_2_LC_15_7_1 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_2_LC_15_7_1 .LUT_INIT=16'b0100110011001100;
    LogicCell40 \reset_module_System.count_2_LC_15_7_1  (
            .in0(N__37317),
            .in1(N__34779),
            .in2(N__33841),
            .in3(N__33787),
            .lcout(\reset_module_System.countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47436),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNI97FD_5_LC_15_7_2 .C_ON=1'b0;
    defparam \reset_module_System.count_RNI97FD_5_LC_15_7_2 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNI97FD_5_LC_15_7_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \reset_module_System.count_RNI97FD_5_LC_15_7_2  (
            .in0(N__34988),
            .in1(N__35003),
            .in2(N__34974),
            .in3(N__35033),
            .lcout(),
            .ltout(\reset_module_System.reset6_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNIA72I1_16_LC_15_7_3 .C_ON=1'b0;
    defparam \reset_module_System.count_RNIA72I1_16_LC_15_7_3 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNIA72I1_16_LC_15_7_3 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \reset_module_System.count_RNIA72I1_16_LC_15_7_3  (
            .in0(N__35105),
            .in1(N__35088),
            .in2(N__33450),
            .in3(N__33447),
            .lcout(\reset_module_System.reset6_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_RNO_0_1_LC_15_7_5 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_RNO_0_1_LC_15_7_5 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNO_0_1_LC_15_7_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart_drone.timer_Count_RNO_0_1_LC_15_7_5  (
            .in0(_gnd_net_),
            .in1(N__33955),
            .in2(_gnd_net_),
            .in3(N__33930),
            .lcout(),
            .ltout(\uart_drone.timer_Count_RNO_0_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_1_LC_15_7_6 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_1_LC_15_7_6 .SEQ_MODE=4'b1000;
    defparam \uart_drone.timer_Count_1_LC_15_7_6 .LUT_INIT=16'b0000000011100000;
    LogicCell40 \uart_drone.timer_Count_1_LC_15_7_6  (
            .in0(N__33869),
            .in1(N__33915),
            .in2(N__33933),
            .in3(N__44128),
            .lcout(\uart_drone.timer_CountZ1Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47436),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_4_LC_15_8_1 .C_ON=1'b0;
    defparam \uart_drone.state_4_LC_15_8_1 .SEQ_MODE=4'b1000;
    defparam \uart_drone.state_4_LC_15_8_1 .LUT_INIT=16'b1100110011101100;
    LogicCell40 \uart_drone.state_4_LC_15_8_1  (
            .in0(N__44538),
            .in1(N__33913),
            .in2(N__36714),
            .in3(N__44123),
            .lcout(\uart_drone.stateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47426),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_RNI40411_2_LC_15_8_3 .C_ON=1'b0;
    defparam \uart_drone.state_RNI40411_2_LC_15_8_3 .SEQ_MODE=4'b0000;
    defparam \uart_drone.state_RNI40411_2_LC_15_8_3 .LUT_INIT=16'b0011001011111010;
    LogicCell40 \uart_drone.state_RNI40411_2_LC_15_8_3  (
            .in0(N__44537),
            .in1(N__36604),
            .in2(N__33752),
            .in3(N__36535),
            .lcout(\uart_drone.timer_Count_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNI9O1P_2_LC_15_8_5 .C_ON=1'b0;
    defparam \reset_module_System.count_RNI9O1P_2_LC_15_8_5 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNI9O1P_2_LC_15_8_5 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \reset_module_System.count_RNI9O1P_2_LC_15_8_5  (
            .in0(N__35019),
            .in1(N__34770),
            .in2(N__35067),
            .in3(N__34791),
            .lcout(\reset_module_System.reset6_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNIMJ304_12_LC_15_9_0 .C_ON=1'b0;
    defparam \reset_module_System.count_RNIMJ304_12_LC_15_9_0 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNIMJ304_12_LC_15_9_0 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \reset_module_System.count_RNIMJ304_12_LC_15_9_0  (
            .in0(N__34831),
            .in1(N__34947),
            .in2(N__35145),
            .in3(N__33801),
            .lcout(\reset_module_System.reset6_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.bit_Count_RNIJOJC1_2_LC_15_9_1 .C_ON=1'b0;
    defparam \uart_drone.bit_Count_RNIJOJC1_2_LC_15_9_1 .SEQ_MODE=4'b0000;
    defparam \uart_drone.bit_Count_RNIJOJC1_2_LC_15_9_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uart_drone.bit_Count_RNIJOJC1_2_LC_15_9_1  (
            .in0(N__36671),
            .in1(N__39496),
            .in2(_gnd_net_),
            .in3(N__44391),
            .lcout(\uart_drone.N_152 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_RNO_0_3_LC_15_9_6 .C_ON=1'b0;
    defparam \uart_drone.state_RNO_0_3_LC_15_9_6 .SEQ_MODE=4'b0000;
    defparam \uart_drone.state_RNO_0_3_LC_15_9_6 .LUT_INIT=16'b0001010101010101;
    LogicCell40 \uart_drone.state_RNO_0_3_LC_15_9_6  (
            .in0(N__44540),
            .in1(N__36606),
            .in2(N__33753),
            .in3(N__36536),
            .lcout(),
            .ltout(\uart_drone.N_145_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_3_LC_15_9_7 .C_ON=1'b0;
    defparam \uart_drone.state_3_LC_15_9_7 .SEQ_MODE=4'b1000;
    defparam \uart_drone.state_3_LC_15_9_7 .LUT_INIT=16'b0000000000001011;
    LogicCell40 \uart_drone.state_3_LC_15_9_7  (
            .in0(N__33751),
            .in1(N__36710),
            .in2(N__33723),
            .in3(N__44124),
            .lcout(\uart_drone.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47416),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.data_Aux_RNO_0_2_LC_15_10_0 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_RNO_0_2_LC_15_10_0 .SEQ_MODE=4'b0000;
    defparam \uart_drone.data_Aux_RNO_0_2_LC_15_10_0 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \uart_drone.data_Aux_RNO_0_2_LC_15_10_0  (
            .in0(N__36677),
            .in1(N__39512),
            .in2(_gnd_net_),
            .in3(N__44405),
            .lcout(\uart_drone.data_Auxce_0_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.data_Aux_RNO_0_6_LC_15_10_1 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_RNO_0_6_LC_15_10_1 .SEQ_MODE=4'b0000;
    defparam \uart_drone.data_Aux_RNO_0_6_LC_15_10_1 .LUT_INIT=16'b0101000000000000;
    LogicCell40 \uart_drone.data_Aux_RNO_0_6_LC_15_10_1  (
            .in0(N__44406),
            .in1(_gnd_net_),
            .in2(N__39519),
            .in3(N__36678),
            .lcout(\uart_drone.data_Auxce_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_LC_15_10_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_LC_15_10_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_LC_15_10_5 .LUT_INIT=16'b0010001000110000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_2_LC_15_10_5  (
            .in0(N__34008),
            .in1(N__44110),
            .in2(N__40926),
            .in3(N__42009),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47405),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_3_12_LC_15_10_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_3_12_LC_15_10_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_3_12_LC_15_10_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_3_12_LC_15_10_6  (
            .in0(N__40131),
            .in1(N__34068),
            .in2(_gnd_net_),
            .in3(N__34044),
            .lcout(\ppm_encoder_1.N_304 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_0_LC_15_11_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_0_LC_15_11_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_0_LC_15_11_0 .LUT_INIT=16'b1111000111111010;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_0_LC_15_11_0  (
            .in0(N__33999),
            .in1(N__42167),
            .in2(N__44136),
            .in3(N__41947),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47389),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_1_LC_15_11_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_1_LC_15_11_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_1_LC_15_11_1 .LUT_INIT=16'b0000000001111000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_1_LC_15_11_1  (
            .in0(N__41945),
            .in1(N__38917),
            .in2(N__33980),
            .in3(N__44116),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47389),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m6_LC_15_11_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m6_LC_15_11_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m6_LC_15_11_2 .LUT_INIT=16'b0000000001101100;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m6_LC_15_11_2  (
            .in0(N__40134),
            .in1(N__40888),
            .in2(N__38946),
            .in3(N__42166),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_ns_2 ),
            .ltout(\ppm_encoder_1.CHOOSE_CHANNEL_ns_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_2_LC_15_11_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_2_LC_15_11_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_2_LC_15_11_3 .LUT_INIT=16'b0011000100100000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_2_LC_15_11_3  (
            .in0(N__41946),
            .in1(N__44112),
            .in2(N__34002),
            .in3(N__35310),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47389),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI6LFQ_0_LC_15_11_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI6LFQ_0_LC_15_11_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI6LFQ_0_LC_15_11_5 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI6LFQ_0_LC_15_11_5  (
            .in0(N__33997),
            .in1(N__35129),
            .in2(N__33979),
            .in3(N__35309),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_d_4 ),
            .ltout(\ppm_encoder_1.CHOOSE_CHANNEL_d_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI5QE01_0_0_LC_15_11_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI5QE01_0_0_LC_15_11_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI5QE01_0_0_LC_15_11_6 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI5QE01_0_0_LC_15_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__34113),
            .in3(N__41943),
            .lcout(\ppm_encoder_1.init_pulses_3_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_LC_15_11_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_LC_15_11_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_LC_15_11_7 .LUT_INIT=16'b0001001000110000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_LC_15_11_7  (
            .in0(N__41944),
            .in1(N__44111),
            .in2(N__40377),
            .in3(N__38916),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47389),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIS5KK2_8_LC_15_12_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIS5KK2_8_LC_15_12_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIS5KK2_8_LC_15_12_0 .LUT_INIT=16'b1011000010111011;
    LogicCell40 \ppm_encoder_1.throttle_RNIS5KK2_8_LC_15_12_0  (
            .in0(N__38401),
            .in1(N__35267),
            .in2(N__34188),
            .in3(N__37552),
            .lcout(\ppm_encoder_1.un2_throttle_iv_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNILS7D_3_LC_15_12_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNILS7D_3_LC_15_12_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNILS7D_3_LC_15_12_1 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNILS7D_3_LC_15_12_1  (
            .in0(N__35128),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35308),
            .lcout(\ppm_encoder_1.N_227 ),
            .ltout(\ppm_encoder_1.N_227_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1_0_LC_15_12_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1_0_LC_15_12_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1_0_LC_15_12_2 .LUT_INIT=16'b0000000000000101;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1_0_LC_15_12_2  (
            .in0(N__34100),
            .in1(_gnd_net_),
            .in2(N__34110),
            .in3(N__42114),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1Z0Z_0 ),
            .ltout(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.PPM_STATE_RNI2APU1_1_LC_15_12_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_RNI2APU1_1_LC_15_12_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.PPM_STATE_RNI2APU1_1_LC_15_12_3 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \ppm_encoder_1.PPM_STATE_RNI2APU1_1_LC_15_12_3  (
            .in0(N__42008),
            .in1(_gnd_net_),
            .in2(N__34107),
            .in3(_gnd_net_),
            .lcout(\ppm_encoder_1.PPM_STATE_RNI2APU1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_esr_RNIMGR62_4_LC_15_12_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_esr_RNIMGR62_4_LC_15_12_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.aileron_esr_RNIMGR62_4_LC_15_12_4 .LUT_INIT=16'b1100010011110101;
    LogicCell40 \ppm_encoder_1.aileron_esr_RNIMGR62_4_LC_15_12_4  (
            .in0(N__35780),
            .in1(N__34139),
            .in2(N__34166),
            .in3(N__35684),
            .lcout(\ppm_encoder_1.un2_throttle_iv_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m9_LC_15_12_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m9_LC_15_12_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m9_LC_15_12_5 .LUT_INIT=16'b0011001110000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m9_LC_15_12_5  (
            .in0(N__40136),
            .in1(N__40958),
            .in2(N__38971),
            .in3(N__39981),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_ns_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIHFK13_0_LC_15_12_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIHFK13_0_LC_15_12_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIHFK13_0_LC_15_12_6 .LUT_INIT=16'b0000000100010001;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIHFK13_0_LC_15_12_6  (
            .in0(N__35779),
            .in1(N__35683),
            .in2(N__34104),
            .in3(N__42007),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIALN65_1_LC_15_12_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIALN65_1_LC_15_12_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIALN65_1_LC_15_12_7 .LUT_INIT=16'b1000111110001111;
    LogicCell40 \ppm_encoder_1.throttle_RNIALN65_1_LC_15_12_7  (
            .in0(N__37553),
            .in1(N__34577),
            .in2(N__34092),
            .in3(N__37973),
            .lcout(\ppm_encoder_1.throttle_RNIALN65Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNI7RM01_LC_15_13_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNI7RM01_LC_15_13_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNI7RM01_LC_15_13_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNI7RM01_LC_15_13_0  (
            .in0(N__40472),
            .in1(N__40407),
            .in2(N__40378),
            .in3(N__41923),
            .lcout(\ppm_encoder_1.init_pulses_2_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_4_LC_15_13_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_4_LC_15_13_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_4_LC_15_13_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_4_LC_15_13_1  (
            .in0(N__34167),
            .in1(N__35378),
            .in2(_gnd_net_),
            .in3(N__40373),
            .lcout(),
            .ltout(\ppm_encoder_1.N_296_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_4_LC_15_13_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_4_LC_15_13_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_4_LC_15_13_2 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_4_LC_15_13_2  (
            .in0(_gnd_net_),
            .in1(N__38918),
            .in2(N__34146),
            .in3(N__34143),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNI7RM01_0_LC_15_13_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNI7RM01_0_LC_15_13_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNI7RM01_0_LC_15_13_4 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNI7RM01_0_LC_15_13_4  (
            .in0(N__40471),
            .in1(N__40406),
            .in2(N__40379),
            .in3(N__41924),
            .lcout(\ppm_encoder_1.init_pulses_0_sqmuxa_0 ),
            .ltout(\ppm_encoder_1.init_pulses_0_sqmuxa_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIO1KK2_6_LC_15_13_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIO1KK2_6_LC_15_13_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIO1KK2_6_LC_15_13_5 .LUT_INIT=16'b1000110010101111;
    LogicCell40 \ppm_encoder_1.throttle_RNIO1KK2_6_LC_15_13_5  (
            .in0(N__34276),
            .in1(N__36212),
            .in2(N__34125),
            .in3(N__35268),
            .lcout(\ppm_encoder_1.un2_throttle_iv_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_esr_RNI81QU2_14_LC_15_13_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_esr_RNI81QU2_14_LC_15_13_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_esr_RNI81QU2_14_LC_15_13_6 .LUT_INIT=16'b0000011101110111;
    LogicCell40 \ppm_encoder_1.throttle_esr_RNI81QU2_14_LC_15_13_6  (
            .in0(N__35269),
            .in1(N__41021),
            .in2(N__35649),
            .in3(N__37568),
            .lcout(\ppm_encoder_1.un2_throttle_iv_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNI8GVN2_6_LC_15_14_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNI8GVN2_6_LC_15_14_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNI8GVN2_6_LC_15_14_0 .LUT_INIT=16'b1010001011110011;
    LogicCell40 \ppm_encoder_1.elevator_RNI8GVN2_6_LC_15_14_0  (
            .in0(N__34366),
            .in1(N__35783),
            .in2(N__34335),
            .in3(N__35730),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_1_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIEDI96_6_LC_15_14_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIEDI96_6_LC_15_14_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIEDI96_6_LC_15_14_1 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ppm_encoder_1.throttle_RNIEDI96_6_LC_15_14_1  (
            .in0(N__37787),
            .in1(_gnd_net_),
            .in2(N__34122),
            .in3(N__34119),
            .lcout(\ppm_encoder_1.throttle_RNIEDI96Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_6_LC_15_14_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_6_LC_15_14_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_6_LC_15_14_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_6_LC_15_14_3  (
            .in0(N__40114),
            .in1(N__34277),
            .in2(_gnd_net_),
            .in3(N__34333),
            .lcout(),
            .ltout(\ppm_encoder_1.N_298_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_6_LC_15_14_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_6_LC_15_14_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_6_LC_15_14_4 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_6_LC_15_14_4  (
            .in0(N__34367),
            .in1(_gnd_net_),
            .in2(N__34371),
            .in3(N__38949),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_6_LC_15_14_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_6_LC_15_14_5 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.aileron_6_LC_15_14_5 .LUT_INIT=16'b0111011100100010;
    LogicCell40 \ppm_encoder_1.aileron_6_LC_15_14_5  (
            .in0(N__37250),
            .in1(N__35600),
            .in2(_gnd_net_),
            .in3(N__34368),
            .lcout(\ppm_encoder_1.aileronZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47350),
            .ce(),
            .sr(N__43870));
    defparam \ppm_encoder_1.elevator_6_LC_15_14_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_6_LC_15_14_6 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.elevator_6_LC_15_14_6 .LUT_INIT=16'b0011001110101010;
    LogicCell40 \ppm_encoder_1.elevator_6_LC_15_14_6  (
            .in0(N__34334),
            .in1(N__34355),
            .in2(_gnd_net_),
            .in3(N__37254),
            .lcout(\ppm_encoder_1.elevatorZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47350),
            .ce(),
            .sr(N__43870));
    defparam \ppm_encoder_1.throttle_6_LC_15_14_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_6_LC_15_14_7 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.throttle_6_LC_15_14_7 .LUT_INIT=16'b1001111110010000;
    LogicCell40 \ppm_encoder_1.throttle_6_LC_15_14_7  (
            .in0(N__34320),
            .in1(N__34308),
            .in2(N__37263),
            .in3(N__34278),
            .lcout(\ppm_encoder_1.throttleZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47350),
            .ce(),
            .sr(N__43870));
    defparam \ppm_encoder_1.elevator_RNICKVN2_8_LC_15_15_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNICKVN2_8_LC_15_15_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNICKVN2_8_LC_15_15_0 .LUT_INIT=16'b1010001011110011;
    LogicCell40 \ppm_encoder_1.elevator_RNICKVN2_8_LC_15_15_0  (
            .in0(N__38800),
            .in1(N__35800),
            .in2(N__34251),
            .in3(N__35734),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_1_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIONI96_8_LC_15_15_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIONI96_8_LC_15_15_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIONI96_8_LC_15_15_1 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ppm_encoder_1.throttle_RNIONI96_8_LC_15_15_1  (
            .in0(N__40623),
            .in1(_gnd_net_),
            .in2(N__34263),
            .in3(N__34260),
            .lcout(\ppm_encoder_1.throttle_RNIONI96Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_8_LC_15_15_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_8_LC_15_15_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_8_LC_15_15_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_8_LC_15_15_3  (
            .in0(N__40113),
            .in1(N__34183),
            .in2(_gnd_net_),
            .in3(N__34250),
            .lcout(\ppm_encoder_1.N_300 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_8_LC_15_15_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_8_LC_15_15_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_8_LC_15_15_5 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.throttle_8_LC_15_15_5  (
            .in0(N__34227),
            .in1(N__34200),
            .in2(N__37256),
            .in3(N__34184),
            .lcout(\ppm_encoder_1.throttleZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47333),
            .ce(),
            .sr(N__43877));
    defparam \ppm_encoder_1.aileron_8_LC_15_15_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_8_LC_15_15_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.aileron_8_LC_15_15_6 .LUT_INIT=16'b0010111011100010;
    LogicCell40 \ppm_encoder_1.aileron_8_LC_15_15_6  (
            .in0(N__38801),
            .in1(N__37214),
            .in2(N__36027),
            .in3(N__36047),
            .lcout(\ppm_encoder_1.aileronZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47333),
            .ce(),
            .sr(N__43877));
    defparam \ppm_encoder_1.rudder_8_LC_15_15_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_8_LC_15_15_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.rudder_8_LC_15_15_7 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.rudder_8_LC_15_15_7  (
            .in0(N__34542),
            .in1(N__34527),
            .in2(N__37255),
            .in3(N__38405),
            .lcout(\ppm_encoder_1.rudderZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47333),
            .ce(),
            .sr(N__43877));
    defparam \ppm_encoder_1.throttle_RNIK8JI2_13_LC_15_16_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIK8JI2_13_LC_15_16_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIK8JI2_13_LC_15_16_0 .LUT_INIT=16'b1011000010111011;
    LogicCell40 \ppm_encoder_1.throttle_RNIK8JI2_13_LC_15_16_0  (
            .in0(N__39001),
            .in1(N__35289),
            .in2(N__34425),
            .in3(N__37583),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNIKVRT5_13_LC_15_16_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNIKVRT5_13_LC_15_16_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNIKVRT5_13_LC_15_16_1 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ppm_encoder_1.elevator_RNIKVRT5_13_LC_15_16_1  (
            .in0(_gnd_net_),
            .in1(N__38045),
            .in2(N__34509),
            .in3(N__34506),
            .lcout(\ppm_encoder_1.elevator_RNIKVRT5Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNI47DH2_13_LC_15_16_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNI47DH2_13_LC_15_16_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNI47DH2_13_LC_15_16_2 .LUT_INIT=16'b1010001011110011;
    LogicCell40 \ppm_encoder_1.elevator_RNI47DH2_13_LC_15_16_2  (
            .in0(N__34384),
            .in1(N__35819),
            .in2(N__34407),
            .in3(N__35744),
            .lcout(\ppm_encoder_1.un2_throttle_iv_1_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_13_LC_15_16_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_13_LC_15_16_5 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.aileron_13_LC_15_16_5 .LUT_INIT=16'b1010010111001100;
    LogicCell40 \ppm_encoder_1.aileron_13_LC_15_16_5  (
            .in0(N__35883),
            .in1(N__34385),
            .in2(N__35907),
            .in3(N__37224),
            .lcout(\ppm_encoder_1.aileronZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47320),
            .ce(),
            .sr(N__43884));
    defparam \ppm_encoder_1.elevator_13_LC_15_16_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_13_LC_15_16_6 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.elevator_13_LC_15_16_6 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \ppm_encoder_1.elevator_13_LC_15_16_6  (
            .in0(N__34405),
            .in1(N__34500),
            .in2(N__37257),
            .in3(N__34476),
            .lcout(\ppm_encoder_1.elevatorZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47320),
            .ce(),
            .sr(N__43884));
    defparam \ppm_encoder_1.throttle_13_LC_15_16_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_13_LC_15_16_7 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.throttle_13_LC_15_16_7 .LUT_INIT=16'b1010010111001100;
    LogicCell40 \ppm_encoder_1.throttle_13_LC_15_16_7  (
            .in0(N__34464),
            .in1(N__34423),
            .in2(N__34440),
            .in3(N__37225),
            .lcout(\ppm_encoder_1.throttleZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47320),
            .ce(),
            .sr(N__43884));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_13_LC_15_17_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_13_LC_15_17_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_13_LC_15_17_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_13_LC_15_17_0  (
            .in0(N__40125),
            .in1(N__34424),
            .in2(_gnd_net_),
            .in3(N__34406),
            .lcout(),
            .ltout(\ppm_encoder_1.N_305_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_13_LC_15_17_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_13_LC_15_17_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_13_LC_15_17_1 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_13_LC_15_17_1  (
            .in0(_gnd_net_),
            .in1(N__38974),
            .in2(N__34389),
            .in3(N__34386),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_3_11_LC_15_17_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_3_11_LC_15_17_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_3_11_LC_15_17_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_3_11_LC_15_17_4  (
            .in0(N__40126),
            .in1(N__34631),
            .in2(_gnd_net_),
            .in3(N__34921),
            .lcout(),
            .ltout(\ppm_encoder_1.N_303_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_11_LC_15_17_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_11_LC_15_17_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_11_LC_15_17_5 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_11_LC_15_17_5  (
            .in0(_gnd_net_),
            .in1(N__38973),
            .in2(N__34614),
            .in3(N__36148),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNISFRP_13_LC_15_17_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNISFRP_13_LC_15_17_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNISFRP_13_LC_15_17_6 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNISFRP_13_LC_15_17_6  (
            .in0(N__41332),
            .in1(N__42233),
            .in2(_gnd_net_),
            .in3(N__41840),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNIALRT5_11_LC_15_17_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNIALRT5_11_LC_15_17_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNIALRT5_11_LC_15_17_7 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \ppm_encoder_1.elevator_RNIALRT5_11_LC_15_17_7  (
            .in0(N__38144),
            .in1(N__34611),
            .in2(_gnd_net_),
            .in3(N__34902),
            .lcout(\ppm_encoder_1.elevator_RNIALRT5Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_11_LC_15_18_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_11_LC_15_18_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_11_LC_15_18_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_11_LC_15_18_2  (
            .in0(N__34601),
            .in1(N__40927),
            .in2(_gnd_net_),
            .in3(N__37762),
            .lcout(),
            .ltout(\ppm_encoder_1.N_319_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_11_LC_15_18_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_11_LC_15_18_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_11_LC_15_18_3 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_11_LC_15_18_3  (
            .in0(_gnd_net_),
            .in1(N__41148),
            .in2(N__34584),
            .in3(N__35527),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_LC_15_18_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_LC_15_18_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_LC_15_18_4 .LUT_INIT=16'b1111000111111100;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_LC_15_18_4  (
            .in0(N__42234),
            .in1(N__40454),
            .in2(N__44137),
            .in3(N__41777),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47300),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_2_LC_15_18_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_2_LC_15_18_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_2_LC_15_18_5 .LUT_INIT=16'b0101000000000000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_2_LC_15_18_5  (
            .in0(N__40092),
            .in1(_gnd_net_),
            .in2(N__38984),
            .in3(N__37630),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_1_LC_15_18_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_1_LC_15_18_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_1_LC_15_18_6 .LUT_INIT=16'b1110111011111111;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_1_LC_15_18_6  (
            .in0(N__34581),
            .in1(N__40091),
            .in2(_gnd_net_),
            .in3(N__38976),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_10_LC_15_18_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_10_LC_15_18_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_10_LC_15_18_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_10_LC_15_18_7  (
            .in0(N__38975),
            .in1(N__34548),
            .in2(_gnd_net_),
            .in3(N__34737),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter_RNIAEV01_8_LC_15_19_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter_RNIAEV01_8_LC_15_19_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter_RNIAEV01_8_LC_15_19_0 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \ppm_encoder_1.counter_RNIAEV01_8_LC_15_19_0  (
            .in0(N__34638),
            .in1(N__42445),
            .in2(N__34647),
            .in3(N__39263),
            .lcout(\ppm_encoder_1.N_145_17 ),
            .ltout(\ppm_encoder_1.N_145_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.PPM_STATE_RNI09RH2_1_LC_15_19_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_RNI09RH2_1_LC_15_19_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.PPM_STATE_RNI09RH2_1_LC_15_19_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \ppm_encoder_1.PPM_STATE_RNI09RH2_1_LC_15_19_1  (
            .in0(N__34892),
            .in1(N__39641),
            .in2(N__34716),
            .in3(N__34653),
            .lcout(\ppm_encoder_1.N_238 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.ppm_output_reg_RNO_2_LC_15_19_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.ppm_output_reg_RNO_2_LC_15_19_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.ppm_output_reg_RNO_2_LC_15_19_2 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \ppm_encoder_1.ppm_output_reg_RNO_2_LC_15_19_2  (
            .in0(N__36371),
            .in1(N__39356),
            .in2(N__40321),
            .in3(N__39385),
            .lcout(\ppm_encoder_1.un1_PPM_STATE_1_sqmuxa_i_a3_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNI5GRT5_10_LC_15_19_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNI5GRT5_10_LC_15_19_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNI5GRT5_10_LC_15_19_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ppm_encoder_1.elevator_RNI5GRT5_10_LC_15_19_3  (
            .in0(N__39030),
            .in1(N__34692),
            .in2(_gnd_net_),
            .in3(N__34686),
            .lcout(\ppm_encoder_1.elevator_RNI5GRT5Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.PPM_STATE_RNISH5F_1_LC_15_19_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_RNISH5F_1_LC_15_19_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.PPM_STATE_RNISH5F_1_LC_15_19_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \ppm_encoder_1.PPM_STATE_RNISH5F_1_LC_15_19_4  (
            .in0(_gnd_net_),
            .in1(N__44084),
            .in2(_gnd_net_),
            .in3(N__41814),
            .lcout(\ppm_encoder_1.N_1330_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.PPM_STATE_RNISL0F_1_LC_15_19_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_RNISL0F_1_LC_15_19_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.PPM_STATE_RNISL0F_1_LC_15_19_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \ppm_encoder_1.PPM_STATE_RNISL0F_1_LC_15_19_5  (
            .in0(N__39355),
            .in1(N__36370),
            .in2(N__39387),
            .in3(N__34675),
            .lcout(\ppm_encoder_1.PPM_STATE_ns_0_a3_0_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter_RNIUS1G_4_LC_15_19_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter_RNIUS1G_4_LC_15_19_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter_RNIUS1G_4_LC_15_19_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \ppm_encoder_1.counter_RNIUS1G_4_LC_15_19_7  (
            .in0(N__42706),
            .in1(N__36320),
            .in2(N__42741),
            .in3(N__36341),
            .lcout(\ppm_encoder_1.PPM_STATE_ns_0_a3_0_17_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_1_c_RNO_LC_15_20_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_1_c_RNO_LC_15_20_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_1_c_RNO_LC_15_20_0 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_1_c_RNO_LC_15_20_0  (
            .in0(N__36081),
            .in1(N__36369),
            .in2(N__36393),
            .in3(N__36057),
            .lcout(\ppm_encoder_1.counter24_0_I_1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter_RNIDBJ8_13_LC_15_20_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter_RNIDBJ8_13_LC_15_20_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter_RNIDBJ8_13_LC_15_20_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \ppm_encoder_1.counter_RNIDBJ8_13_LC_15_20_2  (
            .in0(_gnd_net_),
            .in1(N__39245),
            .in2(_gnd_net_),
            .in3(N__42484),
            .lcout(\ppm_encoder_1.PPM_STATE_ns_0_a3_0_17_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_LC_15_20_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_LC_15_20_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_LC_15_20_3 .LUT_INIT=16'b0001001000100010;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_1_LC_15_20_3  (
            .in0(N__40055),
            .in1(N__44118),
            .in2(N__38985),
            .in3(N__41776),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47286),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNI03DH2_11_LC_15_20_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNI03DH2_11_LC_15_20_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNI03DH2_11_LC_15_20_4 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \ppm_encoder_1.elevator_RNI03DH2_11_LC_15_20_4  (
            .in0(N__36153),
            .in1(N__35820),
            .in2(N__34929),
            .in3(N__35745),
            .lcout(\ppm_encoder_1.un2_throttle_iv_1_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter_RNIK1KG_0_LC_15_20_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter_RNIK1KG_0_LC_15_20_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter_RNIK1KG_0_LC_15_20_5 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \ppm_encoder_1.counter_RNIK1KG_0_LC_15_20_5  (
            .in0(N__36391),
            .in1(N__44620),
            .in2(N__39294),
            .in3(N__44584),
            .lcout(\ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_reg_esr_1_LC_15_21_0 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_1_LC_15_21_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_1_LC_15_21_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_1_LC_15_21_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34881),
            .lcout(\pid_alt.error_i_regZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47277),
            .ce(N__46797),
            .sr(N__46593));
    defparam \reset_module_System.count_1_cry_1_c_LC_16_7_0 .C_ON=1'b1;
    defparam \reset_module_System.count_1_cry_1_c_LC_16_7_0 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_1_cry_1_c_LC_16_7_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \reset_module_System.count_1_cry_1_c_LC_16_7_0  (
            .in0(_gnd_net_),
            .in1(N__34854),
            .in2(N__34833),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_16_7_0_),
            .carryout(\reset_module_System.count_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNO_0_2_LC_16_7_1 .C_ON=1'b1;
    defparam \reset_module_System.count_RNO_0_2_LC_16_7_1 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNO_0_2_LC_16_7_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_RNO_0_2_LC_16_7_1  (
            .in0(_gnd_net_),
            .in1(N__34790),
            .in2(_gnd_net_),
            .in3(N__34773),
            .lcout(\reset_module_System.count_1_2 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_1 ),
            .carryout(\reset_module_System.count_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_3_LC_16_7_2 .C_ON=1'b1;
    defparam \reset_module_System.count_3_LC_16_7_2 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_3_LC_16_7_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_3_LC_16_7_2  (
            .in0(_gnd_net_),
            .in1(N__34769),
            .in2(_gnd_net_),
            .in3(N__34758),
            .lcout(\reset_module_System.countZ0Z_3 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_2 ),
            .carryout(\reset_module_System.count_1_cry_3 ),
            .clk(N__47443),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_4_LC_16_7_3 .C_ON=1'b1;
    defparam \reset_module_System.count_4_LC_16_7_3 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_4_LC_16_7_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_4_LC_16_7_3  (
            .in0(_gnd_net_),
            .in1(N__34754),
            .in2(_gnd_net_),
            .in3(N__34740),
            .lcout(\reset_module_System.countZ0Z_4 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_3 ),
            .carryout(\reset_module_System.count_1_cry_4 ),
            .clk(N__47443),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_5_LC_16_7_4 .C_ON=1'b1;
    defparam \reset_module_System.count_5_LC_16_7_4 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_5_LC_16_7_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_5_LC_16_7_4  (
            .in0(_gnd_net_),
            .in1(N__35034),
            .in2(_gnd_net_),
            .in3(N__35022),
            .lcout(\reset_module_System.countZ0Z_5 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_4 ),
            .carryout(\reset_module_System.count_1_cry_5 ),
            .clk(N__47443),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_6_LC_16_7_5 .C_ON=1'b1;
    defparam \reset_module_System.count_6_LC_16_7_5 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_6_LC_16_7_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_6_LC_16_7_5  (
            .in0(_gnd_net_),
            .in1(N__35018),
            .in2(_gnd_net_),
            .in3(N__35007),
            .lcout(\reset_module_System.countZ0Z_6 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_5 ),
            .carryout(\reset_module_System.count_1_cry_6 ),
            .clk(N__47443),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_7_LC_16_7_6 .C_ON=1'b1;
    defparam \reset_module_System.count_7_LC_16_7_6 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_7_LC_16_7_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_7_LC_16_7_6  (
            .in0(_gnd_net_),
            .in1(N__35004),
            .in2(_gnd_net_),
            .in3(N__34992),
            .lcout(\reset_module_System.countZ0Z_7 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_6 ),
            .carryout(\reset_module_System.count_1_cry_7 ),
            .clk(N__47443),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_8_LC_16_7_7 .C_ON=1'b1;
    defparam \reset_module_System.count_8_LC_16_7_7 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_8_LC_16_7_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_8_LC_16_7_7  (
            .in0(_gnd_net_),
            .in1(N__34989),
            .in2(_gnd_net_),
            .in3(N__34977),
            .lcout(\reset_module_System.countZ0Z_8 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_7 ),
            .carryout(\reset_module_System.count_1_cry_8 ),
            .clk(N__47443),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_9_LC_16_8_0 .C_ON=1'b1;
    defparam \reset_module_System.count_9_LC_16_8_0 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_9_LC_16_8_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_9_LC_16_8_0  (
            .in0(_gnd_net_),
            .in1(N__34970),
            .in2(_gnd_net_),
            .in3(N__34956),
            .lcout(\reset_module_System.countZ0Z_9 ),
            .ltout(),
            .carryin(bfn_16_8_0_),
            .carryout(\reset_module_System.count_1_cry_9 ),
            .clk(N__47437),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_10_LC_16_8_1 .C_ON=1'b1;
    defparam \reset_module_System.count_10_LC_16_8_1 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_10_LC_16_8_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_10_LC_16_8_1  (
            .in0(_gnd_net_),
            .in1(N__37331),
            .in2(_gnd_net_),
            .in3(N__34953),
            .lcout(\reset_module_System.countZ0Z_10 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_9 ),
            .carryout(\reset_module_System.count_1_cry_10 ),
            .clk(N__47437),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_11_LC_16_8_2 .C_ON=1'b1;
    defparam \reset_module_System.count_11_LC_16_8_2 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_11_LC_16_8_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_11_LC_16_8_2  (
            .in0(_gnd_net_),
            .in1(N__37370),
            .in2(_gnd_net_),
            .in3(N__34950),
            .lcout(\reset_module_System.countZ0Z_11 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_10 ),
            .carryout(\reset_module_System.count_1_cry_11 ),
            .clk(N__47437),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_12_LC_16_8_3 .C_ON=1'b1;
    defparam \reset_module_System.count_12_LC_16_8_3 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_12_LC_16_8_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_12_LC_16_8_3  (
            .in0(_gnd_net_),
            .in1(N__34946),
            .in2(_gnd_net_),
            .in3(N__34935),
            .lcout(\reset_module_System.countZ0Z_12 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_11 ),
            .carryout(\reset_module_System.count_1_cry_12 ),
            .clk(N__47437),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_13_LC_16_8_4 .C_ON=1'b1;
    defparam \reset_module_System.count_13_LC_16_8_4 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_13_LC_16_8_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_13_LC_16_8_4  (
            .in0(_gnd_net_),
            .in1(N__35157),
            .in2(_gnd_net_),
            .in3(N__34932),
            .lcout(\reset_module_System.countZ0Z_13 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_12 ),
            .carryout(\reset_module_System.count_1_cry_13 ),
            .clk(N__47437),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_14_LC_16_8_5 .C_ON=1'b1;
    defparam \reset_module_System.count_14_LC_16_8_5 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_14_LC_16_8_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_14_LC_16_8_5  (
            .in0(_gnd_net_),
            .in1(N__37358),
            .in2(_gnd_net_),
            .in3(N__35112),
            .lcout(\reset_module_System.countZ0Z_14 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_13 ),
            .carryout(\reset_module_System.count_1_cry_14 ),
            .clk(N__47437),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_15_LC_16_8_6 .C_ON=1'b1;
    defparam \reset_module_System.count_15_LC_16_8_6 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_15_LC_16_8_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_15_LC_16_8_6  (
            .in0(_gnd_net_),
            .in1(N__35181),
            .in2(_gnd_net_),
            .in3(N__35109),
            .lcout(\reset_module_System.countZ0Z_15 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_14 ),
            .carryout(\reset_module_System.count_1_cry_15 ),
            .clk(N__47437),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_16_LC_16_8_7 .C_ON=1'b1;
    defparam \reset_module_System.count_16_LC_16_8_7 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_16_LC_16_8_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_16_LC_16_8_7  (
            .in0(_gnd_net_),
            .in1(N__35106),
            .in2(_gnd_net_),
            .in3(N__35094),
            .lcout(\reset_module_System.countZ0Z_16 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_15 ),
            .carryout(\reset_module_System.count_1_cry_16 ),
            .clk(N__47437),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_17_LC_16_9_0 .C_ON=1'b1;
    defparam \reset_module_System.count_17_LC_16_9_0 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_17_LC_16_9_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_17_LC_16_9_0  (
            .in0(_gnd_net_),
            .in1(N__37343),
            .in2(_gnd_net_),
            .in3(N__35091),
            .lcout(\reset_module_System.countZ0Z_17 ),
            .ltout(),
            .carryin(bfn_16_9_0_),
            .carryout(\reset_module_System.count_1_cry_17 ),
            .clk(N__47427),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_18_LC_16_9_1 .C_ON=1'b1;
    defparam \reset_module_System.count_18_LC_16_9_1 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_18_LC_16_9_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_18_LC_16_9_1  (
            .in0(_gnd_net_),
            .in1(N__35087),
            .in2(_gnd_net_),
            .in3(N__35073),
            .lcout(\reset_module_System.countZ0Z_18 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_17 ),
            .carryout(\reset_module_System.count_1_cry_18 ),
            .clk(N__47427),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_19_LC_16_9_2 .C_ON=1'b1;
    defparam \reset_module_System.count_19_LC_16_9_2 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_19_LC_16_9_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \reset_module_System.count_19_LC_16_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__35046),
            .in3(N__35070),
            .lcout(\reset_module_System.countZ0Z_19 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_18 ),
            .carryout(\reset_module_System.count_1_cry_19 ),
            .clk(N__47427),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_20_LC_16_9_3 .C_ON=1'b1;
    defparam \reset_module_System.count_20_LC_16_9_3 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_20_LC_16_9_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_20_LC_16_9_3  (
            .in0(_gnd_net_),
            .in1(N__35066),
            .in2(_gnd_net_),
            .in3(N__35052),
            .lcout(\reset_module_System.countZ0Z_20 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_19 ),
            .carryout(\reset_module_System.count_1_cry_20 ),
            .clk(N__47427),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_21_LC_16_9_4 .C_ON=1'b0;
    defparam \reset_module_System.count_21_LC_16_9_4 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_21_LC_16_9_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \reset_module_System.count_21_LC_16_9_4  (
            .in0(N__35168),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35049),
            .lcout(\reset_module_System.countZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47427),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNI34OR1_21_LC_16_9_6 .C_ON=1'b0;
    defparam \reset_module_System.count_RNI34OR1_21_LC_16_9_6 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNI34OR1_21_LC_16_9_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \reset_module_System.count_RNI34OR1_21_LC_16_9_6  (
            .in0(N__35042),
            .in1(N__35180),
            .in2(N__35169),
            .in3(N__35156),
            .lcout(\reset_module_System.reset6_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_5_LC_16_10_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_5_LC_16_10_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_5_LC_16_10_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_5_LC_16_10_4  (
            .in0(N__35222),
            .in1(N__35408),
            .in2(_gnd_net_),
            .in3(N__40362),
            .lcout(),
            .ltout(\ppm_encoder_1.N_297_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_5_LC_16_10_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_5_LC_16_10_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_5_LC_16_10_5 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_5_LC_16_10_5  (
            .in0(_gnd_net_),
            .in1(N__38860),
            .in2(N__35136),
            .in3(N__35430),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNIE3D21_3_LC_16_10_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNIE3D21_3_LC_16_10_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNIE3D21_3_LC_16_10_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_RNIE3D21_3_LC_16_10_6  (
            .in0(N__40363),
            .in1(N__40490),
            .in2(N__40929),
            .in3(N__39993),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_159_d ),
            .ltout(\ppm_encoder_1.CHOOSE_CHANNEL_159_d_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNIGD613_3_LC_16_10_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNIGD613_3_LC_16_10_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNIGD613_3_LC_16_10_7 .LUT_INIT=16'b0000000000001010;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_RNIGD613_3_LC_16_10_7  (
            .in0(N__42038),
            .in1(_gnd_net_),
            .in2(N__35133),
            .in3(N__37704),
            .lcout(\ppm_encoder_1.un1_init_pulses_4_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIAVNR2_0_LC_16_11_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIAVNR2_0_LC_16_11_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIAVNR2_0_LC_16_11_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIAVNR2_0_LC_16_11_0  (
            .in0(N__41978),
            .in1(N__36941),
            .in2(N__37703),
            .in3(N__42337),
            .lcout(\ppm_encoder_1.init_pulses_RNIAVNR2Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_0_LC_16_11_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_0_LC_16_11_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_0_LC_16_11_2 .LUT_INIT=16'b1111111110111011;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_0_LC_16_11_2  (
            .in0(N__40132),
            .in1(N__38857),
            .in2(_gnd_net_),
            .in3(N__36965),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_3_LC_16_11_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_3_LC_16_11_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_3_LC_16_11_3 .LUT_INIT=16'b0101000001000100;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_3_LC_16_11_3  (
            .in0(N__44108),
            .in1(N__35130),
            .in2(N__35196),
            .in3(N__41977),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47406),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_3_LC_16_11_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_3_LC_16_11_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_3_LC_16_11_5 .LUT_INIT=16'b1111111111011101;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_3_LC_16_11_5  (
            .in0(N__38858),
            .in1(N__40133),
            .in2(_gnd_net_),
            .in3(N__35451),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_LC_16_11_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_LC_16_11_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_LC_16_11_6 .LUT_INIT=16'b1101110111001110;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_0_LC_16_11_6  (
            .in0(N__41976),
            .in1(N__44109),
            .in2(N__42231),
            .in3(N__38859),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47406),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.PPM_STATE_RNI2APU1_1_1_LC_16_11_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_RNI2APU1_1_1_LC_16_11_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.PPM_STATE_RNI2APU1_1_1_LC_16_11_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ppm_encoder_1.PPM_STATE_RNI2APU1_1_1_LC_16_11_7  (
            .in0(_gnd_net_),
            .in1(N__37687),
            .in2(_gnd_net_),
            .in3(N__41975),
            .lcout(\ppm_encoder_1.PPM_STATE_RNI2APU1_1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNI33GU_3_LC_16_12_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNI33GU_3_LC_16_12_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNI33GU_3_LC_16_12_0 .LUT_INIT=16'b0001000101010101;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_RNI33GU_3_LC_16_12_0  (
            .in0(N__39975),
            .in1(N__40130),
            .in2(_gnd_net_),
            .in3(N__40485),
            .lcout(\ppm_encoder_1.pulses2count_9_sn_N_10_mux ),
            .ltout(\ppm_encoder_1.pulses2count_9_sn_N_10_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_1_LC_16_12_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_1_LC_16_12_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_1_LC_16_12_1 .LUT_INIT=16'b1010111110001101;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_1_LC_16_12_1  (
            .in0(N__41122),
            .in1(N__40909),
            .in2(N__35385),
            .in3(N__37386),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.rudder_esr_RNITVNJ2_4_LC_16_12_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_esr_RNITVNJ2_4_LC_16_12_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.rudder_esr_RNITVNJ2_4_LC_16_12_2 .LUT_INIT=16'b1011000010111011;
    LogicCell40 \ppm_encoder_1.rudder_esr_RNITVNJ2_4_LC_16_12_2  (
            .in0(N__37454),
            .in1(N__35249),
            .in2(N__35382),
            .in3(N__37550),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_esr_RNIV9IN5_4_LC_16_12_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_esr_RNIV9IN5_4_LC_16_12_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.aileron_esr_RNIV9IN5_4_LC_16_12_3 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ppm_encoder_1.aileron_esr_RNIV9IN5_4_LC_16_12_3  (
            .in0(_gnd_net_),
            .in1(N__37865),
            .in2(N__35349),
            .in3(N__35346),
            .lcout(\ppm_encoder_1.aileron_esr_RNIV9IN5Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIQ3KK2_7_LC_16_12_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIQ3KK2_7_LC_16_12_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIQ3KK2_7_LC_16_12_4 .LUT_INIT=16'b0000011101110111;
    LogicCell40 \ppm_encoder_1.throttle_RNIQ3KK2_7_LC_16_12_4  (
            .in0(N__40691),
            .in1(N__35250),
            .in2(N__35340),
            .in3(N__37551),
            .lcout(\ppm_encoder_1.un2_throttle_iv_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI8J2H_2_LC_16_12_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI8J2H_2_LC_16_12_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI8J2H_2_LC_16_12_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI8J2H_2_LC_16_12_5  (
            .in0(_gnd_net_),
            .in1(N__35307),
            .in2(_gnd_net_),
            .in3(N__39974),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_d_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.rudder_esr_RNIV1OJ2_5_LC_16_12_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_esr_RNIV1OJ2_5_LC_16_12_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.rudder_esr_RNIV1OJ2_5_LC_16_12_6 .LUT_INIT=16'b0000011101110111;
    LogicCell40 \ppm_encoder_1.rudder_esr_RNIV1OJ2_5_LC_16_12_6  (
            .in0(N__37412),
            .in1(N__35248),
            .in2(N__35226),
            .in3(N__37549),
            .lcout(\ppm_encoder_1.un2_throttle_iv_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_3_LC_16_12_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_3_LC_16_12_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_3_LC_16_12_7 .LUT_INIT=16'b0011001000010000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_3_LC_16_12_7  (
            .in0(N__42002),
            .in1(N__44117),
            .in2(N__39991),
            .in3(N__35192),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47390),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_3_LC_16_13_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_3_LC_16_13_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.init_pulses_3_LC_16_13_0 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_3_LC_16_13_0  (
            .in0(N__41611),
            .in1(N__39867),
            .in2(N__41444),
            .in3(N__37887),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47376),
            .ce(),
            .sr(N__43871));
    defparam \ppm_encoder_1.throttle_RNIT9352_3_LC_16_13_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIT9352_3_LC_16_13_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIT9352_3_LC_16_13_1 .LUT_INIT=16'b1001011010011001;
    LogicCell40 \ppm_encoder_1.throttle_RNIT9352_3_LC_16_13_1  (
            .in0(N__35549),
            .in1(N__42327),
            .in2(N__35450),
            .in3(N__37548),
            .lcout(),
            .ltout(\ppm_encoder_1.un1_init_pulses_0_axb_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNI82223_3_LC_16_13_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNI82223_3_LC_16_13_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNI82223_3_LC_16_13_2 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \ppm_encoder_1.throttle_RNI82223_3_LC_16_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__35553),
            .in3(N__37898),
            .lcout(\ppm_encoder_1.throttle_RNI82223Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIBOUS_3_LC_16_13_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIBOUS_3_LC_16_13_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIBOUS_3_LC_16_13_3 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIBOUS_3_LC_16_13_3  (
            .in0(N__35547),
            .in1(N__42151),
            .in2(_gnd_net_),
            .in3(N__41995),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIBOUS_0_3_LC_16_13_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIBOUS_0_3_LC_16_13_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIBOUS_0_3_LC_16_13_4 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIBOUS_0_3_LC_16_13_4  (
            .in0(N__41996),
            .in1(_gnd_net_),
            .in2(N__42228),
            .in3(N__35548),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_3_LC_16_13_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_3_LC_16_13_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_3_LC_16_13_5 .LUT_INIT=16'b1010111110001101;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_3_LC_16_13_5  (
            .in0(N__41124),
            .in1(N__35550),
            .in2(N__35531),
            .in3(N__40948),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_2_LC_16_13_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_2_LC_16_13_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_2_LC_16_13_6 .LUT_INIT=16'b0011101100001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_2_LC_16_13_6  (
            .in0(N__37653),
            .in1(N__41123),
            .in2(N__40977),
            .in3(N__35523),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_3_LC_16_13_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_3_LC_16_13_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_3_LC_16_13_7 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \ppm_encoder_1.throttle_3_LC_16_13_7  (
            .in0(N__35446),
            .in1(N__35490),
            .in2(N__37262),
            .in3(N__35478),
            .lcout(\ppm_encoder_1.throttleZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47376),
            .ce(),
            .sr(N__43871));
    defparam \ppm_encoder_1.aileron_esr_RNIOIR62_5_LC_16_14_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_esr_RNIOIR62_5_LC_16_14_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.aileron_esr_RNIOIR62_5_LC_16_14_0 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \ppm_encoder_1.aileron_esr_RNIOIR62_5_LC_16_14_0  (
            .in0(N__35429),
            .in1(N__35781),
            .in2(N__35409),
            .in3(N__35728),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_1_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_esr_RNI4FIN5_5_LC_16_14_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_esr_RNI4FIN5_5_LC_16_14_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.aileron_esr_RNI4FIN5_5_LC_16_14_1 .LUT_INIT=16'b0000111111111111;
    LogicCell40 \ppm_encoder_1.aileron_esr_RNI4FIN5_5_LC_16_14_1  (
            .in0(N__37833),
            .in1(_gnd_net_),
            .in2(N__35832),
            .in3(N__35829),
            .lcout(\ppm_encoder_1.aileron_esr_RNI4FIN5Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_esr_RNIOVDS2_14_LC_16_14_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_esr_RNIOVDS2_14_LC_16_14_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.aileron_esr_RNIOVDS2_14_LC_16_14_2 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \ppm_encoder_1.aileron_esr_RNIOVDS2_14_LC_16_14_2  (
            .in0(N__38373),
            .in1(N__35782),
            .in2(N__35625),
            .in3(N__35729),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_1_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_esr_RNITH3L6_14_LC_16_14_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_esr_RNITH3L6_14_LC_16_14_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.aileron_esr_RNITH3L6_14_LC_16_14_3 .LUT_INIT=16'b0000111111111111;
    LogicCell40 \ppm_encoder_1.aileron_esr_RNITH3L6_14_LC_16_14_3  (
            .in0(N__41190),
            .in1(_gnd_net_),
            .in2(N__35658),
            .in3(N__35655),
            .lcout(\ppm_encoder_1.aileron_esr_RNITH3L6Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIANUS_2_LC_16_14_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIANUS_2_LC_16_14_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIANUS_2_LC_16_14_4 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIANUS_2_LC_16_14_4  (
            .in0(N__37650),
            .in1(N__42172),
            .in2(_gnd_net_),
            .in3(N__41993),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_14_LC_16_14_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_14_LC_16_14_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_14_LC_16_14_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_14_LC_16_14_5  (
            .in0(N__35645),
            .in1(N__40121),
            .in2(_gnd_net_),
            .in3(N__35624),
            .lcout(\ppm_encoder_1.N_306 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI7O1N_0_2_LC_16_14_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI7O1N_0_2_LC_16_14_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI7O1N_0_2_LC_16_14_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI7O1N_0_2_LC_16_14_6  (
            .in0(_gnd_net_),
            .in1(N__42171),
            .in2(_gnd_net_),
            .in3(N__41992),
            .lcout(\ppm_encoder_1.un1_init_pulses_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIERUS_6_LC_16_14_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIERUS_6_LC_16_14_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIERUS_6_LC_16_14_7 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIERUS_6_LC_16_14_7  (
            .in0(N__41994),
            .in1(_gnd_net_),
            .in2(N__42232),
            .in3(N__37486),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_6_c_LC_16_15_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_6_c_LC_16_15_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_6_c_LC_16_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_6_c_LC_16_15_0  (
            .in0(_gnd_net_),
            .in1(N__35604),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_16_15_0_),
            .carryout(\ppm_encoder_1.un1_aileron_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_6_THRU_LUT4_0_LC_16_15_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_6_THRU_LUT4_0_LC_16_15_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_6_THRU_LUT4_0_LC_16_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_6_THRU_LUT4_0_LC_16_15_1  (
            .in0(_gnd_net_),
            .in1(N__35586),
            .in2(_gnd_net_),
            .in3(N__35556),
            .lcout(\ppm_encoder_1.un1_aileron_cry_6_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_6 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_7_THRU_LUT4_0_LC_16_15_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_7_THRU_LUT4_0_LC_16_15_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_7_THRU_LUT4_0_LC_16_15_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_7_THRU_LUT4_0_LC_16_15_2  (
            .in0(_gnd_net_),
            .in1(N__36048),
            .in2(_gnd_net_),
            .in3(N__36018),
            .lcout(\ppm_encoder_1.un1_aileron_cry_7_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_7 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_8_THRU_LUT4_0_LC_16_15_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_8_THRU_LUT4_0_LC_16_15_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_8_THRU_LUT4_0_LC_16_15_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_8_THRU_LUT4_0_LC_16_15_3  (
            .in0(_gnd_net_),
            .in1(N__36015),
            .in2(_gnd_net_),
            .in3(N__35988),
            .lcout(\ppm_encoder_1.un1_aileron_cry_8_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_8 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_9_THRU_LUT4_0_LC_16_15_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_9_THRU_LUT4_0_LC_16_15_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_9_THRU_LUT4_0_LC_16_15_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_9_THRU_LUT4_0_LC_16_15_4  (
            .in0(_gnd_net_),
            .in1(N__35984),
            .in2(_gnd_net_),
            .in3(N__35952),
            .lcout(\ppm_encoder_1.un1_aileron_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_9 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_10_THRU_LUT4_0_LC_16_15_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_10_THRU_LUT4_0_LC_16_15_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_10_THRU_LUT4_0_LC_16_15_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_10_THRU_LUT4_0_LC_16_15_5  (
            .in0(_gnd_net_),
            .in1(N__36185),
            .in2(_gnd_net_),
            .in3(N__35949),
            .lcout(\ppm_encoder_1.un1_aileron_cry_10_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_10 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_11_THRU_LUT4_0_LC_16_15_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_11_THRU_LUT4_0_LC_16_15_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_11_THRU_LUT4_0_LC_16_15_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_11_THRU_LUT4_0_LC_16_15_6  (
            .in0(_gnd_net_),
            .in1(N__35945),
            .in2(_gnd_net_),
            .in3(N__35910),
            .lcout(\ppm_encoder_1.un1_aileron_cry_11_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_11 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_12_THRU_LUT4_0_LC_16_15_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_12_THRU_LUT4_0_LC_16_15_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_12_THRU_LUT4_0_LC_16_15_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_12_THRU_LUT4_0_LC_16_15_7  (
            .in0(_gnd_net_),
            .in1(N__35906),
            .in2(N__43050),
            .in3(N__35877),
            .lcout(\ppm_encoder_1.un1_aileron_cry_12_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_12 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_esr_14_LC_16_16_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_esr_14_LC_16_16_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.aileron_esr_14_LC_16_16_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ppm_encoder_1.aileron_esr_14_LC_16_16_0  (
            .in0(_gnd_net_),
            .in1(N__35874),
            .in2(_gnd_net_),
            .in3(N__35862),
            .lcout(\ppm_encoder_1.aileronZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47334),
            .ce(N__36227),
            .sr(N__43887));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_10_LC_16_17_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_10_LC_16_17_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_10_LC_16_17_0 .LUT_INIT=16'b1010100000001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_10_LC_16_17_0  (
            .in0(N__41145),
            .in1(N__41247),
            .in2(N__40991),
            .in3(N__35859),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.rudder_13_LC_16_17_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_13_LC_16_17_2 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.rudder_13_LC_16_17_2 .LUT_INIT=16'b1001111110010000;
    LogicCell40 \ppm_encoder_1.rudder_13_LC_16_17_2  (
            .in0(N__36294),
            .in1(N__36279),
            .in2(N__37227),
            .in3(N__39005),
            .lcout(\ppm_encoder_1.rudderZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47321),
            .ce(),
            .sr(N__43892));
    defparam \ppm_encoder_1.rudder_esr_ctle_14_LC_16_17_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_esr_ctle_14_LC_16_17_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.rudder_esr_ctle_14_LC_16_17_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \ppm_encoder_1.rudder_esr_ctle_14_LC_16_17_3  (
            .in0(_gnd_net_),
            .in1(N__37165),
            .in2(_gnd_net_),
            .in3(N__44074),
            .lcout(\ppm_encoder_1.pid_altitude_dv_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_6_LC_16_17_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_6_LC_16_17_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_6_LC_16_17_5 .LUT_INIT=16'b1110010011111111;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_6_LC_16_17_5  (
            .in0(N__40982),
            .in1(N__37494),
            .in2(N__36216),
            .in3(N__41146),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_11_LC_16_17_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_11_LC_16_17_6 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.aileron_11_LC_16_17_6 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.aileron_11_LC_16_17_6  (
            .in0(N__36186),
            .in1(N__36162),
            .in2(N__37226),
            .in3(N__36149),
            .lcout(\ppm_encoder_1.aileronZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47321),
            .ce(),
            .sr(N__43892));
    defparam \ppm_encoder_1.counter24_0_I_15_c_RNO_LC_16_18_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_15_c_RNO_LC_16_18_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_15_c_RNO_LC_16_18_0 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_15_c_RNO_LC_16_18_0  (
            .in0(N__36117),
            .in1(N__36319),
            .in2(N__36099),
            .in3(N__36340),
            .lcout(\ppm_encoder_1.counter24_0_I_15_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_4_LC_16_18_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_4_LC_16_18_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_4_LC_16_18_1 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_4_LC_16_18_1  (
            .in0(N__37440),
            .in1(_gnd_net_),
            .in2(N__42617),
            .in3(N__36129),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47310),
            .ce(N__42540),
            .sr(N__43894));
    defparam \ppm_encoder_1.pulses2count_esr_5_LC_16_18_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_5_LC_16_18_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_5_LC_16_18_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_5_LC_16_18_2  (
            .in0(N__36111),
            .in1(N__42603),
            .in2(_gnd_net_),
            .in3(N__37398),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47310),
            .ce(N__42540),
            .sr(N__43894));
    defparam \ppm_encoder_1.pulses2count_esr_0_LC_16_18_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_0_LC_16_18_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_0_LC_16_18_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_0_LC_16_18_3  (
            .in0(N__42598),
            .in1(N__36090),
            .in2(_gnd_net_),
            .in3(N__36921),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47310),
            .ce(N__42540),
            .sr(N__43894));
    defparam \ppm_encoder_1.pulses2count_esr_1_LC_16_18_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_1_LC_16_18_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_1_LC_16_18_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_1_LC_16_18_5  (
            .in0(N__42599),
            .in1(N__36072),
            .in2(_gnd_net_),
            .in3(N__36066),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47310),
            .ce(N__42540),
            .sr(N__43894));
    defparam \ppm_encoder_1.counter_0_LC_16_19_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_0_LC_16_19_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_0_LC_16_19_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_0_LC_16_19_0  (
            .in0(_gnd_net_),
            .in1(N__36392),
            .in2(N__36417),
            .in3(N__36416),
            .lcout(\ppm_encoder_1.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_16_19_0_),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_0 ),
            .clk(N__47301),
            .ce(),
            .sr(N__36903));
    defparam \ppm_encoder_1.counter_1_LC_16_19_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_1_LC_16_19_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_1_LC_16_19_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_1_LC_16_19_1  (
            .in0(_gnd_net_),
            .in1(N__36372),
            .in2(_gnd_net_),
            .in3(N__36351),
            .lcout(\ppm_encoder_1.counterZ0Z_1 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_0 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_1 ),
            .clk(N__47301),
            .ce(),
            .sr(N__36903));
    defparam \ppm_encoder_1.counter_2_LC_16_19_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_2_LC_16_19_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_2_LC_16_19_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_2_LC_16_19_2  (
            .in0(_gnd_net_),
            .in1(N__39357),
            .in2(_gnd_net_),
            .in3(N__36348),
            .lcout(\ppm_encoder_1.counterZ0Z_2 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_1 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_2 ),
            .clk(N__47301),
            .ce(),
            .sr(N__36903));
    defparam \ppm_encoder_1.counter_3_LC_16_19_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_3_LC_16_19_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_3_LC_16_19_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_3_LC_16_19_3  (
            .in0(_gnd_net_),
            .in1(N__39386),
            .in2(_gnd_net_),
            .in3(N__36345),
            .lcout(\ppm_encoder_1.counterZ0Z_3 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_2 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_3 ),
            .clk(N__47301),
            .ce(),
            .sr(N__36903));
    defparam \ppm_encoder_1.counter_4_LC_16_19_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_4_LC_16_19_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_4_LC_16_19_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_4_LC_16_19_4  (
            .in0(_gnd_net_),
            .in1(N__36342),
            .in2(_gnd_net_),
            .in3(N__36324),
            .lcout(\ppm_encoder_1.counterZ0Z_4 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_3 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_4 ),
            .clk(N__47301),
            .ce(),
            .sr(N__36903));
    defparam \ppm_encoder_1.counter_5_LC_16_19_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_5_LC_16_19_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_5_LC_16_19_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_5_LC_16_19_5  (
            .in0(_gnd_net_),
            .in1(N__36321),
            .in2(_gnd_net_),
            .in3(N__36303),
            .lcout(\ppm_encoder_1.counterZ0Z_5 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_4 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_5 ),
            .clk(N__47301),
            .ce(),
            .sr(N__36903));
    defparam \ppm_encoder_1.counter_6_LC_16_19_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_6_LC_16_19_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_6_LC_16_19_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_6_LC_16_19_6  (
            .in0(_gnd_net_),
            .in1(N__42708),
            .in2(_gnd_net_),
            .in3(N__36300),
            .lcout(\ppm_encoder_1.counterZ0Z_6 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_5 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_6 ),
            .clk(N__47301),
            .ce(),
            .sr(N__36903));
    defparam \ppm_encoder_1.counter_7_LC_16_19_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_7_LC_16_19_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_7_LC_16_19_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_7_LC_16_19_7  (
            .in0(_gnd_net_),
            .in1(N__42740),
            .in2(_gnd_net_),
            .in3(N__36297),
            .lcout(\ppm_encoder_1.counterZ0Z_7 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_6 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_7 ),
            .clk(N__47301),
            .ce(),
            .sr(N__36903));
    defparam \ppm_encoder_1.counter_8_LC_16_20_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_8_LC_16_20_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_8_LC_16_20_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_8_LC_16_20_0  (
            .in0(_gnd_net_),
            .in1(N__39264),
            .in2(_gnd_net_),
            .in3(N__36447),
            .lcout(\ppm_encoder_1.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_16_20_0_),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_8 ),
            .clk(N__47292),
            .ce(),
            .sr(N__36902));
    defparam \ppm_encoder_1.counter_9_LC_16_20_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_9_LC_16_20_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_9_LC_16_20_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_9_LC_16_20_1  (
            .in0(_gnd_net_),
            .in1(N__39293),
            .in2(_gnd_net_),
            .in3(N__36444),
            .lcout(\ppm_encoder_1.counterZ0Z_9 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_8 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_9 ),
            .clk(N__47292),
            .ce(),
            .sr(N__36902));
    defparam \ppm_encoder_1.counter_10_LC_16_20_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_10_LC_16_20_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_10_LC_16_20_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_10_LC_16_20_2  (
            .in0(_gnd_net_),
            .in1(N__44585),
            .in2(_gnd_net_),
            .in3(N__36441),
            .lcout(\ppm_encoder_1.counterZ0Z_10 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_9 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_10 ),
            .clk(N__47292),
            .ce(),
            .sr(N__36902));
    defparam \ppm_encoder_1.counter_11_LC_16_20_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_11_LC_16_20_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_11_LC_16_20_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_11_LC_16_20_3  (
            .in0(_gnd_net_),
            .in1(N__44621),
            .in2(_gnd_net_),
            .in3(N__36438),
            .lcout(\ppm_encoder_1.counterZ0Z_11 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_10 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_11 ),
            .clk(N__47292),
            .ce(),
            .sr(N__36902));
    defparam \ppm_encoder_1.counter_12_LC_16_20_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_12_LC_16_20_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_12_LC_16_20_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_12_LC_16_20_4  (
            .in0(_gnd_net_),
            .in1(N__42446),
            .in2(_gnd_net_),
            .in3(N__36435),
            .lcout(\ppm_encoder_1.counterZ0Z_12 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_11 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_12 ),
            .clk(N__47292),
            .ce(),
            .sr(N__36902));
    defparam \ppm_encoder_1.counter_13_LC_16_20_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_13_LC_16_20_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_13_LC_16_20_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_13_LC_16_20_5  (
            .in0(_gnd_net_),
            .in1(N__42485),
            .in2(_gnd_net_),
            .in3(N__36432),
            .lcout(\ppm_encoder_1.counterZ0Z_13 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_12 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_13 ),
            .clk(N__47292),
            .ce(),
            .sr(N__36902));
    defparam \ppm_encoder_1.counter_14_LC_16_20_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_14_LC_16_20_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_14_LC_16_20_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_14_LC_16_20_6  (
            .in0(_gnd_net_),
            .in1(N__39246),
            .in2(_gnd_net_),
            .in3(N__36429),
            .lcout(\ppm_encoder_1.counterZ0Z_14 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_13 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_14 ),
            .clk(N__47292),
            .ce(),
            .sr(N__36902));
    defparam \ppm_encoder_1.counter_15_LC_16_20_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_15_LC_16_20_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_15_LC_16_20_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_15_LC_16_20_7  (
            .in0(_gnd_net_),
            .in1(N__39699),
            .in2(_gnd_net_),
            .in3(N__36426),
            .lcout(\ppm_encoder_1.counterZ0Z_15 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_14 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_15 ),
            .clk(N__47292),
            .ce(),
            .sr(N__36902));
    defparam \ppm_encoder_1.counter_16_LC_16_21_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_16_LC_16_21_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_16_LC_16_21_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_16_LC_16_21_0  (
            .in0(_gnd_net_),
            .in1(N__39659),
            .in2(_gnd_net_),
            .in3(N__36423),
            .lcout(\ppm_encoder_1.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_16_21_0_),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_16 ),
            .clk(N__47287),
            .ce(),
            .sr(N__36901));
    defparam \ppm_encoder_1.counter_17_LC_16_21_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_17_LC_16_21_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_17_LC_16_21_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_17_LC_16_21_1  (
            .in0(_gnd_net_),
            .in1(N__39682),
            .in2(_gnd_net_),
            .in3(N__36420),
            .lcout(\ppm_encoder_1.counterZ0Z_17 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_16 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_17 ),
            .clk(N__47287),
            .ce(),
            .sr(N__36901));
    defparam \ppm_encoder_1.counter_18_LC_16_21_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter_18_LC_16_21_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_18_LC_16_21_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ppm_encoder_1.counter_18_LC_16_21_2  (
            .in0(_gnd_net_),
            .in1(N__39612),
            .in2(_gnd_net_),
            .in3(N__36906),
            .lcout(\ppm_encoder_1.counterZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47287),
            .ce(),
            .sr(N__36901));
    defparam \Commands_frame_decoder.source_alt_ki_2_LC_16_22_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_ki_2_LC_16_22_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_ki_2_LC_16_22_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_ki_2_LC_16_22_2  (
            .in0(_gnd_net_),
            .in1(N__36887),
            .in2(_gnd_net_),
            .in3(N__46678),
            .lcout(alt_ki_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47278),
            .ce(N__44849),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_reg_esr_2_LC_16_23_6 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_2_LC_16_23_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_2_LC_16_23_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_2_LC_16_23_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36738),
            .lcout(\pid_alt.error_i_regZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47274),
            .ce(N__46795),
            .sr(N__46586));
    defparam \uart_drone.timer_Count_RNIU8TV1_3_LC_17_7_3 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_RNIU8TV1_3_LC_17_7_3 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNIU8TV1_3_LC_17_7_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uart_drone.timer_Count_RNIU8TV1_3_LC_17_7_3  (
            .in0(N__44461),
            .in1(N__36618),
            .in2(_gnd_net_),
            .in3(N__36549),
            .lcout(\uart_drone.N_144_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.bit_Count_2_LC_17_8_2 .C_ON=1'b0;
    defparam \uart_drone.bit_Count_2_LC_17_8_2 .SEQ_MODE=4'b1000;
    defparam \uart_drone.bit_Count_2_LC_17_8_2 .LUT_INIT=16'b0000000001111000;
    LogicCell40 \uart_drone.bit_Count_2_LC_17_8_2  (
            .in0(N__39537),
            .in1(N__39495),
            .in2(N__36686),
            .in3(N__39531),
            .lcout(\uart_drone.bit_CountZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47444),
            .ce(),
            .sr(N__43839));
    defparam \uart_drone.state_RNI62411_4_LC_17_9_2 .C_ON=1'b0;
    defparam \uart_drone.state_RNI62411_4_LC_17_9_2 .SEQ_MODE=4'b0000;
    defparam \uart_drone.state_RNI62411_4_LC_17_9_2 .LUT_INIT=16'b0000000010001111;
    LogicCell40 \uart_drone.state_RNI62411_4_LC_17_9_2  (
            .in0(N__36617),
            .in1(N__36545),
            .in2(N__44552),
            .in3(N__36489),
            .lcout(\uart_drone.un1_state_4_0 ),
            .ltout(\uart_drone.un1_state_4_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_RNI63LK2_3_LC_17_9_3 .C_ON=1'b0;
    defparam \uart_drone.state_RNI63LK2_3_LC_17_9_3 .SEQ_MODE=4'b0000;
    defparam \uart_drone.state_RNI63LK2_3_LC_17_9_3 .LUT_INIT=16'b1111000000110000;
    LogicCell40 \uart_drone.state_RNI63LK2_3_LC_17_9_3  (
            .in0(_gnd_net_),
            .in1(N__44548),
            .in2(N__36450),
            .in3(N__44451),
            .lcout(\uart_drone.un1_state_7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_0_LC_17_9_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNO_0_0_LC_17_9_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_0_LC_17_9_4 .LUT_INIT=16'b0110011000110011;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_0_LC_17_9_4  (
            .in0(N__36966),
            .in1(N__38000),
            .in2(_gnd_net_),
            .in3(N__37596),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNISRMR1_10_LC_17_9_5 .C_ON=1'b0;
    defparam \reset_module_System.count_RNISRMR1_10_LC_17_9_5 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNISRMR1_10_LC_17_9_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \reset_module_System.count_RNISRMR1_10_LC_17_9_5  (
            .in0(N__37371),
            .in1(N__37359),
            .in2(N__37347),
            .in3(N__37332),
            .lcout(\reset_module_System.reset6_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_0_LC_17_10_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNO_1_0_LC_17_10_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_0_LC_17_10_1 .LUT_INIT=16'b1000011101111000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_0_LC_17_10_1  (
            .in0(N__42035),
            .in1(N__37713),
            .in2(N__36945),
            .in3(N__42348),
            .lcout(),
            .ltout(\ppm_encoder_1.un1_init_pulses_11_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_0_LC_17_10_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_0_LC_17_10_2 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_0_LC_17_10_2 .LUT_INIT=16'b0100010001010000;
    LogicCell40 \ppm_encoder_1.init_pulses_0_LC_17_10_2  (
            .in0(N__41615),
            .in1(N__37275),
            .in2(N__37269),
            .in3(N__41380),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47428),
            .ce(),
            .sr(N__43855));
    defparam \ppm_encoder_1.init_pulses_RNI8LUS_0_LC_17_10_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI8LUS_0_LC_17_10_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI8LUS_0_LC_17_10_4 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI8LUS_0_LC_17_10_4  (
            .in0(N__36939),
            .in1(N__42229),
            .in2(_gnd_net_),
            .in3(N__42034),
            .lcout(\ppm_encoder_1.un1_init_pulses_0 ),
            .ltout(\ppm_encoder_1.un1_init_pulses_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIN3352_0_LC_17_10_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIN3352_0_LC_17_10_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIN3352_0_LC_17_10_5 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \ppm_encoder_1.throttle_RNIN3352_0_LC_17_10_5  (
            .in0(_gnd_net_),
            .in1(N__36963),
            .in2(N__37266),
            .in3(N__37592),
            .lcout(\ppm_encoder_1.throttle_RNIN3352Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_0_LC_17_10_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_0_LC_17_10_6 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.throttle_0_LC_17_10_6 .LUT_INIT=16'b0010001011101110;
    LogicCell40 \ppm_encoder_1.throttle_0_LC_17_10_6  (
            .in0(N__36964),
            .in1(N__37203),
            .in2(_gnd_net_),
            .in3(N__36996),
            .lcout(\ppm_encoder_1.throttleZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47428),
            .ce(),
            .sr(N__43855));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_0_LC_17_10_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_0_LC_17_10_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_0_LC_17_10_7 .LUT_INIT=16'b1111111111110101;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_0_LC_17_10_7  (
            .in0(N__41062),
            .in1(_gnd_net_),
            .in2(N__40930),
            .in3(N__36940),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_4_LC_17_11_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_4_LC_17_11_0 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_4_LC_17_11_0 .LUT_INIT=16'b0011001000000010;
    LogicCell40 \ppm_encoder_1.init_pulses_4_LC_17_11_0  (
            .in0(N__39846),
            .in1(N__41616),
            .in2(N__41411),
            .in3(N__37851),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47417),
            .ce(),
            .sr(N__43861));
    defparam \ppm_encoder_1.init_pulses_RNICPUS_0_4_LC_17_11_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNICPUS_0_4_LC_17_11_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNICPUS_0_4_LC_17_11_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNICPUS_0_4_LC_17_11_1  (
            .in0(N__42162),
            .in1(N__37469),
            .in2(_gnd_net_),
            .in3(N__41984),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNICPUS_4_LC_17_11_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNICPUS_4_LC_17_11_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNICPUS_4_LC_17_11_2 .LUT_INIT=16'b0101101010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNICPUS_4_LC_17_11_2  (
            .in0(N__37468),
            .in1(_gnd_net_),
            .in2(N__42037),
            .in3(N__42164),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_4_LC_17_11_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_4_LC_17_11_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_4_LC_17_11_3 .LUT_INIT=16'b1010100000001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_4_LC_17_11_3  (
            .in0(N__41063),
            .in1(N__37470),
            .in2(N__40983),
            .in3(N__37458),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_5_LC_17_11_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_5_LC_17_11_4 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_5_LC_17_11_4 .LUT_INIT=16'b0011001000000010;
    LogicCell40 \ppm_encoder_1.init_pulses_5_LC_17_11_4  (
            .in0(N__39831),
            .in1(N__41617),
            .in2(N__41412),
            .in3(N__37809),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47417),
            .ce(),
            .sr(N__43861));
    defparam \ppm_encoder_1.init_pulses_RNIDQUS_5_LC_17_11_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIDQUS_5_LC_17_11_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIDQUS_5_LC_17_11_5 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIDQUS_5_LC_17_11_5  (
            .in0(N__42165),
            .in1(N__41991),
            .in2(_gnd_net_),
            .in3(N__37426),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIDQUS_0_5_LC_17_11_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIDQUS_0_5_LC_17_11_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIDQUS_0_5_LC_17_11_6 .LUT_INIT=16'b0101101010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIDQUS_0_5_LC_17_11_6  (
            .in0(N__37427),
            .in1(_gnd_net_),
            .in2(N__42036),
            .in3(N__42163),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_5_LC_17_11_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_5_LC_17_11_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_5_LC_17_11_7 .LUT_INIT=16'b1010100000001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_5_LC_17_11_7  (
            .in0(N__41064),
            .in1(N__37428),
            .in2(N__40984),
            .in3(N__37416),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_1_LC_17_12_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_1_LC_17_12_2 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_1_LC_17_12_2 .LUT_INIT=16'b0000000011100100;
    LogicCell40 \ppm_encoder_1.init_pulses_1_LC_17_12_2  (
            .in0(N__41423),
            .in1(N__39924),
            .in2(N__37953),
            .in3(N__41606),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47407),
            .ce(),
            .sr(N__43872));
    defparam \ppm_encoder_1.init_pulses_RNI9MUS_1_LC_17_12_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI9MUS_1_LC_17_12_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI9MUS_1_LC_17_12_3 .LUT_INIT=16'b0101101010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI9MUS_1_LC_17_12_3  (
            .in0(N__37384),
            .in1(_gnd_net_),
            .in2(N__42230),
            .in3(N__41998),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNI9MUS_0_1_LC_17_12_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI9MUS_0_1_LC_17_12_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI9MUS_0_1_LC_17_12_4 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI9MUS_0_1_LC_17_12_4  (
            .in0(N__41997),
            .in1(N__42158),
            .in2(_gnd_net_),
            .in3(N__37385),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_10_LC_17_12_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_10_LC_17_12_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.init_pulses_10_LC_17_12_5 .LUT_INIT=16'b0000111000000010;
    LogicCell40 \ppm_encoder_1.init_pulses_10_LC_17_12_5  (
            .in0(N__40221),
            .in1(N__41419),
            .in2(N__41619),
            .in3(N__38175),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47407),
            .ce(),
            .sr(N__43872));
    defparam \ppm_encoder_1.init_pulses_11_LC_17_12_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_11_LC_17_12_6 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_11_LC_17_12_6 .LUT_INIT=16'b0011001000000010;
    LogicCell40 \ppm_encoder_1.init_pulses_11_LC_17_12_6  (
            .in0(N__40194),
            .in1(N__41602),
            .in2(N__41446),
            .in3(N__38124),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47407),
            .ce(),
            .sr(N__43872));
    defparam \ppm_encoder_1.init_pulses_12_LC_17_12_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_12_LC_17_12_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.init_pulses_12_LC_17_12_7 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_12_LC_17_12_7  (
            .in0(N__41601),
            .in1(N__40173),
            .in2(N__41447),
            .in3(N__38076),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47407),
            .ce(),
            .sr(N__43872));
    defparam \ppm_encoder_1.init_pulses_RNIC1OR2_2_LC_17_13_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIC1OR2_2_LC_17_13_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIC1OR2_2_LC_17_13_0 .LUT_INIT=16'b0110011001100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIC1OR2_2_LC_17_13_0  (
            .in0(N__37652),
            .in1(N__42324),
            .in2(N__37719),
            .in3(N__42003),
            .lcout(\ppm_encoder_1.init_pulses_RNIC1OR2Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIG5OR2_6_LC_17_13_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIG5OR2_6_LC_17_13_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIG5OR2_6_LC_17_13_1 .LUT_INIT=16'b0110011001100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIG5OR2_6_LC_17_13_1  (
            .in0(N__42325),
            .in1(N__37487),
            .in2(N__42039),
            .in3(N__37717),
            .lcout(\ppm_encoder_1.init_pulses_RNIG5OR2Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIUPKO2_13_LC_17_13_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIUPKO2_13_LC_17_13_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIUPKO2_13_LC_17_13_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIUPKO2_13_LC_17_13_2  (
            .in0(N__37718),
            .in1(N__42326),
            .in2(N__42047),
            .in3(N__41337),
            .lcout(\ppm_encoder_1.init_pulses_RNIUPKO2Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_2_LC_17_13_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_2_LC_17_13_3 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_2_LC_17_13_3 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_2_LC_17_13_3  (
            .in0(N__41595),
            .in1(N__39894),
            .in2(N__41448),
            .in3(N__37917),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47391),
            .ce(),
            .sr(N__43878));
    defparam \ppm_encoder_1.throttle_RNIR7352_2_LC_17_13_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIR7352_2_LC_17_13_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIR7352_2_LC_17_13_4 .LUT_INIT=16'b1001011001100110;
    LogicCell40 \ppm_encoder_1.throttle_RNIR7352_2_LC_17_13_4  (
            .in0(N__37651),
            .in1(N__42323),
            .in2(N__37632),
            .in3(N__37574),
            .lcout(),
            .ltout(\ppm_encoder_1.un1_init_pulses_0_axb_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNI5V123_2_LC_17_13_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNI5V123_2_LC_17_13_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNI5V123_2_LC_17_13_5 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \ppm_encoder_1.throttle_RNI5V123_2_LC_17_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__37497),
            .in3(N__37928),
            .lcout(\ppm_encoder_1.throttle_RNI5V123Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_6_LC_17_13_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_6_LC_17_13_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.init_pulses_6_LC_17_13_7 .LUT_INIT=16'b0000111000000010;
    LogicCell40 \ppm_encoder_1.init_pulses_6_LC_17_13_7  (
            .in0(N__39792),
            .in1(N__41445),
            .in2(N__41618),
            .in3(N__37773),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47391),
            .ce(),
            .sr(N__43878));
    defparam \ppm_encoder_1.throttle_RNIVO123_0_LC_17_14_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.throttle_RNIVO123_0_LC_17_14_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIVO123_0_LC_17_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.throttle_RNIVO123_0_LC_17_14_0  (
            .in0(_gnd_net_),
            .in1(N__38016),
            .in2(N__38004),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_17_14_0_),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_1_LC_17_14_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_1_LC_17_14_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_1_LC_17_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_1_LC_17_14_1  (
            .in0(_gnd_net_),
            .in1(N__37986),
            .in2(N__37974),
            .in3(N__37941),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_1 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_0 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_2_LC_17_14_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_2_LC_17_14_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_2_LC_17_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_2_LC_17_14_2  (
            .in0(_gnd_net_),
            .in1(N__37938),
            .in2(N__37932),
            .in3(N__37911),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_2 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_1 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_3_LC_17_14_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_3_LC_17_14_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_3_LC_17_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_3_LC_17_14_3  (
            .in0(_gnd_net_),
            .in1(N__37908),
            .in2(N__37902),
            .in3(N__37881),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_3 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_2 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_4_LC_17_14_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_4_LC_17_14_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_4_LC_17_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_4_LC_17_14_4  (
            .in0(_gnd_net_),
            .in1(N__37878),
            .in2(N__37869),
            .in3(N__37842),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_4 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_3 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_5_LC_17_14_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_5_LC_17_14_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_5_LC_17_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_5_LC_17_14_5  (
            .in0(_gnd_net_),
            .in1(N__37839),
            .in2(N__37832),
            .in3(N__37800),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_5 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_4 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_6_LC_17_14_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_6_LC_17_14_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_6_LC_17_14_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_6_LC_17_14_6  (
            .in0(_gnd_net_),
            .in1(N__37797),
            .in2(N__37788),
            .in3(N__37767),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_6 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_5 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_7_LC_17_14_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_7_LC_17_14_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_7_LC_17_14_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_7_LC_17_14_7  (
            .in0(_gnd_net_),
            .in1(N__38226),
            .in2(N__40247),
            .in3(N__38214),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_7 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_6 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_8_LC_17_15_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_8_LC_17_15_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_8_LC_17_15_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_8_LC_17_15_0  (
            .in0(_gnd_net_),
            .in1(N__38211),
            .in2(N__40622),
            .in3(N__38202),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_8 ),
            .ltout(),
            .carryin(bfn_17_15_0_),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_9_LC_17_15_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_9_LC_17_15_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_9_LC_17_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_9_LC_17_15_1  (
            .in0(_gnd_net_),
            .in1(N__38199),
            .in2(N__40575),
            .in3(N__38190),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_9 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_8 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_10_LC_17_15_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_10_LC_17_15_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_10_LC_17_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_10_LC_17_15_2  (
            .in0(_gnd_net_),
            .in1(N__38187),
            .in2(N__39029),
            .in3(N__38166),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_10 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_9 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_11_LC_17_15_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_11_LC_17_15_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_11_LC_17_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_11_LC_17_15_3  (
            .in0(_gnd_net_),
            .in1(N__38163),
            .in2(N__38151),
            .in3(N__38115),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_11 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_10 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_12_LC_17_15_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_12_LC_17_15_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_12_LC_17_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_12_LC_17_15_4  (
            .in0(_gnd_net_),
            .in1(N__38112),
            .in2(N__38100),
            .in3(N__38067),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_12 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_11 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_13_LC_17_15_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_13_LC_17_15_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_13_LC_17_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_13_LC_17_15_5  (
            .in0(_gnd_net_),
            .in1(N__38064),
            .in2(N__38052),
            .in3(N__38031),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_13 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_12 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_14_LC_17_15_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_14_LC_17_15_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_14_LC_17_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_14_LC_17_15_6  (
            .in0(_gnd_net_),
            .in1(N__41183),
            .in2(N__38028),
            .in3(N__38019),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_14 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_13 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_15_LC_17_15_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_15_LC_17_15_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_15_LC_17_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_15_LC_17_15_7  (
            .in0(_gnd_net_),
            .in1(N__42405),
            .in2(N__38451),
            .in3(N__38433),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_15 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_14 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_16_LC_17_16_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_16_LC_17_16_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_16_LC_17_16_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_16_LC_17_16_0  (
            .in0(_gnd_net_),
            .in1(N__38379),
            .in2(_gnd_net_),
            .in3(N__38430),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_16 ),
            .ltout(),
            .carryin(bfn_17_16_0_),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_17_LC_17_16_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_17_LC_17_16_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_17_LC_17_16_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_17_LC_17_16_1  (
            .in0(_gnd_net_),
            .in1(N__38427),
            .in2(_gnd_net_),
            .in3(N__38412),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_17 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_16 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_18_LC_17_16_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNO_0_18_LC_17_16_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_18_LC_17_16_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_18_LC_17_16_2  (
            .in0(N__41673),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38409),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_8_LC_17_16_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_8_LC_17_16_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_8_LC_17_16_3 .LUT_INIT=16'b1100100000001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_8_LC_17_16_3  (
            .in0(N__40644),
            .in1(N__41132),
            .in2(N__40992),
            .in3(N__38406),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIVIRP_0_16_LC_17_16_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIVIRP_0_16_LC_17_16_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIVIRP_0_16_LC_17_16_4 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIVIRP_0_16_LC_17_16_4  (
            .in0(N__40798),
            .in1(N__42273),
            .in2(_gnd_net_),
            .in3(N__41939),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_14_LC_17_16_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_14_LC_17_16_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_14_LC_17_16_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_14_LC_17_16_7  (
            .in0(N__38972),
            .in1(N__38372),
            .in2(_gnd_net_),
            .in3(N__38358),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un9_error_filt_add_1_axb_0_LC_17_17_0 .C_ON=1'b1;
    defparam \pid_alt.un9_error_filt_add_1_axb_0_LC_17_17_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un9_error_filt_add_1_axb_0_LC_17_17_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \pid_alt.un9_error_filt_add_1_axb_0_LC_17_17_0  (
            .in0(_gnd_net_),
            .in1(N__38349),
            .in2(N__38334),
            .in3(_gnd_net_),
            .lcout(\pid_alt.un9_error_filt_add_1_axbZ0Z_0 ),
            .ltout(),
            .carryin(bfn_17_17_0_),
            .carryout(\pid_alt.un9_error_filt_add_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un9_error_filt_add_1_cry_1_s_LC_17_17_1 .C_ON=1'b1;
    defparam \pid_alt.un9_error_filt_add_1_cry_1_s_LC_17_17_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un9_error_filt_add_1_cry_1_s_LC_17_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.un9_error_filt_add_1_cry_1_s_LC_17_17_1  (
            .in0(_gnd_net_),
            .in1(N__38289),
            .in2(N__38274),
            .in3(N__38229),
            .lcout(\pid_alt.un9_error_filt_add_1_cry_1_sZ0 ),
            .ltout(),
            .carryin(\pid_alt.un9_error_filt_add_1_cry_0 ),
            .carryout(\pid_alt.un9_error_filt_add_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un9_error_filt_add_1_cry_2_s_LC_17_17_2 .C_ON=1'b1;
    defparam \pid_alt.un9_error_filt_add_1_cry_2_s_LC_17_17_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un9_error_filt_add_1_cry_2_s_LC_17_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.un9_error_filt_add_1_cry_2_s_LC_17_17_2  (
            .in0(_gnd_net_),
            .in1(N__38775),
            .in2(N__38760),
            .in3(N__38718),
            .lcout(\pid_alt.un9_error_filt_add_1_cry_2_sZ0 ),
            .ltout(),
            .carryin(\pid_alt.un9_error_filt_add_1_cry_1 ),
            .carryout(\pid_alt.un9_error_filt_add_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un9_error_filt_add_1_cry_3_s_LC_17_17_3 .C_ON=1'b1;
    defparam \pid_alt.un9_error_filt_add_1_cry_3_s_LC_17_17_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un9_error_filt_add_1_cry_3_s_LC_17_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.un9_error_filt_add_1_cry_3_s_LC_17_17_3  (
            .in0(_gnd_net_),
            .in1(N__38715),
            .in2(N__38700),
            .in3(N__38658),
            .lcout(\pid_alt.un9_error_filt_add_1_cry_3_sZ0 ),
            .ltout(),
            .carryin(\pid_alt.un9_error_filt_add_1_cry_2 ),
            .carryout(\pid_alt.un9_error_filt_add_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un9_error_filt_add_1_cry_4_s_LC_17_17_4 .C_ON=1'b1;
    defparam \pid_alt.un9_error_filt_add_1_cry_4_s_LC_17_17_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un9_error_filt_add_1_cry_4_s_LC_17_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.un9_error_filt_add_1_cry_4_s_LC_17_17_4  (
            .in0(_gnd_net_),
            .in1(N__39107),
            .in2(N__38655),
            .in3(N__38625),
            .lcout(\pid_alt.un9_error_filt_add_1_cry_4_sZ0 ),
            .ltout(),
            .carryin(\pid_alt.un9_error_filt_add_1_cry_3 ),
            .carryout(\pid_alt.un9_error_filt_add_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un9_error_filt_add_1_cry_5_s_LC_17_17_5 .C_ON=1'b1;
    defparam \pid_alt.un9_error_filt_add_1_cry_5_s_LC_17_17_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un9_error_filt_add_1_cry_5_s_LC_17_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.un9_error_filt_add_1_cry_5_s_LC_17_17_5  (
            .in0(_gnd_net_),
            .in1(N__38622),
            .in2(N__39124),
            .in3(N__38592),
            .lcout(\pid_alt.un9_error_filt_add_1_cry_5_sZ0 ),
            .ltout(),
            .carryin(\pid_alt.un9_error_filt_add_1_cry_4 ),
            .carryout(\pid_alt.un9_error_filt_add_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un9_error_filt_add_1_cry_6_s_LC_17_17_6 .C_ON=1'b1;
    defparam \pid_alt.un9_error_filt_add_1_cry_6_s_LC_17_17_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un9_error_filt_add_1_cry_6_s_LC_17_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.un9_error_filt_add_1_cry_6_s_LC_17_17_6  (
            .in0(_gnd_net_),
            .in1(N__39111),
            .in2(N__38589),
            .in3(N__38547),
            .lcout(\pid_alt.un9_error_filt_add_1_cry_6_sZ0 ),
            .ltout(),
            .carryin(\pid_alt.un9_error_filt_add_1_cry_5 ),
            .carryout(\pid_alt.un9_error_filt_add_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un9_error_filt_add_1_cry_7_s_LC_17_17_7 .C_ON=1'b1;
    defparam \pid_alt.un9_error_filt_add_1_cry_7_s_LC_17_17_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un9_error_filt_add_1_cry_7_s_LC_17_17_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.un9_error_filt_add_1_cry_7_s_LC_17_17_7  (
            .in0(_gnd_net_),
            .in1(N__38544),
            .in2(N__39125),
            .in3(N__38502),
            .lcout(\pid_alt.un9_error_filt_add_1_cry_7_sZ0 ),
            .ltout(),
            .carryin(\pid_alt.un9_error_filt_add_1_cry_6 ),
            .carryout(\pid_alt.un9_error_filt_add_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un9_error_filt_add_1_cry_8_s_LC_17_18_0 .C_ON=1'b1;
    defparam \pid_alt.un9_error_filt_add_1_cry_8_s_LC_17_18_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un9_error_filt_add_1_cry_8_s_LC_17_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.un9_error_filt_add_1_cry_8_s_LC_17_18_0  (
            .in0(_gnd_net_),
            .in1(N__39126),
            .in2(N__38499),
            .in3(N__38454),
            .lcout(\pid_alt.un9_error_filt_add_1_cry_8_sZ0 ),
            .ltout(),
            .carryin(bfn_17_18_0_),
            .carryout(\pid_alt.un9_error_filt_add_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un9_error_filt_add_1_cry_9_s_LC_17_18_1 .C_ON=1'b1;
    defparam \pid_alt.un9_error_filt_add_1_cry_9_s_LC_17_18_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un9_error_filt_add_1_cry_9_s_LC_17_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.un9_error_filt_add_1_cry_9_s_LC_17_18_1  (
            .in0(_gnd_net_),
            .in1(N__39216),
            .in2(N__39132),
            .in3(N__39180),
            .lcout(\pid_alt.un9_error_filt_add_1_cry_9_sZ0 ),
            .ltout(),
            .carryin(\pid_alt.un9_error_filt_add_1_cry_8 ),
            .carryout(\pid_alt.un9_error_filt_add_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un9_error_filt_add_1_cry_10_s_LC_17_18_2 .C_ON=1'b1;
    defparam \pid_alt.un9_error_filt_add_1_cry_10_s_LC_17_18_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un9_error_filt_add_1_cry_10_s_LC_17_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.un9_error_filt_add_1_cry_10_s_LC_17_18_2  (
            .in0(_gnd_net_),
            .in1(N__39130),
            .in2(N__39177),
            .in3(N__39135),
            .lcout(\pid_alt.un9_error_filt_add_1_cry_10_sZ0 ),
            .ltout(),
            .carryin(\pid_alt.un9_error_filt_add_1_cry_9 ),
            .carryout(\pid_alt.un9_error_filt_add_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un9_error_filt_add_1_s_11_LC_17_18_3 .C_ON=1'b0;
    defparam \pid_alt.un9_error_filt_add_1_s_11_LC_17_18_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un9_error_filt_add_1_s_11_LC_17_18_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.un9_error_filt_add_1_s_11_LC_17_18_3  (
            .in0(N__39131),
            .in1(N__39081),
            .in2(_gnd_net_),
            .in3(N__39063),
            .lcout(\pid_alt.un9_error_filt_add_1_sZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.ppm_output_reg_RNO_0_LC_17_18_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.ppm_output_reg_RNO_0_LC_17_18_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.ppm_output_reg_RNO_0_LC_17_18_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ppm_encoder_1.ppm_output_reg_RNO_0_LC_17_18_4  (
            .in0(N__44661),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40325),
            .lcout(\ppm_encoder_1.N_140_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIPCRP_10_LC_17_18_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIPCRP_10_LC_17_18_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIPCRP_10_LC_17_18_5 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIPCRP_10_LC_17_18_5  (
            .in0(N__41246),
            .in1(N__42289),
            .in2(_gnd_net_),
            .in3(N__41921),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNIC2521_1_LC_17_18_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNIC2521_1_LC_17_18_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNIC2521_1_LC_17_18_6 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_RNIC2521_1_LC_17_18_6  (
            .in0(N__38947),
            .in1(N__40129),
            .in2(_gnd_net_),
            .in3(N__40425),
            .lcout(\ppm_encoder_1.pulses2count_9_sn_N_11_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_13_LC_17_18_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_13_LC_17_18_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_13_LC_17_18_7 .LUT_INIT=16'b1011100011111111;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_13_LC_17_18_7  (
            .in0(N__39006),
            .in1(N__40990),
            .in2(N__41336),
            .in3(N__41147),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_8_LC_17_19_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_8_LC_17_19_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_8_LC_17_19_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_8_LC_17_19_0  (
            .in0(N__38948),
            .in1(N__38823),
            .in2(_gnd_net_),
            .in3(N__38808),
            .lcout(),
            .ltout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_8_LC_17_19_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_8_LC_17_19_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_8_LC_17_19_1 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_8_LC_17_19_1  (
            .in0(_gnd_net_),
            .in1(N__42610),
            .in2(N__38787),
            .in3(N__38784),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47311),
            .ce(N__42531),
            .sr(N__43897));
    defparam \ppm_encoder_1.pulses2count_esr_9_LC_17_19_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_9_LC_17_19_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_9_LC_17_19_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_9_LC_17_19_2  (
            .in0(N__42611),
            .in1(N__39447),
            .in2(_gnd_net_),
            .in3(N__40515),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47311),
            .ce(N__42531),
            .sr(N__43897));
    defparam \ppm_encoder_1.pulses2count_esr_13_LC_17_19_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_13_LC_17_19_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_13_LC_17_19_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_13_LC_17_19_3  (
            .in0(N__39432),
            .in1(N__42607),
            .in2(_gnd_net_),
            .in3(N__39417),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47311),
            .ce(N__42531),
            .sr(N__43897));
    defparam \ppm_encoder_1.pulses2count_esr_2_LC_17_19_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_2_LC_17_19_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_2_LC_17_19_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_2_LC_17_19_4  (
            .in0(N__42608),
            .in1(N__39411),
            .in2(_gnd_net_),
            .in3(N__39399),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47311),
            .ce(N__42531),
            .sr(N__43897));
    defparam \ppm_encoder_1.counter24_0_I_9_c_RNO_LC_17_19_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_9_c_RNO_LC_17_19_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_9_c_RNO_LC_17_19_5 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_9_c_RNO_LC_17_19_5  (
            .in0(N__39381),
            .in1(N__39363),
            .in2(N__39309),
            .in3(N__39354),
            .lcout(\ppm_encoder_1.counter24_0_I_9_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_3_LC_17_19_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_3_LC_17_19_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_3_LC_17_19_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_3_LC_17_19_6  (
            .in0(N__42609),
            .in1(N__39336),
            .in2(_gnd_net_),
            .in3(N__39321),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47311),
            .ce(N__42531),
            .sr(N__43897));
    defparam \ppm_encoder_1.counter24_0_I_27_c_RNO_LC_17_19_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_27_c_RNO_LC_17_19_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_27_c_RNO_LC_17_19_7 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_27_c_RNO_LC_17_19_7  (
            .in0(N__39300),
            .in1(N__39289),
            .in2(N__39273),
            .in3(N__39262),
            .lcout(\ppm_encoder_1.counter24_0_I_27_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_45_c_RNO_LC_17_20_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_45_c_RNO_LC_17_20_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_45_c_RNO_LC_17_20_0 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_45_c_RNO_LC_17_20_0  (
            .in0(N__41289),
            .in1(N__39697),
            .in2(N__39228),
            .in3(N__39244),
            .lcout(\ppm_encoder_1.counter24_0_I_45_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_15_LC_17_20_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_15_LC_17_20_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_15_LC_17_20_1 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \ppm_encoder_1.pulses2count_15_LC_17_20_1  (
            .in0(N__42369),
            .in1(N__39227),
            .in2(N__39746),
            .in3(N__41941),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47302),
            .ce(),
            .sr(N__43900));
    defparam \ppm_encoder_1.counter24_0_I_51_c_RNO_LC_17_20_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_51_c_RNO_LC_17_20_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_51_c_RNO_LC_17_20_3 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_51_c_RNO_LC_17_20_3  (
            .in0(N__39655),
            .in1(N__39755),
            .in2(N__39683),
            .in3(N__39780),
            .lcout(\ppm_encoder_1.counter24_0_I_51_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_17_LC_17_20_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_17_LC_17_20_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_17_LC_17_20_4 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \ppm_encoder_1.pulses2count_17_LC_17_20_4  (
            .in0(N__41940),
            .in1(N__39742),
            .in2(N__39759),
            .in3(N__40754),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47302),
            .ce(),
            .sr(N__43900));
    defparam \ppm_encoder_1.pulses2count_18_LC_17_20_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_18_LC_17_20_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_18_LC_17_20_5 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \ppm_encoder_1.pulses2count_18_LC_17_20_5  (
            .in0(N__41651),
            .in1(N__39624),
            .in2(N__39747),
            .in3(N__41942),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47302),
            .ce(),
            .sr(N__43900));
    defparam \ppm_encoder_1.counter_RNI637H_18_LC_17_20_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter_RNI637H_18_LC_17_20_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter_RNI637H_18_LC_17_20_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \ppm_encoder_1.counter_RNI637H_18_LC_17_20_7  (
            .in0(N__39698),
            .in1(N__39684),
            .in2(N__39660),
            .in3(N__39611),
            .lcout(\ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNO_LC_17_21_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNO_LC_17_21_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNO_LC_17_21_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ppm_encoder_1.counter24_0_I_57_c_RNO_LC_17_21_2  (
            .in0(_gnd_net_),
            .in1(N__39623),
            .in2(_gnd_net_),
            .in3(N__39610),
            .lcout(\ppm_encoder_1.counter24_0_I_57_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_reg_esr_0_LC_17_23_5 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_0_LC_17_23_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_0_LC_17_23_5 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \pid_alt.error_i_reg_esr_0_LC_17_23_5  (
            .in0(_gnd_net_),
            .in1(N__39594),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_i_regZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47279),
            .ce(N__46798),
            .sr(N__46585));
    defparam \pid_alt.error_i_reg_esr_3_LC_17_23_6 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_3_LC_17_23_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_3_LC_17_23_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_3_LC_17_23_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39561),
            .lcout(\pid_alt.error_i_regZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47279),
            .ce(N__46798),
            .sr(N__46585));
    defparam \uart_drone.bit_Count_RNO_0_2_LC_18_8_0 .C_ON=1'b0;
    defparam \uart_drone.bit_Count_RNO_0_2_LC_18_8_0 .SEQ_MODE=4'b0000;
    defparam \uart_drone.bit_Count_RNO_0_2_LC_18_8_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uart_drone.bit_Count_RNO_0_2_LC_18_8_0  (
            .in0(_gnd_net_),
            .in1(N__44485),
            .in2(_gnd_net_),
            .in3(N__44382),
            .lcout(\uart_drone.CO0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.bit_Count_1_LC_18_9_3 .C_ON=1'b0;
    defparam \uart_drone.bit_Count_1_LC_18_9_3 .SEQ_MODE=4'b1000;
    defparam \uart_drone.bit_Count_1_LC_18_9_3 .LUT_INIT=16'b0001001000100010;
    LogicCell40 \uart_drone.bit_Count_1_LC_18_9_3  (
            .in0(N__39494),
            .in1(N__39530),
            .in2(N__44495),
            .in3(N__44392),
            .lcout(\uart_drone.bit_CountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47445),
            .ce(),
            .sr(N__43856));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNI33GU_0_3_LC_18_10_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNI33GU_0_3_LC_18_10_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNI33GU_0_3_LC_18_10_5 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_RNI33GU_0_3_LC_18_10_5  (
            .in0(N__40140),
            .in1(N__40491),
            .in2(_gnd_net_),
            .in3(N__39992),
            .lcout(\ppm_encoder_1.pulses2count_9_sn_N_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIC9HQ4_0_LC_18_11_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNIC9HQ4_0_LC_18_11_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIC9HQ4_0_LC_18_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIC9HQ4_0_LC_18_11_0  (
            .in0(_gnd_net_),
            .in1(N__39951),
            .in2(N__39942),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_18_11_0_),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_1_LC_18_11_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_1_LC_18_11_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_1_LC_18_11_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_1_LC_18_11_1  (
            .in0(_gnd_net_),
            .in1(N__39930),
            .in2(_gnd_net_),
            .in3(N__39918),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_1 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_0 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_2_LC_18_11_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_2_LC_18_11_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_2_LC_18_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_2_LC_18_11_2  (
            .in0(_gnd_net_),
            .in1(N__39915),
            .in2(N__39906),
            .in3(N__39882),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_2 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_1 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_3_LC_18_11_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_3_LC_18_11_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_3_LC_18_11_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_3_LC_18_11_3  (
            .in0(_gnd_net_),
            .in1(N__39879),
            .in2(_gnd_net_),
            .in3(N__39855),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_3 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_2 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_4_LC_18_11_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_4_LC_18_11_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_4_LC_18_11_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_4_LC_18_11_4  (
            .in0(_gnd_net_),
            .in1(N__39852),
            .in2(_gnd_net_),
            .in3(N__39840),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_4 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_3 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_5_LC_18_11_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_5_LC_18_11_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_5_LC_18_11_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_5_LC_18_11_5  (
            .in0(_gnd_net_),
            .in1(N__39837),
            .in2(_gnd_net_),
            .in3(N__39825),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_5 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_4 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_6_LC_18_11_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_6_LC_18_11_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_6_LC_18_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_6_LC_18_11_6  (
            .in0(_gnd_net_),
            .in1(N__39822),
            .in2(N__39804),
            .in3(N__39783),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_6 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_5 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_7_LC_18_11_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_7_LC_18_11_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_7_LC_18_11_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_7_LC_18_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__40722),
            .in3(N__40230),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_7 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_6 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_8_LC_18_12_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_8_LC_18_12_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_8_LC_18_12_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_8_LC_18_12_0  (
            .in0(_gnd_net_),
            .in1(N__40272),
            .in2(_gnd_net_),
            .in3(N__40227),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_8 ),
            .ltout(),
            .carryin(bfn_18_12_0_),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_9_LC_18_12_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_9_LC_18_12_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_9_LC_18_12_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_9_LC_18_12_1  (
            .in0(_gnd_net_),
            .in1(N__40584),
            .in2(_gnd_net_),
            .in3(N__40224),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_9 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_8 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_10_LC_18_12_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_10_LC_18_12_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_10_LC_18_12_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_10_LC_18_12_2  (
            .in0(_gnd_net_),
            .in1(N__41217),
            .in2(_gnd_net_),
            .in3(N__40215),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_10 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_9 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_11_LC_18_12_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_11_LC_18_12_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_11_LC_18_12_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_11_LC_18_12_3  (
            .in0(_gnd_net_),
            .in1(N__40212),
            .in2(_gnd_net_),
            .in3(N__40188),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_11 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_10 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_12_LC_18_12_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_12_LC_18_12_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_12_LC_18_12_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_12_LC_18_12_4  (
            .in0(_gnd_net_),
            .in1(N__40185),
            .in2(_gnd_net_),
            .in3(N__40167),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_12 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_11 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_13_LC_18_12_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_13_LC_18_12_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_13_LC_18_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_13_LC_18_12_5  (
            .in0(_gnd_net_),
            .in1(N__40164),
            .in2(N__40158),
            .in3(N__40146),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_13 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_12 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_14_LC_18_12_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_14_LC_18_12_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_14_LC_18_12_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_14_LC_18_12_6  (
            .in0(_gnd_net_),
            .in1(N__41172),
            .in2(_gnd_net_),
            .in3(N__40143),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_14 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_13 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_15_LC_18_12_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_15_LC_18_12_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_15_LC_18_12_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_15_LC_18_12_7  (
            .in0(_gnd_net_),
            .in1(N__42396),
            .in2(_gnd_net_),
            .in3(N__40503),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_15 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_14 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_16_LC_18_13_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_16_LC_18_13_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_16_LC_18_13_0 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_16_LC_18_13_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__40782),
            .in3(N__40500),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_16 ),
            .ltout(),
            .carryin(bfn_18_13_0_),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_17_LC_18_13_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_17_LC_18_13_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_17_LC_18_13_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_17_LC_18_13_1  (
            .in0(_gnd_net_),
            .in1(N__41256),
            .in2(_gnd_net_),
            .in3(N__40497),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_17 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_16 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_18_LC_18_13_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNO_1_18_LC_18_13_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_18_LC_18_13_2 .LUT_INIT=16'b1000011101111000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_18_LC_18_13_2  (
            .in0(N__42259),
            .in1(N__42023),
            .in2(N__41652),
            .in3(N__40494),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.PPM_STATE_RNI78NT_0_LC_18_13_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_RNI78NT_0_LC_18_13_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.PPM_STATE_RNI78NT_0_LC_18_13_3 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \ppm_encoder_1.PPM_STATE_RNI78NT_0_LC_18_13_3  (
            .in0(N__40489),
            .in1(N__40421),
            .in2(N__40383),
            .in3(N__40326),
            .lcout(),
            .ltout(\ppm_encoder_1.init_pulses_0_sqmuxa_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNIRCE81_LC_18_13_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNIRCE81_LC_18_13_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNIRCE81_LC_18_13_4 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_57_c_RNIRCE81_LC_18_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__40275),
            .in3(N__44670),
            .lcout(\ppm_encoder_1.init_pulses_0_sqmuxa_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIGTUS_0_8_LC_18_13_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIGTUS_0_8_LC_18_13_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIGTUS_0_8_LC_18_13_7 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIGTUS_0_8_LC_18_13_7  (
            .in0(N__42022),
            .in1(N__40640),
            .in2(_gnd_net_),
            .in3(N__42258),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_7_LC_18_14_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_7_LC_18_14_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.init_pulses_7_LC_18_14_0 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_7_LC_18_14_0  (
            .in0(N__41599),
            .in1(N__40266),
            .in2(N__41473),
            .in3(N__40257),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47392),
            .ce(),
            .sr(N__43888));
    defparam \ppm_encoder_1.init_pulses_RNIFSUS_7_LC_18_14_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIFSUS_7_LC_18_14_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIFSUS_7_LC_18_14_1 .LUT_INIT=16'b0101101010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIFSUS_7_LC_18_14_1  (
            .in0(N__40708),
            .in1(_gnd_net_),
            .in2(N__42040),
            .in3(N__42248),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIFSUS_0_7_LC_18_14_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIFSUS_0_7_LC_18_14_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIFSUS_0_7_LC_18_14_2 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIFSUS_0_7_LC_18_14_2  (
            .in0(N__42247),
            .in1(N__42011),
            .in2(_gnd_net_),
            .in3(N__40709),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_7_LC_18_14_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_7_LC_18_14_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_7_LC_18_14_3 .LUT_INIT=16'b1110000000100000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_7_LC_18_14_3  (
            .in0(N__40710),
            .in1(N__40978),
            .in2(N__41121),
            .in3(N__40695),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_8_LC_18_14_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_8_LC_18_14_4 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_8_LC_18_14_4 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_8_LC_18_14_4  (
            .in0(N__41600),
            .in1(N__40659),
            .in2(N__41474),
            .in3(N__40650),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47392),
            .ce(),
            .sr(N__43888));
    defparam \ppm_encoder_1.init_pulses_RNIGTUS_8_LC_18_14_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIGTUS_8_LC_18_14_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIGTUS_8_LC_18_14_5 .LUT_INIT=16'b0101101010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIGTUS_8_LC_18_14_5  (
            .in0(N__40639),
            .in1(_gnd_net_),
            .in2(N__42041),
            .in3(N__42249),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_9_LC_18_15_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_9_LC_18_15_0 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_9_LC_18_15_0 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \ppm_encoder_1.init_pulses_9_LC_18_15_0  (
            .in0(N__41610),
            .in1(N__40599),
            .in2(N__41496),
            .in3(N__40593),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47377),
            .ce(),
            .sr(N__43893));
    defparam \ppm_encoder_1.init_pulses_RNIHUUS_0_9_LC_18_15_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIHUUS_0_9_LC_18_15_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIHUUS_0_9_LC_18_15_1 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIHUUS_0_9_LC_18_15_1  (
            .in0(N__42019),
            .in1(_gnd_net_),
            .in2(N__42284),
            .in3(N__40553),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIHUUS_9_LC_18_15_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIHUUS_9_LC_18_15_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIHUUS_9_LC_18_15_2 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIHUUS_9_LC_18_15_2  (
            .in0(N__40552),
            .in1(N__42254),
            .in2(_gnd_net_),
            .in3(N__42020),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_9_LC_18_15_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_9_LC_18_15_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_9_LC_18_15_3 .LUT_INIT=16'b1010000010001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_9_LC_18_15_3  (
            .in0(N__41094),
            .in1(N__40554),
            .in2(N__40542),
            .in3(N__40988),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNI0KRP_17_LC_18_15_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI0KRP_17_LC_18_15_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI0KRP_17_LC_18_15_5 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI0KRP_17_LC_18_15_5  (
            .in0(N__42021),
            .in1(_gnd_net_),
            .in2(N__42285),
            .in3(N__40741),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIPCRP_0_10_LC_18_15_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIPCRP_0_10_LC_18_15_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIPCRP_0_10_LC_18_15_6 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIPCRP_0_10_LC_18_15_6  (
            .in0(N__41242),
            .in1(N__42250),
            .in2(_gnd_net_),
            .in3(N__42018),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_14_LC_18_16_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_14_LC_18_16_0 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_14_LC_18_16_0 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_14_LC_18_16_0  (
            .in0(N__41612),
            .in1(N__41205),
            .in2(N__41497),
            .in3(N__41196),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47365),
            .ce(),
            .sr(N__43895));
    defparam \ppm_encoder_1.init_pulses_RNITGRP_14_LC_18_16_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNITGRP_14_LC_18_16_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNITGRP_14_LC_18_16_1 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNITGRP_14_LC_18_16_1  (
            .in0(N__41158),
            .in1(N__42272),
            .in2(_gnd_net_),
            .in3(N__41938),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNITGRP_0_14_LC_18_16_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNITGRP_0_14_LC_18_16_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNITGRP_0_14_LC_18_16_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNITGRP_0_14_LC_18_16_2  (
            .in0(N__41936),
            .in1(N__41159),
            .in2(_gnd_net_),
            .in3(N__42270),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_14_LC_18_16_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_14_LC_18_16_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_14_LC_18_16_3 .LUT_INIT=16'b1100000010001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_14_LC_18_16_3  (
            .in0(N__41160),
            .in1(N__41128),
            .in2(N__41025),
            .in3(N__40989),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_16_LC_18_16_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_16_LC_18_16_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.init_pulses_16_LC_18_16_4 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_16_LC_18_16_4  (
            .in0(N__41613),
            .in1(N__40824),
            .in2(N__41498),
            .in3(N__40815),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47365),
            .ce(),
            .sr(N__43895));
    defparam \ppm_encoder_1.init_pulses_RNIVIRP_16_LC_18_16_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIVIRP_16_LC_18_16_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIVIRP_16_LC_18_16_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIVIRP_16_LC_18_16_6  (
            .in0(N__41937),
            .in1(N__40799),
            .in2(_gnd_net_),
            .in3(N__42271),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_17_LC_18_16_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_17_LC_18_16_7 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_17_LC_18_16_7 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_17_LC_18_16_7  (
            .in0(N__41614),
            .in1(N__40770),
            .in2(N__41499),
            .in3(N__40761),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47365),
            .ce(),
            .sr(N__43895));
    defparam \ppm_encoder_1.init_pulses_RNI5ATG1_15_LC_18_17_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI5ATG1_15_LC_18_17_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI5ATG1_15_LC_18_17_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI5ATG1_15_LC_18_17_0  (
            .in0(N__42288),
            .in1(N__42361),
            .in2(N__42048),
            .in3(N__42346),
            .lcout(\ppm_encoder_1.init_pulses_RNI5ATG1Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIUHRP_15_LC_18_17_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIUHRP_15_LC_18_17_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIUHRP_15_LC_18_17_1 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIUHRP_15_LC_18_17_1  (
            .in0(N__42362),
            .in1(N__42286),
            .in2(_gnd_net_),
            .in3(N__42042),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_15_LC_18_17_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_15_LC_18_17_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.init_pulses_15_LC_18_17_2 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_15_LC_18_17_2  (
            .in0(N__41608),
            .in1(N__42387),
            .in2(N__41501),
            .in3(N__42378),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47351),
            .ce(),
            .sr(N__43896));
    defparam \ppm_encoder_1.init_pulses_RNO_2_18_LC_18_17_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNO_2_18_LC_18_17_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_2_18_LC_18_17_3 .LUT_INIT=16'b1001011001011010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_2_18_LC_18_17_3  (
            .in0(N__42347),
            .in1(N__42287),
            .in2(N__41641),
            .in3(N__42043),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_axb_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_18_LC_18_17_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_18_LC_18_17_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.init_pulses_18_LC_18_17_4 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_18_LC_18_17_4  (
            .in0(N__41609),
            .in1(N__41667),
            .in2(N__41502),
            .in3(N__41658),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47351),
            .ce(),
            .sr(N__43896));
    defparam \ppm_encoder_1.init_pulses_13_LC_18_17_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_13_LC_18_17_6 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_13_LC_18_17_6 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_13_LC_18_17_6  (
            .in0(N__41607),
            .in1(N__41514),
            .in2(N__41500),
            .in3(N__41346),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47351),
            .ce(),
            .sr(N__43896));
    defparam \ppm_encoder_1.pulses2count_esr_14_LC_18_18_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_14_LC_18_18_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_14_LC_18_18_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_14_LC_18_18_0  (
            .in0(N__42605),
            .in1(N__41307),
            .in2(_gnd_net_),
            .in3(N__41298),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47335),
            .ce(N__42539),
            .sr(N__43898));
    defparam \ppm_encoder_1.pulses2count_esr_10_LC_18_18_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_10_LC_18_18_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_10_LC_18_18_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_10_LC_18_18_4  (
            .in0(N__42604),
            .in1(N__41280),
            .in2(_gnd_net_),
            .in3(N__41268),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47335),
            .ce(N__42539),
            .sr(N__43898));
    defparam \ppm_encoder_1.pulses2count_esr_7_LC_18_18_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_7_LC_18_18_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_7_LC_18_18_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_7_LC_18_18_7  (
            .in0(N__42762),
            .in1(N__42606),
            .in2(_gnd_net_),
            .in3(N__42750),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47335),
            .ce(N__42539),
            .sr(N__43898));
    defparam \ppm_encoder_1.counter24_0_I_21_c_RNO_LC_18_19_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_21_c_RNO_LC_18_19_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_21_c_RNO_LC_18_19_0 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_21_c_RNO_LC_18_19_0  (
            .in0(N__42736),
            .in1(N__42660),
            .in2(N__42717),
            .in3(N__42707),
            .lcout(\ppm_encoder_1.counter24_0_I_21_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_6_LC_18_19_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_6_LC_18_19_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_6_LC_18_19_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_6_LC_18_19_1  (
            .in0(N__42616),
            .in1(N__42687),
            .in2(_gnd_net_),
            .in3(N__42672),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47322),
            .ce(N__42538),
            .sr(N__43901));
    defparam \ppm_encoder_1.pulses2count_esr_11_LC_18_19_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_11_LC_18_19_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_11_LC_18_19_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_11_LC_18_19_3  (
            .in0(N__42612),
            .in1(N__42654),
            .in2(_gnd_net_),
            .in3(N__42642),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47322),
            .ce(N__42538),
            .sr(N__43901));
    defparam \ppm_encoder_1.pulses2count_esr_12_LC_18_19_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_12_LC_18_19_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_12_LC_18_19_5 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_12_LC_18_19_5  (
            .in0(N__42630),
            .in1(_gnd_net_),
            .in2(N__42618),
            .in3(N__42555),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47322),
            .ce(N__42538),
            .sr(N__43901));
    defparam \ppm_encoder_1.counter24_0_I_39_c_RNO_LC_18_19_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_39_c_RNO_LC_18_19_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_39_c_RNO_LC_18_19_6 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_39_c_RNO_LC_18_19_6  (
            .in0(N__42489),
            .in1(N__42465),
            .in2(N__42459),
            .in3(N__42450),
            .lcout(\ppm_encoder_1.counter24_0_I_39_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_1_c_LC_18_20_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_1_c_LC_18_20_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_1_c_LC_18_20_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_1_c_LC_18_20_0  (
            .in0(_gnd_net_),
            .in1(N__42426),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_18_20_0_),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_9_c_LC_18_20_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_9_c_LC_18_20_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_9_c_LC_18_20_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_9_c_LC_18_20_1  (
            .in0(_gnd_net_),
            .in1(N__43008),
            .in2(N__42417),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ppm_encoder_1.counter24_0_data_tmp_0 ),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_15_c_LC_18_20_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_15_c_LC_18_20_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_15_c_LC_18_20_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_15_c_LC_18_20_2  (
            .in0(_gnd_net_),
            .in1(N__43191),
            .in2(N__43068),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ppm_encoder_1.counter24_0_data_tmp_1 ),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_21_c_LC_18_20_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_21_c_LC_18_20_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_21_c_LC_18_20_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_21_c_LC_18_20_3  (
            .in0(_gnd_net_),
            .in1(N__42999),
            .in2(N__43179),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ppm_encoder_1.counter24_0_data_tmp_2 ),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_27_c_LC_18_20_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_27_c_LC_18_20_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_27_c_LC_18_20_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_27_c_LC_18_20_4  (
            .in0(_gnd_net_),
            .in1(N__43167),
            .in2(N__43069),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ppm_encoder_1.counter24_0_data_tmp_3 ),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_33_c_LC_18_20_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_33_c_LC_18_20_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_33_c_LC_18_20_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_33_c_LC_18_20_5  (
            .in0(_gnd_net_),
            .in1(N__43003),
            .in2(N__44565),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ppm_encoder_1.counter24_0_data_tmp_4 ),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_39_c_LC_18_20_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_39_c_LC_18_20_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_39_c_LC_18_20_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_39_c_LC_18_20_6  (
            .in0(_gnd_net_),
            .in1(N__43161),
            .in2(N__43070),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ppm_encoder_1.counter24_0_data_tmp_5 ),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_45_c_LC_18_20_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_45_c_LC_18_20_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_45_c_LC_18_20_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_45_c_LC_18_20_7  (
            .in0(_gnd_net_),
            .in1(N__43007),
            .in2(N__43155),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ppm_encoder_1.counter24_0_data_tmp_6 ),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_51_c_LC_18_21_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_51_c_LC_18_21_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_51_c_LC_18_21_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_51_c_LC_18_21_0  (
            .in0(_gnd_net_),
            .in1(N__43146),
            .in2(N__43118),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_18_21_0_),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_57_c_LC_18_21_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_57_c_LC_18_21_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_57_c_LC_18_21_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_57_c_LC_18_21_1  (
            .in0(_gnd_net_),
            .in1(N__43074),
            .in2(N__42771),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ppm_encoder_1.counter24_0_data_tmp_8 ),
            .carryout(\ppm_encoder_1.counter24_0_N_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_N_2_THRU_LUT4_0_LC_18_21_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_N_2_THRU_LUT4_0_LC_18_21_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_N_2_THRU_LUT4_0_LC_18_21_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.counter24_0_N_2_THRU_LUT4_0_LC_18_21_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44673),
            .lcout(\ppm_encoder_1.counter24_0_N_2_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_33_c_RNO_LC_18_21_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_33_c_RNO_LC_18_21_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_33_c_RNO_LC_18_21_3 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_33_c_RNO_LC_18_21_3  (
            .in0(N__44634),
            .in1(N__44625),
            .in2(N__44601),
            .in3(N__44589),
            .lcout(\ppm_encoder_1.counter24_0_I_33_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.bit_Count_0_LC_20_8_1 .C_ON=1'b0;
    defparam \uart_drone.bit_Count_0_LC_20_8_1 .SEQ_MODE=4'b1000;
    defparam \uart_drone.bit_Count_0_LC_20_8_1 .LUT_INIT=16'b0000110000101100;
    LogicCell40 \uart_drone.bit_Count_0_LC_20_8_1  (
            .in0(N__44556),
            .in1(N__44378),
            .in2(N__44499),
            .in3(N__44469),
            .lcout(\uart_drone.bit_CountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47465),
            .ce(),
            .sr(N__43862));
    defparam \pid_alt.error_filt_prev_esr_21_LC_20_10_1 .C_ON=1'b0;
    defparam \pid_alt.error_filt_prev_esr_21_LC_20_10_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_filt_prev_esr_21_LC_20_10_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_filt_prev_esr_21_LC_20_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44343),
            .lcout(\pid_alt.error_filt_prevZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47453),
            .ce(N__46819),
            .sr(N__46600));
    defparam \Commands_frame_decoder.source_alt_ki_5_LC_20_23_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_ki_5_LC_20_23_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_ki_5_LC_20_23_7 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_ki_5_LC_20_23_7  (
            .in0(_gnd_net_),
            .in1(N__44283),
            .in2(_gnd_net_),
            .in3(N__46675),
            .lcout(alt_ki_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47303),
            .ce(N__44865),
            .sr(_gnd_net_));
    defparam GB_BUFFER_reset_system_g_THRU_LUT4_0_LC_20_30_0.C_ON=1'b0;
    defparam GB_BUFFER_reset_system_g_THRU_LUT4_0_LC_20_30_0.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_reset_system_g_THRU_LUT4_0_LC_20_30_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 GB_BUFFER_reset_system_g_THRU_LUT4_0_LC_20_30_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44065),
            .lcout(GB_BUFFER_reset_system_g_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_ki_3_LC_21_20_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_ki_3_LC_21_20_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_ki_3_LC_21_20_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_ki_3_LC_21_20_2  (
            .in0(_gnd_net_),
            .in1(N__43364),
            .in2(_gnd_net_),
            .in3(N__46680),
            .lcout(alt_ki_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47353),
            .ce(N__44860),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_reg_esr_4_LC_21_21_2 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_4_LC_21_21_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_4_LC_21_21_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_4_LC_21_21_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43218),
            .lcout(\pid_alt.error_i_regZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47337),
            .ce(N__46806),
            .sr(N__46589));
    defparam \pid_alt.error_i_reg_esr_5_LC_21_21_7 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_5_LC_21_21_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_5_LC_21_21_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_5_LC_21_21_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45420),
            .lcout(\pid_alt.error_i_regZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47337),
            .ce(N__46806),
            .sr(N__46589));
    defparam \pid_alt.error_i_reg_esr_8_LC_21_22_0 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_8_LC_21_22_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_8_LC_21_22_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_8_LC_21_22_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45396),
            .lcout(\pid_alt.error_i_regZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47324),
            .ce(N__46802),
            .sr(N__46587));
    defparam \Commands_frame_decoder.source_alt_ki_4_LC_21_23_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_ki_4_LC_21_23_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_ki_4_LC_21_23_2 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Commands_frame_decoder.source_alt_ki_4_LC_21_23_2  (
            .in0(N__46677),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45366),
            .lcout(alt_ki_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47312),
            .ce(N__44856),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_ki_1_LC_21_23_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_ki_1_LC_21_23_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_ki_1_LC_21_23_5 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_ki_1_LC_21_23_5  (
            .in0(_gnd_net_),
            .in1(N__45224),
            .in2(_gnd_net_),
            .in3(N__46676),
            .lcout(alt_ki_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47312),
            .ce(N__44856),
            .sr(_gnd_net_));
    defparam \pid_alt.error_filt_prev_esr_19_LC_22_10_4 .C_ON=1'b0;
    defparam \pid_alt.error_filt_prev_esr_19_LC_22_10_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_filt_prev_esr_19_LC_22_10_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_filt_prev_esr_19_LC_22_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45066),
            .lcout(\pid_alt.error_filt_prevZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47466),
            .ce(N__46822),
            .sr(N__46604));
    defparam \Commands_frame_decoder.source_alt_ki_7_LC_22_22_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_ki_7_LC_22_22_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_ki_7_LC_22_22_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_ki_7_LC_22_22_2  (
            .in0(_gnd_net_),
            .in1(N__45013),
            .in2(_gnd_net_),
            .in3(N__46679),
            .lcout(alt_ki_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47338),
            .ce(N__44864),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_reg_esr_10_LC_22_23_1 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_10_LC_22_23_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_10_LC_22_23_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_10_LC_22_23_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44772),
            .lcout(\pid_alt.error_i_regZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47325),
            .ce(N__46803),
            .sr(N__46588));
    defparam \pid_alt.error_i_reg_esr_11_LC_23_23_0 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_11_LC_23_23_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_11_LC_23_23_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_11_LC_23_23_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44739),
            .lcout(\pid_alt.error_i_regZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47339),
            .ce(N__46807),
            .sr(N__46590));
    defparam \pid_alt.error_i_reg_esr_12_LC_23_23_1 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_12_LC_23_23_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_12_LC_23_23_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_12_LC_23_23_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44706),
            .lcout(\pid_alt.error_i_regZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47339),
            .ce(N__46807),
            .sr(N__46590));
    defparam \pid_alt.error_i_reg_esr_13_LC_23_23_4 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_13_LC_23_23_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_13_LC_23_23_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_13_LC_23_23_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45831),
            .lcout(\pid_alt.error_i_regZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47339),
            .ce(N__46807),
            .sr(N__46590));
    defparam \pid_alt.error_filt_prev_esr_17_LC_24_10_0 .C_ON=1'b0;
    defparam \pid_alt.error_filt_prev_esr_17_LC_24_10_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_filt_prev_esr_17_LC_24_10_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_filt_prev_esr_17_LC_24_10_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45798),
            .lcout(\pid_alt.error_filt_prevZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47473),
            .ce(N__46824),
            .sr(N__46611));
    defparam \pid_alt.error_filt_prev_esr_18_LC_24_10_1 .C_ON=1'b0;
    defparam \pid_alt.error_filt_prev_esr_18_LC_24_10_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_filt_prev_esr_18_LC_24_10_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_filt_prev_esr_18_LC_24_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45750),
            .lcout(\pid_alt.error_filt_prevZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47473),
            .ce(N__46824),
            .sr(N__46611));
    defparam \pid_alt.error_filt_prev_esr_22_LC_24_10_2 .C_ON=1'b0;
    defparam \pid_alt.error_filt_prev_esr_22_LC_24_10_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_filt_prev_esr_22_LC_24_10_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_filt_prev_esr_22_LC_24_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45702),
            .lcout(\pid_alt.error_filt_prevZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47473),
            .ce(N__46824),
            .sr(N__46611));
    defparam \pid_alt.error_filt_prev_esr_20_LC_24_11_1 .C_ON=1'b0;
    defparam \pid_alt.error_filt_prev_esr_20_LC_24_11_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_filt_prev_esr_20_LC_24_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_filt_prev_esr_20_LC_24_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45600),
            .lcout(\pid_alt.error_filt_prevZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47471),
            .ce(N__46823),
            .sr(N__46607));
    defparam \pid_alt.error_filt_prev_esr_8_LC_24_13_6 .C_ON=1'b0;
    defparam \pid_alt.error_filt_prev_esr_8_LC_24_13_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_filt_prev_esr_8_LC_24_13_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_filt_prev_esr_8_LC_24_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45561),
            .lcout(\pid_alt.error_filt_prevZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47460),
            .ce(N__46821),
            .sr(N__46603));
    defparam \pid_alt.error_d_reg_esr_4_LC_24_14_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_4_LC_24_14_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_4_LC_24_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_4_LC_24_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45522),
            .lcout(\pid_alt.error_d_regZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47454),
            .ce(N__46820),
            .sr(N__46601));
    defparam \pid_alt.error_filt_prev_esr_1_LC_24_14_4 .C_ON=1'b0;
    defparam \pid_alt.error_filt_prev_esr_1_LC_24_14_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_filt_prev_esr_1_LC_24_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_filt_prev_esr_1_LC_24_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45462),
            .lcout(\pid_alt.error_filt_prevZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47454),
            .ce(N__46820),
            .sr(N__46601));
    defparam \pid_alt.error_filt_prev_esr_2_LC_24_14_5 .C_ON=1'b0;
    defparam \pid_alt.error_filt_prev_esr_2_LC_24_14_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_filt_prev_esr_2_LC_24_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_filt_prev_esr_2_LC_24_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46176),
            .lcout(\pid_alt.error_filt_prevZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47454),
            .ce(N__46820),
            .sr(N__46601));
    defparam \pid_alt.error_filt_prev_esr_10_LC_24_15_0 .C_ON=1'b0;
    defparam \pid_alt.error_filt_prev_esr_10_LC_24_15_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_filt_prev_esr_10_LC_24_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_filt_prev_esr_10_LC_24_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46140),
            .lcout(\pid_alt.error_filt_prevZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47446),
            .ce(N__46818),
            .sr(N__46599));
    defparam \pid_alt.error_filt_prev_esr_11_LC_24_15_2 .C_ON=1'b0;
    defparam \pid_alt.error_filt_prev_esr_11_LC_24_15_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_filt_prev_esr_11_LC_24_15_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_filt_prev_esr_11_LC_24_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46104),
            .lcout(\pid_alt.error_filt_prevZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47446),
            .ce(N__46818),
            .sr(N__46599));
    defparam \pid_alt.error_filt_prev_esr_12_LC_24_15_3 .C_ON=1'b0;
    defparam \pid_alt.error_filt_prev_esr_12_LC_24_15_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_filt_prev_esr_12_LC_24_15_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_filt_prev_esr_12_LC_24_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46062),
            .lcout(\pid_alt.error_filt_prevZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47446),
            .ce(N__46818),
            .sr(N__46599));
    defparam \pid_alt.error_filt_prev_esr_13_LC_24_15_5 .C_ON=1'b0;
    defparam \pid_alt.error_filt_prev_esr_13_LC_24_15_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_filt_prev_esr_13_LC_24_15_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_filt_prev_esr_13_LC_24_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46023),
            .lcout(\pid_alt.error_filt_prevZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47446),
            .ce(N__46818),
            .sr(N__46599));
    defparam \pid_alt.error_filt_prev_esr_15_LC_24_15_6 .C_ON=1'b0;
    defparam \pid_alt.error_filt_prev_esr_15_LC_24_15_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_filt_prev_esr_15_LC_24_15_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_filt_prev_esr_15_LC_24_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45987),
            .lcout(\pid_alt.error_filt_prevZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47446),
            .ce(N__46818),
            .sr(N__46599));
    defparam \pid_alt.error_filt_prev_esr_16_LC_24_15_7 .C_ON=1'b0;
    defparam \pid_alt.error_filt_prev_esr_16_LC_24_15_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_filt_prev_esr_16_LC_24_15_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_filt_prev_esr_16_LC_24_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45942),
            .lcout(\pid_alt.error_filt_prevZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47446),
            .ce(N__46818),
            .sr(N__46599));
    defparam \pid_alt.error_filt_prev_esr_4_LC_24_16_0 .C_ON=1'b0;
    defparam \pid_alt.error_filt_prev_esr_4_LC_24_16_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_filt_prev_esr_4_LC_24_16_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_filt_prev_esr_4_LC_24_16_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45894),
            .lcout(\pid_alt.error_filt_prevZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47439),
            .ce(N__46817),
            .sr(N__46597));
    defparam \pid_alt.error_filt_prev_esr_5_LC_24_16_1 .C_ON=1'b0;
    defparam \pid_alt.error_filt_prev_esr_5_LC_24_16_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_filt_prev_esr_5_LC_24_16_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_filt_prev_esr_5_LC_24_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45864),
            .lcout(\pid_alt.error_filt_prevZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47439),
            .ce(N__46817),
            .sr(N__46597));
    defparam \pid_alt.error_filt_prev_esr_6_LC_24_16_2 .C_ON=1'b0;
    defparam \pid_alt.error_filt_prev_esr_6_LC_24_16_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_filt_prev_esr_6_LC_24_16_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_filt_prev_esr_6_LC_24_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46425),
            .lcout(\pid_alt.error_filt_prevZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47439),
            .ce(N__46817),
            .sr(N__46597));
    defparam \pid_alt.error_filt_prev_esr_7_LC_24_16_3 .C_ON=1'b0;
    defparam \pid_alt.error_filt_prev_esr_7_LC_24_16_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_filt_prev_esr_7_LC_24_16_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_filt_prev_esr_7_LC_24_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46392),
            .lcout(\pid_alt.error_filt_prevZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47439),
            .ce(N__46817),
            .sr(N__46597));
    defparam \pid_alt.error_filt_prev_esr_9_LC_24_16_5 .C_ON=1'b0;
    defparam \pid_alt.error_filt_prev_esr_9_LC_24_16_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_filt_prev_esr_9_LC_24_16_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_filt_prev_esr_9_LC_24_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46359),
            .lcout(\pid_alt.error_filt_prevZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47439),
            .ce(N__46817),
            .sr(N__46597));
    defparam \pid_alt.error_filt_prev_esr_3_LC_24_16_7 .C_ON=1'b0;
    defparam \pid_alt.error_filt_prev_esr_3_LC_24_16_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_filt_prev_esr_3_LC_24_16_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_filt_prev_esr_3_LC_24_16_7  (
            .in0(N__46314),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_filt_prevZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47439),
            .ce(N__46817),
            .sr(N__46597));
    defparam \pid_alt.error_filt_prev_esr_14_LC_24_17_5 .C_ON=1'b0;
    defparam \pid_alt.error_filt_prev_esr_14_LC_24_17_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_filt_prev_esr_14_LC_24_17_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_filt_prev_esr_14_LC_24_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46281),
            .lcout(\pid_alt.error_filt_prevZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47429),
            .ce(N__46816),
            .sr(N__46596));
    defparam \pid_alt.error_i_reg_esr_7_LC_24_21_2 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_7_LC_24_21_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_7_LC_24_21_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_i_reg_esr_7_LC_24_21_2  (
            .in0(N__46248),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_i_regZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47379),
            .ce(N__46813),
            .sr(N__46595));
    defparam \pid_alt.error_i_reg_esr_6_LC_24_21_4 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_6_LC_24_21_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_6_LC_24_21_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_i_reg_esr_6_LC_24_21_4  (
            .in0(N__46224),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_i_regZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47379),
            .ce(N__46813),
            .sr(N__46595));
    defparam \pid_alt.error_i_reg_esr_15_LC_24_22_1 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_15_LC_24_22_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_15_LC_24_22_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_15_LC_24_22_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46203),
            .lcout(\pid_alt.error_i_regZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47367),
            .ce(N__46811),
            .sr(N__46594));
    defparam \pid_alt.error_i_reg_esr_9_LC_24_22_3 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_9_LC_24_22_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_9_LC_24_22_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_9_LC_24_22_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47625),
            .lcout(\pid_alt.error_i_regZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47367),
            .ce(N__46811),
            .sr(N__46594));
    defparam \pid_alt.error_i_reg_esr_14_LC_24_22_7 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_14_LC_24_22_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_14_LC_24_22_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_14_LC_24_22_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47604),
            .lcout(\pid_alt.error_i_regZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47367),
            .ce(N__46811),
            .sr(N__46594));
    defparam \pid_alt.error_i_reg_esr_20_LC_24_23_0 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_20_LC_24_23_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_20_LC_24_23_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_20_LC_24_23_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47586),
            .lcout(\pid_alt.error_i_regZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47354),
            .ce(N__46810),
            .sr(N__46592));
    defparam \pid_alt.error_i_reg_esr_17_LC_24_23_4 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_17_LC_24_23_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_17_LC_24_23_4 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \pid_alt.error_i_reg_esr_17_LC_24_23_4  (
            .in0(_gnd_net_),
            .in1(N__47562),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_i_regZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47354),
            .ce(N__46810),
            .sr(N__46592));
    defparam \pid_alt.error_i_reg_esr_18_LC_24_23_6 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_18_LC_24_23_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_18_LC_24_23_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_i_reg_esr_18_LC_24_23_6  (
            .in0(N__47541),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_i_regZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47354),
            .ce(N__46810),
            .sr(N__46592));
    defparam \pid_alt.error_i_reg_esr_16_LC_24_23_7 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_16_LC_24_23_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_16_LC_24_23_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_16_LC_24_23_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47520),
            .lcout(\pid_alt.error_i_regZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47354),
            .ce(N__46810),
            .sr(N__46592));
    defparam \pid_alt.error_i_reg_esr_19_LC_24_24_2 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_19_LC_24_24_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_19_LC_24_24_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_19_LC_24_24_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47502),
            .lcout(\pid_alt.error_i_regZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47340),
            .ce(N__46808),
            .sr(N__46591));
endmodule // Pc2drone
