// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 11 2017 17:30:03

// File Generated:     Jun 2 2019 13:25:24

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "Pc2drone" view "INTERFACE"

module Pc2drone (
    uart_input_pc,
    debug_CH5_31B,
    debug_CH3_20A,
    debug_CH0_16A,
    uart_input_drone,
    ppm_output,
    debug_CH6_5B,
    debug_CH2_18A,
    debug_CH4_2A,
    debug_CH1_0A,
    clk_system);

    input uart_input_pc;
    output debug_CH5_31B;
    output debug_CH3_20A;
    output debug_CH0_16A;
    input uart_input_drone;
    output ppm_output;
    output debug_CH6_5B;
    output debug_CH2_18A;
    output debug_CH4_2A;
    output debug_CH1_0A;
    input clk_system;

    wire N__87702;
    wire N__87688;
    wire N__87687;
    wire N__87686;
    wire N__87679;
    wire N__87678;
    wire N__87677;
    wire N__87670;
    wire N__87669;
    wire N__87668;
    wire N__87661;
    wire N__87660;
    wire N__87659;
    wire N__87652;
    wire N__87651;
    wire N__87650;
    wire N__87643;
    wire N__87642;
    wire N__87641;
    wire N__87634;
    wire N__87633;
    wire N__87632;
    wire N__87625;
    wire N__87624;
    wire N__87623;
    wire N__87616;
    wire N__87615;
    wire N__87614;
    wire N__87607;
    wire N__87606;
    wire N__87605;
    wire N__87588;
    wire N__87585;
    wire N__87582;
    wire N__87579;
    wire N__87578;
    wire N__87577;
    wire N__87570;
    wire N__87567;
    wire N__87564;
    wire N__87561;
    wire N__87558;
    wire N__87555;
    wire N__87552;
    wire N__87549;
    wire N__87546;
    wire N__87545;
    wire N__87540;
    wire N__87539;
    wire N__87536;
    wire N__87533;
    wire N__87530;
    wire N__87527;
    wire N__87524;
    wire N__87521;
    wire N__87516;
    wire N__87513;
    wire N__87510;
    wire N__87507;
    wire N__87504;
    wire N__87503;
    wire N__87502;
    wire N__87499;
    wire N__87494;
    wire N__87491;
    wire N__87488;
    wire N__87485;
    wire N__87482;
    wire N__87477;
    wire N__87474;
    wire N__87471;
    wire N__87468;
    wire N__87465;
    wire N__87464;
    wire N__87463;
    wire N__87460;
    wire N__87455;
    wire N__87450;
    wire N__87447;
    wire N__87444;
    wire N__87441;
    wire N__87438;
    wire N__87435;
    wire N__87432;
    wire N__87429;
    wire N__87426;
    wire N__87425;
    wire N__87424;
    wire N__87423;
    wire N__87422;
    wire N__87421;
    wire N__87420;
    wire N__87419;
    wire N__87418;
    wire N__87417;
    wire N__87416;
    wire N__87415;
    wire N__87414;
    wire N__87409;
    wire N__87404;
    wire N__87403;
    wire N__87398;
    wire N__87389;
    wire N__87382;
    wire N__87379;
    wire N__87376;
    wire N__87373;
    wire N__87366;
    wire N__87363;
    wire N__87360;
    wire N__87355;
    wire N__87352;
    wire N__87347;
    wire N__87344;
    wire N__87341;
    wire N__87338;
    wire N__87333;
    wire N__87330;
    wire N__87327;
    wire N__87324;
    wire N__87323;
    wire N__87322;
    wire N__87315;
    wire N__87312;
    wire N__87309;
    wire N__87306;
    wire N__87303;
    wire N__87300;
    wire N__87297;
    wire N__87296;
    wire N__87295;
    wire N__87288;
    wire N__87285;
    wire N__87282;
    wire N__87279;
    wire N__87278;
    wire N__87277;
    wire N__87276;
    wire N__87275;
    wire N__87274;
    wire N__87273;
    wire N__87272;
    wire N__87271;
    wire N__87270;
    wire N__87269;
    wire N__87268;
    wire N__87267;
    wire N__87266;
    wire N__87265;
    wire N__87264;
    wire N__87263;
    wire N__87262;
    wire N__87261;
    wire N__87260;
    wire N__87259;
    wire N__87258;
    wire N__87257;
    wire N__87256;
    wire N__87255;
    wire N__87254;
    wire N__87253;
    wire N__87252;
    wire N__87251;
    wire N__87250;
    wire N__87249;
    wire N__87248;
    wire N__87247;
    wire N__87246;
    wire N__87245;
    wire N__87244;
    wire N__87243;
    wire N__87242;
    wire N__87241;
    wire N__87240;
    wire N__87239;
    wire N__87238;
    wire N__87237;
    wire N__87236;
    wire N__87235;
    wire N__87234;
    wire N__87233;
    wire N__87232;
    wire N__87231;
    wire N__87230;
    wire N__87229;
    wire N__87228;
    wire N__87227;
    wire N__87226;
    wire N__87225;
    wire N__87224;
    wire N__87223;
    wire N__87222;
    wire N__87221;
    wire N__87220;
    wire N__87219;
    wire N__87218;
    wire N__87217;
    wire N__87216;
    wire N__87215;
    wire N__87214;
    wire N__87213;
    wire N__87212;
    wire N__87211;
    wire N__87210;
    wire N__87209;
    wire N__87208;
    wire N__87207;
    wire N__87206;
    wire N__87205;
    wire N__87204;
    wire N__87203;
    wire N__87202;
    wire N__87201;
    wire N__87200;
    wire N__87199;
    wire N__87198;
    wire N__87197;
    wire N__87196;
    wire N__87195;
    wire N__87194;
    wire N__87193;
    wire N__87192;
    wire N__87191;
    wire N__87190;
    wire N__87189;
    wire N__87188;
    wire N__87187;
    wire N__87186;
    wire N__87185;
    wire N__87184;
    wire N__87183;
    wire N__87182;
    wire N__87181;
    wire N__87180;
    wire N__87179;
    wire N__87178;
    wire N__87177;
    wire N__87176;
    wire N__87175;
    wire N__87174;
    wire N__87173;
    wire N__87172;
    wire N__87171;
    wire N__87170;
    wire N__87169;
    wire N__87168;
    wire N__87167;
    wire N__87166;
    wire N__87165;
    wire N__87164;
    wire N__87163;
    wire N__87162;
    wire N__87161;
    wire N__87160;
    wire N__87159;
    wire N__87158;
    wire N__87157;
    wire N__87156;
    wire N__87155;
    wire N__87154;
    wire N__87153;
    wire N__87152;
    wire N__87151;
    wire N__87150;
    wire N__87149;
    wire N__87148;
    wire N__87147;
    wire N__87146;
    wire N__87145;
    wire N__87144;
    wire N__87143;
    wire N__87142;
    wire N__87141;
    wire N__87140;
    wire N__87139;
    wire N__87138;
    wire N__87137;
    wire N__87136;
    wire N__87135;
    wire N__87134;
    wire N__87133;
    wire N__87132;
    wire N__87131;
    wire N__87130;
    wire N__87129;
    wire N__87128;
    wire N__87127;
    wire N__87126;
    wire N__87125;
    wire N__87124;
    wire N__87123;
    wire N__87122;
    wire N__87121;
    wire N__87120;
    wire N__87119;
    wire N__87118;
    wire N__87117;
    wire N__87116;
    wire N__87115;
    wire N__87114;
    wire N__87113;
    wire N__87112;
    wire N__87111;
    wire N__87110;
    wire N__87109;
    wire N__87108;
    wire N__87107;
    wire N__87106;
    wire N__87105;
    wire N__87104;
    wire N__87103;
    wire N__87102;
    wire N__87101;
    wire N__87100;
    wire N__87099;
    wire N__87098;
    wire N__87097;
    wire N__87096;
    wire N__87095;
    wire N__87094;
    wire N__87093;
    wire N__87092;
    wire N__87091;
    wire N__87090;
    wire N__87089;
    wire N__87088;
    wire N__87087;
    wire N__87086;
    wire N__87085;
    wire N__87084;
    wire N__87083;
    wire N__87082;
    wire N__87081;
    wire N__87080;
    wire N__87079;
    wire N__87078;
    wire N__87077;
    wire N__87076;
    wire N__87075;
    wire N__87074;
    wire N__87073;
    wire N__87072;
    wire N__87071;
    wire N__87070;
    wire N__87069;
    wire N__87068;
    wire N__87067;
    wire N__87066;
    wire N__87065;
    wire N__87064;
    wire N__87063;
    wire N__87062;
    wire N__87061;
    wire N__87060;
    wire N__87059;
    wire N__87058;
    wire N__87057;
    wire N__87056;
    wire N__87055;
    wire N__87054;
    wire N__87053;
    wire N__87052;
    wire N__87051;
    wire N__87050;
    wire N__87049;
    wire N__87048;
    wire N__87047;
    wire N__87046;
    wire N__87045;
    wire N__87044;
    wire N__87043;
    wire N__87042;
    wire N__87041;
    wire N__87040;
    wire N__87039;
    wire N__87038;
    wire N__87037;
    wire N__87036;
    wire N__87035;
    wire N__87034;
    wire N__87033;
    wire N__87032;
    wire N__87031;
    wire N__87030;
    wire N__87029;
    wire N__87028;
    wire N__87027;
    wire N__87026;
    wire N__87025;
    wire N__87024;
    wire N__87023;
    wire N__87022;
    wire N__87021;
    wire N__87020;
    wire N__87019;
    wire N__87018;
    wire N__87017;
    wire N__87016;
    wire N__87015;
    wire N__87014;
    wire N__87013;
    wire N__87012;
    wire N__87011;
    wire N__87010;
    wire N__87009;
    wire N__87008;
    wire N__87007;
    wire N__87006;
    wire N__87005;
    wire N__87004;
    wire N__87003;
    wire N__87002;
    wire N__87001;
    wire N__87000;
    wire N__86999;
    wire N__86998;
    wire N__86997;
    wire N__86996;
    wire N__86995;
    wire N__86994;
    wire N__86993;
    wire N__86992;
    wire N__86991;
    wire N__86990;
    wire N__86989;
    wire N__86988;
    wire N__86987;
    wire N__86986;
    wire N__86985;
    wire N__86984;
    wire N__86983;
    wire N__86982;
    wire N__86981;
    wire N__86980;
    wire N__86979;
    wire N__86978;
    wire N__86977;
    wire N__86976;
    wire N__86975;
    wire N__86974;
    wire N__86973;
    wire N__86972;
    wire N__86971;
    wire N__86970;
    wire N__86969;
    wire N__86346;
    wire N__86343;
    wire N__86340;
    wire N__86339;
    wire N__86338;
    wire N__86337;
    wire N__86336;
    wire N__86333;
    wire N__86330;
    wire N__86329;
    wire N__86326;
    wire N__86323;
    wire N__86320;
    wire N__86319;
    wire N__86318;
    wire N__86317;
    wire N__86314;
    wire N__86311;
    wire N__86308;
    wire N__86307;
    wire N__86304;
    wire N__86299;
    wire N__86296;
    wire N__86293;
    wire N__86292;
    wire N__86289;
    wire N__86288;
    wire N__86283;
    wire N__86280;
    wire N__86277;
    wire N__86276;
    wire N__86269;
    wire N__86266;
    wire N__86263;
    wire N__86260;
    wire N__86257;
    wire N__86252;
    wire N__86249;
    wire N__86246;
    wire N__86243;
    wire N__86240;
    wire N__86237;
    wire N__86232;
    wire N__86225;
    wire N__86222;
    wire N__86219;
    wire N__86216;
    wire N__86213;
    wire N__86210;
    wire N__86207;
    wire N__86204;
    wire N__86197;
    wire N__86190;
    wire N__86189;
    wire N__86188;
    wire N__86187;
    wire N__86186;
    wire N__86185;
    wire N__86184;
    wire N__86183;
    wire N__86182;
    wire N__86181;
    wire N__86180;
    wire N__86179;
    wire N__86178;
    wire N__86177;
    wire N__86176;
    wire N__86175;
    wire N__86174;
    wire N__86173;
    wire N__86172;
    wire N__86171;
    wire N__86170;
    wire N__86169;
    wire N__86168;
    wire N__86167;
    wire N__86166;
    wire N__86165;
    wire N__86164;
    wire N__86163;
    wire N__86162;
    wire N__86161;
    wire N__86160;
    wire N__86159;
    wire N__86158;
    wire N__86157;
    wire N__86156;
    wire N__86155;
    wire N__86154;
    wire N__86153;
    wire N__86152;
    wire N__86151;
    wire N__86150;
    wire N__86149;
    wire N__86148;
    wire N__86137;
    wire N__86134;
    wire N__86129;
    wire N__86112;
    wire N__86107;
    wire N__86092;
    wire N__86089;
    wire N__86080;
    wire N__86077;
    wire N__86072;
    wire N__86069;
    wire N__86064;
    wire N__86061;
    wire N__86058;
    wire N__86055;
    wire N__86052;
    wire N__86045;
    wire N__86044;
    wire N__86043;
    wire N__86042;
    wire N__86041;
    wire N__86040;
    wire N__86039;
    wire N__86038;
    wire N__86037;
    wire N__86036;
    wire N__86035;
    wire N__86034;
    wire N__86033;
    wire N__86032;
    wire N__86031;
    wire N__86030;
    wire N__86029;
    wire N__86028;
    wire N__86027;
    wire N__86026;
    wire N__86025;
    wire N__86024;
    wire N__86023;
    wire N__86022;
    wire N__86021;
    wire N__86020;
    wire N__86019;
    wire N__86018;
    wire N__86017;
    wire N__86016;
    wire N__86015;
    wire N__86014;
    wire N__86013;
    wire N__86012;
    wire N__86011;
    wire N__86010;
    wire N__86009;
    wire N__86008;
    wire N__86007;
    wire N__86006;
    wire N__86005;
    wire N__86004;
    wire N__86003;
    wire N__86002;
    wire N__85999;
    wire N__85996;
    wire N__85993;
    wire N__85990;
    wire N__85987;
    wire N__85984;
    wire N__85981;
    wire N__85978;
    wire N__85975;
    wire N__85972;
    wire N__85969;
    wire N__85966;
    wire N__85963;
    wire N__85960;
    wire N__85957;
    wire N__85954;
    wire N__85951;
    wire N__85830;
    wire N__85827;
    wire N__85824;
    wire N__85821;
    wire N__85818;
    wire N__85815;
    wire N__85812;
    wire N__85811;
    wire N__85810;
    wire N__85809;
    wire N__85806;
    wire N__85799;
    wire N__85798;
    wire N__85795;
    wire N__85792;
    wire N__85789;
    wire N__85782;
    wire N__85779;
    wire N__85776;
    wire N__85773;
    wire N__85772;
    wire N__85767;
    wire N__85766;
    wire N__85763;
    wire N__85760;
    wire N__85755;
    wire N__85754;
    wire N__85753;
    wire N__85752;
    wire N__85751;
    wire N__85748;
    wire N__85747;
    wire N__85746;
    wire N__85745;
    wire N__85742;
    wire N__85741;
    wire N__85738;
    wire N__85735;
    wire N__85732;
    wire N__85729;
    wire N__85728;
    wire N__85725;
    wire N__85724;
    wire N__85723;
    wire N__85720;
    wire N__85717;
    wire N__85714;
    wire N__85711;
    wire N__85710;
    wire N__85709;
    wire N__85708;
    wire N__85705;
    wire N__85702;
    wire N__85699;
    wire N__85696;
    wire N__85693;
    wire N__85690;
    wire N__85687;
    wire N__85684;
    wire N__85681;
    wire N__85676;
    wire N__85673;
    wire N__85670;
    wire N__85667;
    wire N__85664;
    wire N__85657;
    wire N__85652;
    wire N__85647;
    wire N__85644;
    wire N__85631;
    wire N__85620;
    wire N__85617;
    wire N__85614;
    wire N__85611;
    wire N__85610;
    wire N__85609;
    wire N__85608;
    wire N__85605;
    wire N__85602;
    wire N__85597;
    wire N__85594;
    wire N__85593;
    wire N__85592;
    wire N__85587;
    wire N__85586;
    wire N__85585;
    wire N__85582;
    wire N__85577;
    wire N__85574;
    wire N__85571;
    wire N__85568;
    wire N__85557;
    wire N__85556;
    wire N__85553;
    wire N__85552;
    wire N__85549;
    wire N__85548;
    wire N__85543;
    wire N__85538;
    wire N__85537;
    wire N__85534;
    wire N__85531;
    wire N__85530;
    wire N__85529;
    wire N__85526;
    wire N__85521;
    wire N__85518;
    wire N__85515;
    wire N__85506;
    wire N__85505;
    wire N__85504;
    wire N__85503;
    wire N__85500;
    wire N__85495;
    wire N__85492;
    wire N__85491;
    wire N__85490;
    wire N__85489;
    wire N__85486;
    wire N__85483;
    wire N__85480;
    wire N__85475;
    wire N__85472;
    wire N__85469;
    wire N__85466;
    wire N__85463;
    wire N__85458;
    wire N__85455;
    wire N__85448;
    wire N__85443;
    wire N__85440;
    wire N__85437;
    wire N__85434;
    wire N__85431;
    wire N__85428;
    wire N__85425;
    wire N__85422;
    wire N__85421;
    wire N__85420;
    wire N__85413;
    wire N__85410;
    wire N__85407;
    wire N__85404;
    wire N__85401;
    wire N__85400;
    wire N__85397;
    wire N__85396;
    wire N__85393;
    wire N__85390;
    wire N__85387;
    wire N__85384;
    wire N__85381;
    wire N__85380;
    wire N__85379;
    wire N__85378;
    wire N__85375;
    wire N__85374;
    wire N__85371;
    wire N__85368;
    wire N__85365;
    wire N__85364;
    wire N__85363;
    wire N__85362;
    wire N__85361;
    wire N__85358;
    wire N__85357;
    wire N__85356;
    wire N__85353;
    wire N__85350;
    wire N__85347;
    wire N__85340;
    wire N__85337;
    wire N__85334;
    wire N__85331;
    wire N__85328;
    wire N__85325;
    wire N__85322;
    wire N__85321;
    wire N__85318;
    wire N__85315;
    wire N__85312;
    wire N__85309;
    wire N__85308;
    wire N__85305;
    wire N__85302;
    wire N__85295;
    wire N__85292;
    wire N__85289;
    wire N__85288;
    wire N__85285;
    wire N__85280;
    wire N__85277;
    wire N__85274;
    wire N__85271;
    wire N__85268;
    wire N__85259;
    wire N__85254;
    wire N__85251;
    wire N__85236;
    wire N__85233;
    wire N__85232;
    wire N__85229;
    wire N__85226;
    wire N__85223;
    wire N__85220;
    wire N__85215;
    wire N__85214;
    wire N__85211;
    wire N__85210;
    wire N__85209;
    wire N__85206;
    wire N__85203;
    wire N__85200;
    wire N__85199;
    wire N__85198;
    wire N__85195;
    wire N__85192;
    wire N__85189;
    wire N__85188;
    wire N__85187;
    wire N__85184;
    wire N__85181;
    wire N__85178;
    wire N__85177;
    wire N__85174;
    wire N__85169;
    wire N__85168;
    wire N__85165;
    wire N__85162;
    wire N__85159;
    wire N__85158;
    wire N__85155;
    wire N__85152;
    wire N__85149;
    wire N__85146;
    wire N__85143;
    wire N__85140;
    wire N__85133;
    wire N__85132;
    wire N__85131;
    wire N__85130;
    wire N__85127;
    wire N__85122;
    wire N__85119;
    wire N__85116;
    wire N__85113;
    wire N__85110;
    wire N__85107;
    wire N__85104;
    wire N__85099;
    wire N__85098;
    wire N__85097;
    wire N__85086;
    wire N__85079;
    wire N__85076;
    wire N__85071;
    wire N__85062;
    wire N__85061;
    wire N__85058;
    wire N__85055;
    wire N__85052;
    wire N__85049;
    wire N__85044;
    wire N__85041;
    wire N__85040;
    wire N__85039;
    wire N__85036;
    wire N__85033;
    wire N__85030;
    wire N__85029;
    wire N__85028;
    wire N__85027;
    wire N__85026;
    wire N__85023;
    wire N__85020;
    wire N__85019;
    wire N__85016;
    wire N__85013;
    wire N__85010;
    wire N__85009;
    wire N__85006;
    wire N__85003;
    wire N__85000;
    wire N__84997;
    wire N__84994;
    wire N__84991;
    wire N__84988;
    wire N__84987;
    wire N__84984;
    wire N__84983;
    wire N__84980;
    wire N__84979;
    wire N__84974;
    wire N__84971;
    wire N__84968;
    wire N__84961;
    wire N__84960;
    wire N__84957;
    wire N__84954;
    wire N__84951;
    wire N__84948;
    wire N__84945;
    wire N__84940;
    wire N__84937;
    wire N__84936;
    wire N__84933;
    wire N__84930;
    wire N__84927;
    wire N__84924;
    wire N__84913;
    wire N__84910;
    wire N__84907;
    wire N__84894;
    wire N__84893;
    wire N__84890;
    wire N__84887;
    wire N__84884;
    wire N__84881;
    wire N__84876;
    wire N__84873;
    wire N__84870;
    wire N__84869;
    wire N__84868;
    wire N__84867;
    wire N__84866;
    wire N__84863;
    wire N__84860;
    wire N__84857;
    wire N__84854;
    wire N__84851;
    wire N__84846;
    wire N__84839;
    wire N__84834;
    wire N__84831;
    wire N__84830;
    wire N__84827;
    wire N__84824;
    wire N__84819;
    wire N__84816;
    wire N__84813;
    wire N__84810;
    wire N__84807;
    wire N__84806;
    wire N__84805;
    wire N__84804;
    wire N__84801;
    wire N__84800;
    wire N__84799;
    wire N__84798;
    wire N__84793;
    wire N__84788;
    wire N__84785;
    wire N__84780;
    wire N__84775;
    wire N__84772;
    wire N__84769;
    wire N__84766;
    wire N__84763;
    wire N__84760;
    wire N__84757;
    wire N__84750;
    wire N__84747;
    wire N__84744;
    wire N__84741;
    wire N__84738;
    wire N__84737;
    wire N__84736;
    wire N__84729;
    wire N__84726;
    wire N__84723;
    wire N__84720;
    wire N__84717;
    wire N__84716;
    wire N__84715;
    wire N__84708;
    wire N__84705;
    wire N__84702;
    wire N__84699;
    wire N__84696;
    wire N__84693;
    wire N__84692;
    wire N__84691;
    wire N__84684;
    wire N__84681;
    wire N__84678;
    wire N__84675;
    wire N__84672;
    wire N__84669;
    wire N__84666;
    wire N__84665;
    wire N__84664;
    wire N__84657;
    wire N__84654;
    wire N__84651;
    wire N__84648;
    wire N__84645;
    wire N__84642;
    wire N__84639;
    wire N__84636;
    wire N__84633;
    wire N__84632;
    wire N__84631;
    wire N__84630;
    wire N__84629;
    wire N__84626;
    wire N__84625;
    wire N__84624;
    wire N__84623;
    wire N__84622;
    wire N__84621;
    wire N__84614;
    wire N__84605;
    wire N__84598;
    wire N__84595;
    wire N__84594;
    wire N__84593;
    wire N__84592;
    wire N__84591;
    wire N__84588;
    wire N__84585;
    wire N__84582;
    wire N__84573;
    wire N__84570;
    wire N__84567;
    wire N__84564;
    wire N__84561;
    wire N__84558;
    wire N__84555;
    wire N__84546;
    wire N__84543;
    wire N__84540;
    wire N__84537;
    wire N__84536;
    wire N__84535;
    wire N__84530;
    wire N__84527;
    wire N__84524;
    wire N__84519;
    wire N__84516;
    wire N__84513;
    wire N__84510;
    wire N__84507;
    wire N__84504;
    wire N__84501;
    wire N__84500;
    wire N__84497;
    wire N__84494;
    wire N__84489;
    wire N__84486;
    wire N__84483;
    wire N__84480;
    wire N__84477;
    wire N__84474;
    wire N__84471;
    wire N__84468;
    wire N__84465;
    wire N__84462;
    wire N__84459;
    wire N__84458;
    wire N__84457;
    wire N__84456;
    wire N__84453;
    wire N__84450;
    wire N__84445;
    wire N__84442;
    wire N__84439;
    wire N__84436;
    wire N__84431;
    wire N__84428;
    wire N__84423;
    wire N__84420;
    wire N__84417;
    wire N__84416;
    wire N__84413;
    wire N__84410;
    wire N__84405;
    wire N__84402;
    wire N__84399;
    wire N__84396;
    wire N__84393;
    wire N__84390;
    wire N__84387;
    wire N__84384;
    wire N__84383;
    wire N__84378;
    wire N__84375;
    wire N__84372;
    wire N__84369;
    wire N__84366;
    wire N__84363;
    wire N__84360;
    wire N__84357;
    wire N__84354;
    wire N__84351;
    wire N__84350;
    wire N__84345;
    wire N__84342;
    wire N__84339;
    wire N__84336;
    wire N__84333;
    wire N__84330;
    wire N__84329;
    wire N__84324;
    wire N__84321;
    wire N__84318;
    wire N__84315;
    wire N__84312;
    wire N__84309;
    wire N__84308;
    wire N__84305;
    wire N__84302;
    wire N__84297;
    wire N__84294;
    wire N__84291;
    wire N__84288;
    wire N__84285;
    wire N__84284;
    wire N__84281;
    wire N__84278;
    wire N__84275;
    wire N__84272;
    wire N__84267;
    wire N__84264;
    wire N__84261;
    wire N__84260;
    wire N__84257;
    wire N__84254;
    wire N__84253;
    wire N__84252;
    wire N__84247;
    wire N__84242;
    wire N__84239;
    wire N__84234;
    wire N__84231;
    wire N__84228;
    wire N__84225;
    wire N__84222;
    wire N__84221;
    wire N__84216;
    wire N__84215;
    wire N__84214;
    wire N__84211;
    wire N__84210;
    wire N__84209;
    wire N__84208;
    wire N__84205;
    wire N__84204;
    wire N__84201;
    wire N__84198;
    wire N__84195;
    wire N__84192;
    wire N__84189;
    wire N__84186;
    wire N__84183;
    wire N__84182;
    wire N__84179;
    wire N__84174;
    wire N__84171;
    wire N__84168;
    wire N__84165;
    wire N__84162;
    wire N__84161;
    wire N__84160;
    wire N__84157;
    wire N__84156;
    wire N__84151;
    wire N__84148;
    wire N__84147;
    wire N__84144;
    wire N__84139;
    wire N__84136;
    wire N__84133;
    wire N__84132;
    wire N__84131;
    wire N__84128;
    wire N__84125;
    wire N__84124;
    wire N__84123;
    wire N__84120;
    wire N__84117;
    wire N__84114;
    wire N__84109;
    wire N__84106;
    wire N__84103;
    wire N__84098;
    wire N__84093;
    wire N__84090;
    wire N__84087;
    wire N__84078;
    wire N__84073;
    wire N__84070;
    wire N__84065;
    wire N__84054;
    wire N__84053;
    wire N__84050;
    wire N__84047;
    wire N__84044;
    wire N__84041;
    wire N__84038;
    wire N__84035;
    wire N__84030;
    wire N__84029;
    wire N__84028;
    wire N__84025;
    wire N__84022;
    wire N__84021;
    wire N__84020;
    wire N__84019;
    wire N__84016;
    wire N__84013;
    wire N__84010;
    wire N__84003;
    wire N__84002;
    wire N__84001;
    wire N__84000;
    wire N__83997;
    wire N__83994;
    wire N__83989;
    wire N__83988;
    wire N__83985;
    wire N__83984;
    wire N__83981;
    wire N__83980;
    wire N__83977;
    wire N__83974;
    wire N__83969;
    wire N__83968;
    wire N__83965;
    wire N__83962;
    wire N__83959;
    wire N__83956;
    wire N__83953;
    wire N__83948;
    wire N__83947;
    wire N__83946;
    wire N__83945;
    wire N__83942;
    wire N__83939;
    wire N__83938;
    wire N__83935;
    wire N__83932;
    wire N__83929;
    wire N__83926;
    wire N__83923;
    wire N__83920;
    wire N__83915;
    wire N__83912;
    wire N__83907;
    wire N__83904;
    wire N__83893;
    wire N__83888;
    wire N__83885;
    wire N__83874;
    wire N__83871;
    wire N__83870;
    wire N__83867;
    wire N__83864;
    wire N__83861;
    wire N__83858;
    wire N__83853;
    wire N__83850;
    wire N__83849;
    wire N__83848;
    wire N__83841;
    wire N__83838;
    wire N__83837;
    wire N__83836;
    wire N__83835;
    wire N__83832;
    wire N__83829;
    wire N__83828;
    wire N__83825;
    wire N__83822;
    wire N__83817;
    wire N__83814;
    wire N__83811;
    wire N__83808;
    wire N__83807;
    wire N__83804;
    wire N__83801;
    wire N__83798;
    wire N__83797;
    wire N__83796;
    wire N__83795;
    wire N__83794;
    wire N__83791;
    wire N__83788;
    wire N__83787;
    wire N__83782;
    wire N__83779;
    wire N__83776;
    wire N__83773;
    wire N__83770;
    wire N__83769;
    wire N__83766;
    wire N__83761;
    wire N__83758;
    wire N__83757;
    wire N__83756;
    wire N__83755;
    wire N__83750;
    wire N__83747;
    wire N__83744;
    wire N__83741;
    wire N__83738;
    wire N__83735;
    wire N__83732;
    wire N__83729;
    wire N__83724;
    wire N__83723;
    wire N__83720;
    wire N__83717;
    wire N__83714;
    wire N__83707;
    wire N__83698;
    wire N__83695;
    wire N__83682;
    wire N__83681;
    wire N__83678;
    wire N__83675;
    wire N__83672;
    wire N__83669;
    wire N__83666;
    wire N__83663;
    wire N__83658;
    wire N__83655;
    wire N__83652;
    wire N__83649;
    wire N__83646;
    wire N__83643;
    wire N__83642;
    wire N__83641;
    wire N__83636;
    wire N__83633;
    wire N__83630;
    wire N__83627;
    wire N__83624;
    wire N__83621;
    wire N__83618;
    wire N__83615;
    wire N__83612;
    wire N__83607;
    wire N__83604;
    wire N__83601;
    wire N__83598;
    wire N__83597;
    wire N__83592;
    wire N__83589;
    wire N__83586;
    wire N__83583;
    wire N__83580;
    wire N__83577;
    wire N__83574;
    wire N__83573;
    wire N__83570;
    wire N__83569;
    wire N__83568;
    wire N__83567;
    wire N__83566;
    wire N__83563;
    wire N__83562;
    wire N__83553;
    wire N__83552;
    wire N__83551;
    wire N__83550;
    wire N__83549;
    wire N__83548;
    wire N__83541;
    wire N__83538;
    wire N__83537;
    wire N__83534;
    wire N__83533;
    wire N__83532;
    wire N__83523;
    wire N__83520;
    wire N__83517;
    wire N__83508;
    wire N__83505;
    wire N__83502;
    wire N__83499;
    wire N__83496;
    wire N__83493;
    wire N__83490;
    wire N__83485;
    wire N__83480;
    wire N__83475;
    wire N__83472;
    wire N__83469;
    wire N__83466;
    wire N__83465;
    wire N__83460;
    wire N__83457;
    wire N__83454;
    wire N__83451;
    wire N__83450;
    wire N__83445;
    wire N__83442;
    wire N__83441;
    wire N__83436;
    wire N__83433;
    wire N__83430;
    wire N__83427;
    wire N__83424;
    wire N__83423;
    wire N__83418;
    wire N__83415;
    wire N__83412;
    wire N__83409;
    wire N__83406;
    wire N__83405;
    wire N__83404;
    wire N__83403;
    wire N__83402;
    wire N__83401;
    wire N__83400;
    wire N__83399;
    wire N__83398;
    wire N__83397;
    wire N__83394;
    wire N__83393;
    wire N__83392;
    wire N__83389;
    wire N__83386;
    wire N__83385;
    wire N__83382;
    wire N__83379;
    wire N__83376;
    wire N__83373;
    wire N__83370;
    wire N__83367;
    wire N__83364;
    wire N__83361;
    wire N__83358;
    wire N__83355;
    wire N__83350;
    wire N__83347;
    wire N__83342;
    wire N__83339;
    wire N__83336;
    wire N__83333;
    wire N__83330;
    wire N__83329;
    wire N__83326;
    wire N__83321;
    wire N__83316;
    wire N__83313;
    wire N__83308;
    wire N__83303;
    wire N__83300;
    wire N__83297;
    wire N__83290;
    wire N__83285;
    wire N__83282;
    wire N__83279;
    wire N__83274;
    wire N__83271;
    wire N__83262;
    wire N__83261;
    wire N__83258;
    wire N__83257;
    wire N__83256;
    wire N__83255;
    wire N__83254;
    wire N__83251;
    wire N__83248;
    wire N__83245;
    wire N__83244;
    wire N__83241;
    wire N__83240;
    wire N__83237;
    wire N__83236;
    wire N__83233;
    wire N__83230;
    wire N__83229;
    wire N__83228;
    wire N__83223;
    wire N__83220;
    wire N__83219;
    wire N__83218;
    wire N__83215;
    wire N__83212;
    wire N__83209;
    wire N__83206;
    wire N__83201;
    wire N__83198;
    wire N__83195;
    wire N__83190;
    wire N__83187;
    wire N__83184;
    wire N__83183;
    wire N__83178;
    wire N__83177;
    wire N__83174;
    wire N__83171;
    wire N__83166;
    wire N__83159;
    wire N__83156;
    wire N__83153;
    wire N__83150;
    wire N__83147;
    wire N__83142;
    wire N__83139;
    wire N__83136;
    wire N__83131;
    wire N__83128;
    wire N__83125;
    wire N__83120;
    wire N__83115;
    wire N__83110;
    wire N__83103;
    wire N__83102;
    wire N__83097;
    wire N__83094;
    wire N__83093;
    wire N__83090;
    wire N__83087;
    wire N__83084;
    wire N__83081;
    wire N__83078;
    wire N__83075;
    wire N__83072;
    wire N__83069;
    wire N__83064;
    wire N__83061;
    wire N__83058;
    wire N__83055;
    wire N__83052;
    wire N__83049;
    wire N__83046;
    wire N__83045;
    wire N__83044;
    wire N__83043;
    wire N__83042;
    wire N__83041;
    wire N__83038;
    wire N__83029;
    wire N__83026;
    wire N__83021;
    wire N__83016;
    wire N__83013;
    wire N__83012;
    wire N__83011;
    wire N__83008;
    wire N__83003;
    wire N__83002;
    wire N__82999;
    wire N__82996;
    wire N__82993;
    wire N__82986;
    wire N__82983;
    wire N__82980;
    wire N__82977;
    wire N__82976;
    wire N__82973;
    wire N__82970;
    wire N__82965;
    wire N__82962;
    wire N__82961;
    wire N__82958;
    wire N__82955;
    wire N__82952;
    wire N__82949;
    wire N__82946;
    wire N__82943;
    wire N__82938;
    wire N__82937;
    wire N__82934;
    wire N__82931;
    wire N__82928;
    wire N__82923;
    wire N__82920;
    wire N__82919;
    wire N__82914;
    wire N__82911;
    wire N__82908;
    wire N__82905;
    wire N__82902;
    wire N__82899;
    wire N__82896;
    wire N__82893;
    wire N__82892;
    wire N__82891;
    wire N__82890;
    wire N__82889;
    wire N__82882;
    wire N__82877;
    wire N__82872;
    wire N__82869;
    wire N__82868;
    wire N__82865;
    wire N__82862;
    wire N__82857;
    wire N__82854;
    wire N__82851;
    wire N__82850;
    wire N__82847;
    wire N__82844;
    wire N__82843;
    wire N__82842;
    wire N__82841;
    wire N__82838;
    wire N__82835;
    wire N__82834;
    wire N__82833;
    wire N__82832;
    wire N__82831;
    wire N__82828;
    wire N__82827;
    wire N__82822;
    wire N__82819;
    wire N__82816;
    wire N__82811;
    wire N__82802;
    wire N__82799;
    wire N__82788;
    wire N__82785;
    wire N__82782;
    wire N__82779;
    wire N__82776;
    wire N__82775;
    wire N__82772;
    wire N__82771;
    wire N__82770;
    wire N__82769;
    wire N__82766;
    wire N__82763;
    wire N__82760;
    wire N__82757;
    wire N__82754;
    wire N__82747;
    wire N__82744;
    wire N__82741;
    wire N__82738;
    wire N__82733;
    wire N__82730;
    wire N__82727;
    wire N__82724;
    wire N__82721;
    wire N__82716;
    wire N__82713;
    wire N__82712;
    wire N__82709;
    wire N__82706;
    wire N__82703;
    wire N__82700;
    wire N__82697;
    wire N__82692;
    wire N__82689;
    wire N__82688;
    wire N__82685;
    wire N__82682;
    wire N__82679;
    wire N__82676;
    wire N__82675;
    wire N__82672;
    wire N__82669;
    wire N__82666;
    wire N__82659;
    wire N__82656;
    wire N__82653;
    wire N__82650;
    wire N__82649;
    wire N__82646;
    wire N__82643;
    wire N__82640;
    wire N__82637;
    wire N__82632;
    wire N__82629;
    wire N__82626;
    wire N__82625;
    wire N__82622;
    wire N__82619;
    wire N__82614;
    wire N__82611;
    wire N__82608;
    wire N__82607;
    wire N__82604;
    wire N__82601;
    wire N__82596;
    wire N__82593;
    wire N__82590;
    wire N__82587;
    wire N__82584;
    wire N__82583;
    wire N__82580;
    wire N__82577;
    wire N__82574;
    wire N__82571;
    wire N__82566;
    wire N__82565;
    wire N__82564;
    wire N__82563;
    wire N__82560;
    wire N__82553;
    wire N__82548;
    wire N__82545;
    wire N__82542;
    wire N__82539;
    wire N__82536;
    wire N__82535;
    wire N__82534;
    wire N__82527;
    wire N__82524;
    wire N__82521;
    wire N__82518;
    wire N__82515;
    wire N__82512;
    wire N__82511;
    wire N__82508;
    wire N__82505;
    wire N__82504;
    wire N__82503;
    wire N__82500;
    wire N__82493;
    wire N__82488;
    wire N__82485;
    wire N__82482;
    wire N__82481;
    wire N__82480;
    wire N__82477;
    wire N__82474;
    wire N__82469;
    wire N__82464;
    wire N__82461;
    wire N__82458;
    wire N__82455;
    wire N__82452;
    wire N__82449;
    wire N__82446;
    wire N__82445;
    wire N__82442;
    wire N__82439;
    wire N__82438;
    wire N__82435;
    wire N__82432;
    wire N__82429;
    wire N__82422;
    wire N__82421;
    wire N__82418;
    wire N__82415;
    wire N__82410;
    wire N__82407;
    wire N__82406;
    wire N__82403;
    wire N__82400;
    wire N__82397;
    wire N__82394;
    wire N__82391;
    wire N__82388;
    wire N__82385;
    wire N__82382;
    wire N__82377;
    wire N__82376;
    wire N__82371;
    wire N__82368;
    wire N__82365;
    wire N__82362;
    wire N__82359;
    wire N__82356;
    wire N__82353;
    wire N__82350;
    wire N__82347;
    wire N__82344;
    wire N__82341;
    wire N__82340;
    wire N__82339;
    wire N__82336;
    wire N__82333;
    wire N__82332;
    wire N__82329;
    wire N__82328;
    wire N__82321;
    wire N__82316;
    wire N__82311;
    wire N__82308;
    wire N__82305;
    wire N__82302;
    wire N__82299;
    wire N__82298;
    wire N__82297;
    wire N__82290;
    wire N__82287;
    wire N__82284;
    wire N__82281;
    wire N__82278;
    wire N__82277;
    wire N__82274;
    wire N__82273;
    wire N__82272;
    wire N__82271;
    wire N__82270;
    wire N__82269;
    wire N__82266;
    wire N__82261;
    wire N__82258;
    wire N__82257;
    wire N__82254;
    wire N__82251;
    wire N__82248;
    wire N__82243;
    wire N__82238;
    wire N__82227;
    wire N__82226;
    wire N__82223;
    wire N__82220;
    wire N__82215;
    wire N__82212;
    wire N__82209;
    wire N__82206;
    wire N__82203;
    wire N__82200;
    wire N__82199;
    wire N__82196;
    wire N__82193;
    wire N__82190;
    wire N__82187;
    wire N__82182;
    wire N__82179;
    wire N__82176;
    wire N__82173;
    wire N__82170;
    wire N__82167;
    wire N__82166;
    wire N__82163;
    wire N__82162;
    wire N__82159;
    wire N__82156;
    wire N__82153;
    wire N__82150;
    wire N__82147;
    wire N__82144;
    wire N__82141;
    wire N__82134;
    wire N__82131;
    wire N__82128;
    wire N__82125;
    wire N__82122;
    wire N__82119;
    wire N__82116;
    wire N__82113;
    wire N__82110;
    wire N__82109;
    wire N__82106;
    wire N__82103;
    wire N__82102;
    wire N__82099;
    wire N__82096;
    wire N__82093;
    wire N__82092;
    wire N__82087;
    wire N__82082;
    wire N__82077;
    wire N__82076;
    wire N__82075;
    wire N__82074;
    wire N__82071;
    wire N__82066;
    wire N__82063;
    wire N__82056;
    wire N__82053;
    wire N__82052;
    wire N__82051;
    wire N__82048;
    wire N__82045;
    wire N__82042;
    wire N__82035;
    wire N__82032;
    wire N__82029;
    wire N__82026;
    wire N__82023;
    wire N__82022;
    wire N__82021;
    wire N__82018;
    wire N__82015;
    wire N__82012;
    wire N__82009;
    wire N__82006;
    wire N__82003;
    wire N__82000;
    wire N__81997;
    wire N__81994;
    wire N__81989;
    wire N__81984;
    wire N__81983;
    wire N__81982;
    wire N__81979;
    wire N__81976;
    wire N__81975;
    wire N__81972;
    wire N__81969;
    wire N__81966;
    wire N__81963;
    wire N__81960;
    wire N__81957;
    wire N__81952;
    wire N__81949;
    wire N__81944;
    wire N__81939;
    wire N__81936;
    wire N__81933;
    wire N__81930;
    wire N__81927;
    wire N__81926;
    wire N__81923;
    wire N__81920;
    wire N__81915;
    wire N__81912;
    wire N__81909;
    wire N__81906;
    wire N__81903;
    wire N__81902;
    wire N__81901;
    wire N__81900;
    wire N__81897;
    wire N__81894;
    wire N__81889;
    wire N__81882;
    wire N__81879;
    wire N__81876;
    wire N__81873;
    wire N__81870;
    wire N__81869;
    wire N__81866;
    wire N__81865;
    wire N__81864;
    wire N__81861;
    wire N__81858;
    wire N__81853;
    wire N__81846;
    wire N__81843;
    wire N__81842;
    wire N__81837;
    wire N__81834;
    wire N__81831;
    wire N__81830;
    wire N__81829;
    wire N__81828;
    wire N__81827;
    wire N__81820;
    wire N__81815;
    wire N__81810;
    wire N__81807;
    wire N__81804;
    wire N__81801;
    wire N__81798;
    wire N__81795;
    wire N__81792;
    wire N__81789;
    wire N__81786;
    wire N__81783;
    wire N__81780;
    wire N__81777;
    wire N__81776;
    wire N__81775;
    wire N__81770;
    wire N__81767;
    wire N__81764;
    wire N__81761;
    wire N__81758;
    wire N__81753;
    wire N__81750;
    wire N__81747;
    wire N__81744;
    wire N__81741;
    wire N__81738;
    wire N__81735;
    wire N__81734;
    wire N__81731;
    wire N__81728;
    wire N__81725;
    wire N__81722;
    wire N__81719;
    wire N__81716;
    wire N__81711;
    wire N__81710;
    wire N__81705;
    wire N__81702;
    wire N__81699;
    wire N__81698;
    wire N__81695;
    wire N__81692;
    wire N__81687;
    wire N__81684;
    wire N__81681;
    wire N__81678;
    wire N__81675;
    wire N__81672;
    wire N__81671;
    wire N__81666;
    wire N__81663;
    wire N__81660;
    wire N__81657;
    wire N__81654;
    wire N__81653;
    wire N__81650;
    wire N__81647;
    wire N__81642;
    wire N__81639;
    wire N__81636;
    wire N__81633;
    wire N__81630;
    wire N__81627;
    wire N__81626;
    wire N__81623;
    wire N__81620;
    wire N__81619;
    wire N__81616;
    wire N__81611;
    wire N__81606;
    wire N__81605;
    wire N__81602;
    wire N__81599;
    wire N__81596;
    wire N__81593;
    wire N__81588;
    wire N__81585;
    wire N__81582;
    wire N__81579;
    wire N__81576;
    wire N__81573;
    wire N__81570;
    wire N__81567;
    wire N__81564;
    wire N__81563;
    wire N__81560;
    wire N__81557;
    wire N__81552;
    wire N__81549;
    wire N__81548;
    wire N__81545;
    wire N__81542;
    wire N__81537;
    wire N__81534;
    wire N__81531;
    wire N__81528;
    wire N__81525;
    wire N__81524;
    wire N__81521;
    wire N__81520;
    wire N__81517;
    wire N__81514;
    wire N__81511;
    wire N__81508;
    wire N__81501;
    wire N__81498;
    wire N__81495;
    wire N__81492;
    wire N__81489;
    wire N__81486;
    wire N__81483;
    wire N__81482;
    wire N__81481;
    wire N__81478;
    wire N__81473;
    wire N__81470;
    wire N__81467;
    wire N__81462;
    wire N__81459;
    wire N__81456;
    wire N__81453;
    wire N__81450;
    wire N__81447;
    wire N__81444;
    wire N__81441;
    wire N__81440;
    wire N__81437;
    wire N__81434;
    wire N__81431;
    wire N__81426;
    wire N__81423;
    wire N__81422;
    wire N__81417;
    wire N__81414;
    wire N__81413;
    wire N__81408;
    wire N__81405;
    wire N__81402;
    wire N__81399;
    wire N__81396;
    wire N__81393;
    wire N__81390;
    wire N__81387;
    wire N__81384;
    wire N__81381;
    wire N__81380;
    wire N__81377;
    wire N__81374;
    wire N__81371;
    wire N__81368;
    wire N__81367;
    wire N__81366;
    wire N__81365;
    wire N__81362;
    wire N__81359;
    wire N__81352;
    wire N__81345;
    wire N__81342;
    wire N__81339;
    wire N__81336;
    wire N__81333;
    wire N__81330;
    wire N__81327;
    wire N__81324;
    wire N__81321;
    wire N__81318;
    wire N__81315;
    wire N__81312;
    wire N__81309;
    wire N__81308;
    wire N__81303;
    wire N__81302;
    wire N__81301;
    wire N__81300;
    wire N__81299;
    wire N__81296;
    wire N__81287;
    wire N__81282;
    wire N__81279;
    wire N__81276;
    wire N__81273;
    wire N__81270;
    wire N__81269;
    wire N__81268;
    wire N__81267;
    wire N__81258;
    wire N__81255;
    wire N__81252;
    wire N__81249;
    wire N__81246;
    wire N__81243;
    wire N__81240;
    wire N__81237;
    wire N__81234;
    wire N__81233;
    wire N__81230;
    wire N__81229;
    wire N__81228;
    wire N__81225;
    wire N__81222;
    wire N__81217;
    wire N__81214;
    wire N__81211;
    wire N__81208;
    wire N__81205;
    wire N__81202;
    wire N__81199;
    wire N__81196;
    wire N__81193;
    wire N__81188;
    wire N__81183;
    wire N__81180;
    wire N__81177;
    wire N__81174;
    wire N__81171;
    wire N__81170;
    wire N__81169;
    wire N__81166;
    wire N__81163;
    wire N__81162;
    wire N__81153;
    wire N__81150;
    wire N__81147;
    wire N__81144;
    wire N__81141;
    wire N__81138;
    wire N__81135;
    wire N__81132;
    wire N__81129;
    wire N__81128;
    wire N__81127;
    wire N__81120;
    wire N__81119;
    wire N__81118;
    wire N__81115;
    wire N__81110;
    wire N__81105;
    wire N__81102;
    wire N__81099;
    wire N__81096;
    wire N__81093;
    wire N__81090;
    wire N__81087;
    wire N__81084;
    wire N__81081;
    wire N__81078;
    wire N__81075;
    wire N__81072;
    wire N__81071;
    wire N__81068;
    wire N__81067;
    wire N__81064;
    wire N__81061;
    wire N__81060;
    wire N__81059;
    wire N__81058;
    wire N__81057;
    wire N__81054;
    wire N__81051;
    wire N__81048;
    wire N__81047;
    wire N__81044;
    wire N__81041;
    wire N__81038;
    wire N__81035;
    wire N__81032;
    wire N__81027;
    wire N__81024;
    wire N__81021;
    wire N__81018;
    wire N__81015;
    wire N__81012;
    wire N__81009;
    wire N__81004;
    wire N__81001;
    wire N__80998;
    wire N__80989;
    wire N__80982;
    wire N__80981;
    wire N__80980;
    wire N__80977;
    wire N__80976;
    wire N__80975;
    wire N__80974;
    wire N__80973;
    wire N__80972;
    wire N__80971;
    wire N__80968;
    wire N__80965;
    wire N__80964;
    wire N__80963;
    wire N__80962;
    wire N__80961;
    wire N__80960;
    wire N__80959;
    wire N__80956;
    wire N__80953;
    wire N__80948;
    wire N__80945;
    wire N__80944;
    wire N__80943;
    wire N__80940;
    wire N__80939;
    wire N__80938;
    wire N__80935;
    wire N__80932;
    wire N__80931;
    wire N__80924;
    wire N__80919;
    wire N__80914;
    wire N__80907;
    wire N__80904;
    wire N__80899;
    wire N__80896;
    wire N__80893;
    wire N__80888;
    wire N__80885;
    wire N__80882;
    wire N__80879;
    wire N__80876;
    wire N__80871;
    wire N__80868;
    wire N__80865;
    wire N__80858;
    wire N__80857;
    wire N__80854;
    wire N__80851;
    wire N__80846;
    wire N__80843;
    wire N__80840;
    wire N__80835;
    wire N__80832;
    wire N__80829;
    wire N__80826;
    wire N__80823;
    wire N__80820;
    wire N__80817;
    wire N__80814;
    wire N__80809;
    wire N__80796;
    wire N__80795;
    wire N__80794;
    wire N__80793;
    wire N__80792;
    wire N__80791;
    wire N__80788;
    wire N__80787;
    wire N__80786;
    wire N__80781;
    wire N__80780;
    wire N__80779;
    wire N__80778;
    wire N__80775;
    wire N__80774;
    wire N__80771;
    wire N__80768;
    wire N__80767;
    wire N__80766;
    wire N__80765;
    wire N__80764;
    wire N__80759;
    wire N__80756;
    wire N__80755;
    wire N__80754;
    wire N__80751;
    wire N__80748;
    wire N__80745;
    wire N__80742;
    wire N__80739;
    wire N__80738;
    wire N__80735;
    wire N__80732;
    wire N__80729;
    wire N__80726;
    wire N__80725;
    wire N__80722;
    wire N__80721;
    wire N__80718;
    wire N__80715;
    wire N__80710;
    wire N__80705;
    wire N__80704;
    wire N__80703;
    wire N__80702;
    wire N__80699;
    wire N__80694;
    wire N__80689;
    wire N__80686;
    wire N__80683;
    wire N__80680;
    wire N__80675;
    wire N__80670;
    wire N__80667;
    wire N__80664;
    wire N__80659;
    wire N__80656;
    wire N__80649;
    wire N__80646;
    wire N__80639;
    wire N__80616;
    wire N__80615;
    wire N__80614;
    wire N__80613;
    wire N__80612;
    wire N__80611;
    wire N__80610;
    wire N__80609;
    wire N__80608;
    wire N__80607;
    wire N__80604;
    wire N__80603;
    wire N__80600;
    wire N__80599;
    wire N__80596;
    wire N__80595;
    wire N__80594;
    wire N__80591;
    wire N__80586;
    wire N__80583;
    wire N__80580;
    wire N__80577;
    wire N__80572;
    wire N__80569;
    wire N__80568;
    wire N__80567;
    wire N__80564;
    wire N__80561;
    wire N__80558;
    wire N__80555;
    wire N__80554;
    wire N__80551;
    wire N__80542;
    wire N__80539;
    wire N__80538;
    wire N__80537;
    wire N__80536;
    wire N__80535;
    wire N__80534;
    wire N__80533;
    wire N__80532;
    wire N__80529;
    wire N__80526;
    wire N__80523;
    wire N__80522;
    wire N__80521;
    wire N__80520;
    wire N__80519;
    wire N__80516;
    wire N__80515;
    wire N__80512;
    wire N__80507;
    wire N__80502;
    wire N__80497;
    wire N__80494;
    wire N__80491;
    wire N__80484;
    wire N__80479;
    wire N__80476;
    wire N__80475;
    wire N__80472;
    wire N__80467;
    wire N__80460;
    wire N__80453;
    wire N__80450;
    wire N__80441;
    wire N__80436;
    wire N__80431;
    wire N__80428;
    wire N__80423;
    wire N__80418;
    wire N__80413;
    wire N__80408;
    wire N__80397;
    wire N__80396;
    wire N__80395;
    wire N__80394;
    wire N__80391;
    wire N__80390;
    wire N__80387;
    wire N__80384;
    wire N__80383;
    wire N__80382;
    wire N__80379;
    wire N__80378;
    wire N__80377;
    wire N__80372;
    wire N__80369;
    wire N__80366;
    wire N__80365;
    wire N__80364;
    wire N__80363;
    wire N__80360;
    wire N__80357;
    wire N__80354;
    wire N__80351;
    wire N__80348;
    wire N__80347;
    wire N__80344;
    wire N__80341;
    wire N__80340;
    wire N__80339;
    wire N__80338;
    wire N__80335;
    wire N__80330;
    wire N__80327;
    wire N__80324;
    wire N__80321;
    wire N__80318;
    wire N__80313;
    wire N__80310;
    wire N__80305;
    wire N__80304;
    wire N__80301;
    wire N__80298;
    wire N__80295;
    wire N__80288;
    wire N__80287;
    wire N__80284;
    wire N__80281;
    wire N__80278;
    wire N__80275;
    wire N__80270;
    wire N__80267;
    wire N__80264;
    wire N__80261;
    wire N__80256;
    wire N__80253;
    wire N__80250;
    wire N__80239;
    wire N__80230;
    wire N__80223;
    wire N__80222;
    wire N__80217;
    wire N__80214;
    wire N__80213;
    wire N__80210;
    wire N__80207;
    wire N__80202;
    wire N__80201;
    wire N__80198;
    wire N__80195;
    wire N__80190;
    wire N__80187;
    wire N__80184;
    wire N__80181;
    wire N__80178;
    wire N__80175;
    wire N__80172;
    wire N__80169;
    wire N__80166;
    wire N__80163;
    wire N__80160;
    wire N__80157;
    wire N__80156;
    wire N__80151;
    wire N__80148;
    wire N__80145;
    wire N__80142;
    wire N__80139;
    wire N__80136;
    wire N__80133;
    wire N__80130;
    wire N__80127;
    wire N__80126;
    wire N__80123;
    wire N__80118;
    wire N__80115;
    wire N__80112;
    wire N__80111;
    wire N__80108;
    wire N__80105;
    wire N__80104;
    wire N__80101;
    wire N__80096;
    wire N__80091;
    wire N__80088;
    wire N__80085;
    wire N__80082;
    wire N__80079;
    wire N__80076;
    wire N__80073;
    wire N__80070;
    wire N__80067;
    wire N__80064;
    wire N__80061;
    wire N__80058;
    wire N__80057;
    wire N__80056;
    wire N__80053;
    wire N__80048;
    wire N__80043;
    wire N__80040;
    wire N__80037;
    wire N__80034;
    wire N__80031;
    wire N__80028;
    wire N__80025;
    wire N__80022;
    wire N__80019;
    wire N__80016;
    wire N__80015;
    wire N__80012;
    wire N__80009;
    wire N__80006;
    wire N__80001;
    wire N__80000;
    wire N__79999;
    wire N__79998;
    wire N__79997;
    wire N__79996;
    wire N__79995;
    wire N__79994;
    wire N__79993;
    wire N__79992;
    wire N__79991;
    wire N__79990;
    wire N__79987;
    wire N__79986;
    wire N__79985;
    wire N__79984;
    wire N__79983;
    wire N__79982;
    wire N__79981;
    wire N__79980;
    wire N__79979;
    wire N__79978;
    wire N__79977;
    wire N__79976;
    wire N__79975;
    wire N__79974;
    wire N__79973;
    wire N__79970;
    wire N__79969;
    wire N__79968;
    wire N__79967;
    wire N__79966;
    wire N__79965;
    wire N__79964;
    wire N__79963;
    wire N__79962;
    wire N__79961;
    wire N__79960;
    wire N__79959;
    wire N__79958;
    wire N__79957;
    wire N__79956;
    wire N__79955;
    wire N__79954;
    wire N__79953;
    wire N__79952;
    wire N__79951;
    wire N__79950;
    wire N__79949;
    wire N__79948;
    wire N__79947;
    wire N__79946;
    wire N__79945;
    wire N__79944;
    wire N__79943;
    wire N__79942;
    wire N__79941;
    wire N__79938;
    wire N__79937;
    wire N__79936;
    wire N__79935;
    wire N__79934;
    wire N__79933;
    wire N__79932;
    wire N__79931;
    wire N__79930;
    wire N__79929;
    wire N__79928;
    wire N__79927;
    wire N__79926;
    wire N__79925;
    wire N__79924;
    wire N__79923;
    wire N__79922;
    wire N__79921;
    wire N__79920;
    wire N__79919;
    wire N__79918;
    wire N__79917;
    wire N__79916;
    wire N__79915;
    wire N__79912;
    wire N__79909;
    wire N__79904;
    wire N__79901;
    wire N__79896;
    wire N__79893;
    wire N__79888;
    wire N__79885;
    wire N__79882;
    wire N__79879;
    wire N__79876;
    wire N__79871;
    wire N__79864;
    wire N__79857;
    wire N__79850;
    wire N__79845;
    wire N__79842;
    wire N__79839;
    wire N__79836;
    wire N__79831;
    wire N__79826;
    wire N__79823;
    wire N__79820;
    wire N__79813;
    wire N__79810;
    wire N__79805;
    wire N__79800;
    wire N__79793;
    wire N__79784;
    wire N__79779;
    wire N__79776;
    wire N__79771;
    wire N__79768;
    wire N__79765;
    wire N__79762;
    wire N__79759;
    wire N__79752;
    wire N__79747;
    wire N__79740;
    wire N__79737;
    wire N__79732;
    wire N__79725;
    wire N__79722;
    wire N__79719;
    wire N__79716;
    wire N__79713;
    wire N__79712;
    wire N__79711;
    wire N__79710;
    wire N__79709;
    wire N__79708;
    wire N__79707;
    wire N__79706;
    wire N__79705;
    wire N__79704;
    wire N__79703;
    wire N__79702;
    wire N__79701;
    wire N__79700;
    wire N__79699;
    wire N__79698;
    wire N__79697;
    wire N__79696;
    wire N__79695;
    wire N__79694;
    wire N__79693;
    wire N__79692;
    wire N__79691;
    wire N__79690;
    wire N__79689;
    wire N__79688;
    wire N__79687;
    wire N__79686;
    wire N__79685;
    wire N__79684;
    wire N__79683;
    wire N__79682;
    wire N__79681;
    wire N__79680;
    wire N__79679;
    wire N__79678;
    wire N__79677;
    wire N__79676;
    wire N__79675;
    wire N__79674;
    wire N__79673;
    wire N__79672;
    wire N__79671;
    wire N__79670;
    wire N__79669;
    wire N__79668;
    wire N__79667;
    wire N__79666;
    wire N__79665;
    wire N__79664;
    wire N__79663;
    wire N__79662;
    wire N__79661;
    wire N__79660;
    wire N__79659;
    wire N__79658;
    wire N__79657;
    wire N__79656;
    wire N__79655;
    wire N__79654;
    wire N__79653;
    wire N__79652;
    wire N__79651;
    wire N__79650;
    wire N__79649;
    wire N__79648;
    wire N__79647;
    wire N__79646;
    wire N__79645;
    wire N__79644;
    wire N__79643;
    wire N__79642;
    wire N__79641;
    wire N__79640;
    wire N__79639;
    wire N__79638;
    wire N__79637;
    wire N__79636;
    wire N__79635;
    wire N__79634;
    wire N__79633;
    wire N__79632;
    wire N__79631;
    wire N__79630;
    wire N__79629;
    wire N__79628;
    wire N__79627;
    wire N__79626;
    wire N__79625;
    wire N__79624;
    wire N__79623;
    wire N__79622;
    wire N__79621;
    wire N__79620;
    wire N__79619;
    wire N__79618;
    wire N__79617;
    wire N__79616;
    wire N__79615;
    wire N__79614;
    wire N__79613;
    wire N__79612;
    wire N__79611;
    wire N__79610;
    wire N__79609;
    wire N__79608;
    wire N__79607;
    wire N__79606;
    wire N__79605;
    wire N__79604;
    wire N__79603;
    wire N__79602;
    wire N__79601;
    wire N__79600;
    wire N__79599;
    wire N__79598;
    wire N__79597;
    wire N__79596;
    wire N__79595;
    wire N__79594;
    wire N__79593;
    wire N__79592;
    wire N__79591;
    wire N__79590;
    wire N__79589;
    wire N__79588;
    wire N__79587;
    wire N__79586;
    wire N__79585;
    wire N__79584;
    wire N__79583;
    wire N__79582;
    wire N__79581;
    wire N__79580;
    wire N__79579;
    wire N__79578;
    wire N__79577;
    wire N__79576;
    wire N__79575;
    wire N__79574;
    wire N__79573;
    wire N__79572;
    wire N__79571;
    wire N__79570;
    wire N__79569;
    wire N__79568;
    wire N__79567;
    wire N__79566;
    wire N__79565;
    wire N__79564;
    wire N__79563;
    wire N__79562;
    wire N__79561;
    wire N__79560;
    wire N__79559;
    wire N__79558;
    wire N__79557;
    wire N__79556;
    wire N__79553;
    wire N__79550;
    wire N__79547;
    wire N__79544;
    wire N__79541;
    wire N__79538;
    wire N__79535;
    wire N__79532;
    wire N__79529;
    wire N__79526;
    wire N__79523;
    wire N__79520;
    wire N__79517;
    wire N__79514;
    wire N__79511;
    wire N__79508;
    wire N__79505;
    wire N__79502;
    wire N__79499;
    wire N__79496;
    wire N__79493;
    wire N__79490;
    wire N__79487;
    wire N__79484;
    wire N__79481;
    wire N__79478;
    wire N__79475;
    wire N__79472;
    wire N__79469;
    wire N__79466;
    wire N__79463;
    wire N__79460;
    wire N__79457;
    wire N__79454;
    wire N__79451;
    wire N__79448;
    wire N__79445;
    wire N__79442;
    wire N__79439;
    wire N__79436;
    wire N__79433;
    wire N__79430;
    wire N__79427;
    wire N__79424;
    wire N__79421;
    wire N__79418;
    wire N__79011;
    wire N__79008;
    wire N__79005;
    wire N__79002;
    wire N__78999;
    wire N__78996;
    wire N__78993;
    wire N__78990;
    wire N__78989;
    wire N__78986;
    wire N__78983;
    wire N__78982;
    wire N__78979;
    wire N__78976;
    wire N__78973;
    wire N__78968;
    wire N__78963;
    wire N__78960;
    wire N__78959;
    wire N__78956;
    wire N__78953;
    wire N__78948;
    wire N__78947;
    wire N__78942;
    wire N__78939;
    wire N__78938;
    wire N__78933;
    wire N__78930;
    wire N__78927;
    wire N__78924;
    wire N__78921;
    wire N__78918;
    wire N__78915;
    wire N__78912;
    wire N__78909;
    wire N__78906;
    wire N__78903;
    wire N__78900;
    wire N__78897;
    wire N__78896;
    wire N__78895;
    wire N__78892;
    wire N__78889;
    wire N__78886;
    wire N__78881;
    wire N__78876;
    wire N__78875;
    wire N__78874;
    wire N__78871;
    wire N__78870;
    wire N__78867;
    wire N__78864;
    wire N__78861;
    wire N__78858;
    wire N__78855;
    wire N__78852;
    wire N__78849;
    wire N__78846;
    wire N__78841;
    wire N__78836;
    wire N__78831;
    wire N__78828;
    wire N__78825;
    wire N__78822;
    wire N__78819;
    wire N__78816;
    wire N__78815;
    wire N__78814;
    wire N__78807;
    wire N__78806;
    wire N__78803;
    wire N__78800;
    wire N__78795;
    wire N__78792;
    wire N__78789;
    wire N__78786;
    wire N__78783;
    wire N__78782;
    wire N__78781;
    wire N__78778;
    wire N__78773;
    wire N__78770;
    wire N__78767;
    wire N__78762;
    wire N__78759;
    wire N__78756;
    wire N__78753;
    wire N__78752;
    wire N__78749;
    wire N__78746;
    wire N__78741;
    wire N__78738;
    wire N__78735;
    wire N__78732;
    wire N__78729;
    wire N__78726;
    wire N__78723;
    wire N__78720;
    wire N__78717;
    wire N__78714;
    wire N__78711;
    wire N__78710;
    wire N__78707;
    wire N__78704;
    wire N__78703;
    wire N__78700;
    wire N__78697;
    wire N__78694;
    wire N__78691;
    wire N__78690;
    wire N__78687;
    wire N__78684;
    wire N__78681;
    wire N__78678;
    wire N__78675;
    wire N__78672;
    wire N__78667;
    wire N__78666;
    wire N__78663;
    wire N__78660;
    wire N__78657;
    wire N__78654;
    wire N__78651;
    wire N__78646;
    wire N__78643;
    wire N__78636;
    wire N__78633;
    wire N__78630;
    wire N__78627;
    wire N__78624;
    wire N__78621;
    wire N__78618;
    wire N__78615;
    wire N__78612;
    wire N__78611;
    wire N__78610;
    wire N__78609;
    wire N__78602;
    wire N__78599;
    wire N__78596;
    wire N__78591;
    wire N__78588;
    wire N__78585;
    wire N__78584;
    wire N__78581;
    wire N__78578;
    wire N__78575;
    wire N__78572;
    wire N__78567;
    wire N__78564;
    wire N__78561;
    wire N__78558;
    wire N__78555;
    wire N__78552;
    wire N__78549;
    wire N__78546;
    wire N__78543;
    wire N__78540;
    wire N__78539;
    wire N__78538;
    wire N__78535;
    wire N__78532;
    wire N__78529;
    wire N__78524;
    wire N__78521;
    wire N__78518;
    wire N__78513;
    wire N__78512;
    wire N__78511;
    wire N__78510;
    wire N__78507;
    wire N__78500;
    wire N__78497;
    wire N__78494;
    wire N__78489;
    wire N__78486;
    wire N__78485;
    wire N__78482;
    wire N__78479;
    wire N__78474;
    wire N__78471;
    wire N__78468;
    wire N__78467;
    wire N__78464;
    wire N__78461;
    wire N__78456;
    wire N__78453;
    wire N__78450;
    wire N__78447;
    wire N__78446;
    wire N__78443;
    wire N__78442;
    wire N__78441;
    wire N__78436;
    wire N__78431;
    wire N__78428;
    wire N__78423;
    wire N__78420;
    wire N__78419;
    wire N__78418;
    wire N__78417;
    wire N__78416;
    wire N__78415;
    wire N__78412;
    wire N__78411;
    wire N__78408;
    wire N__78407;
    wire N__78404;
    wire N__78403;
    wire N__78400;
    wire N__78399;
    wire N__78396;
    wire N__78393;
    wire N__78390;
    wire N__78385;
    wire N__78382;
    wire N__78381;
    wire N__78380;
    wire N__78377;
    wire N__78374;
    wire N__78373;
    wire N__78372;
    wire N__78369;
    wire N__78366;
    wire N__78361;
    wire N__78360;
    wire N__78359;
    wire N__78354;
    wire N__78351;
    wire N__78348;
    wire N__78347;
    wire N__78344;
    wire N__78341;
    wire N__78338;
    wire N__78335;
    wire N__78334;
    wire N__78331;
    wire N__78330;
    wire N__78325;
    wire N__78322;
    wire N__78317;
    wire N__78314;
    wire N__78311;
    wire N__78306;
    wire N__78303;
    wire N__78298;
    wire N__78293;
    wire N__78288;
    wire N__78281;
    wire N__78278;
    wire N__78271;
    wire N__78266;
    wire N__78259;
    wire N__78252;
    wire N__78251;
    wire N__78250;
    wire N__78249;
    wire N__78248;
    wire N__78247;
    wire N__78246;
    wire N__78245;
    wire N__78244;
    wire N__78243;
    wire N__78240;
    wire N__78235;
    wire N__78232;
    wire N__78227;
    wire N__78222;
    wire N__78221;
    wire N__78220;
    wire N__78219;
    wire N__78218;
    wire N__78217;
    wire N__78216;
    wire N__78215;
    wire N__78214;
    wire N__78213;
    wire N__78210;
    wire N__78209;
    wire N__78208;
    wire N__78205;
    wire N__78194;
    wire N__78191;
    wire N__78188;
    wire N__78185;
    wire N__78180;
    wire N__78173;
    wire N__78170;
    wire N__78167;
    wire N__78166;
    wire N__78163;
    wire N__78160;
    wire N__78157;
    wire N__78152;
    wire N__78143;
    wire N__78140;
    wire N__78137;
    wire N__78134;
    wire N__78131;
    wire N__78126;
    wire N__78121;
    wire N__78118;
    wire N__78105;
    wire N__78104;
    wire N__78103;
    wire N__78100;
    wire N__78099;
    wire N__78098;
    wire N__78097;
    wire N__78094;
    wire N__78093;
    wire N__78092;
    wire N__78091;
    wire N__78090;
    wire N__78089;
    wire N__78086;
    wire N__78085;
    wire N__78084;
    wire N__78083;
    wire N__78082;
    wire N__78079;
    wire N__78076;
    wire N__78073;
    wire N__78072;
    wire N__78071;
    wire N__78068;
    wire N__78065;
    wire N__78062;
    wire N__78061;
    wire N__78058;
    wire N__78057;
    wire N__78054;
    wire N__78047;
    wire N__78046;
    wire N__78045;
    wire N__78042;
    wire N__78041;
    wire N__78040;
    wire N__78039;
    wire N__78036;
    wire N__78035;
    wire N__78032;
    wire N__78029;
    wire N__78026;
    wire N__78023;
    wire N__78018;
    wire N__78015;
    wire N__78012;
    wire N__78009;
    wire N__78006;
    wire N__78001;
    wire N__77998;
    wire N__77993;
    wire N__77988;
    wire N__77983;
    wire N__77976;
    wire N__77971;
    wire N__77964;
    wire N__77961;
    wire N__77956;
    wire N__77953;
    wire N__77948;
    wire N__77947;
    wire N__77940;
    wire N__77937;
    wire N__77930;
    wire N__77921;
    wire N__77918;
    wire N__77915;
    wire N__77904;
    wire N__77903;
    wire N__77902;
    wire N__77901;
    wire N__77898;
    wire N__77897;
    wire N__77896;
    wire N__77893;
    wire N__77892;
    wire N__77891;
    wire N__77890;
    wire N__77889;
    wire N__77886;
    wire N__77881;
    wire N__77878;
    wire N__77875;
    wire N__77874;
    wire N__77871;
    wire N__77868;
    wire N__77863;
    wire N__77860;
    wire N__77855;
    wire N__77850;
    wire N__77849;
    wire N__77846;
    wire N__77841;
    wire N__77838;
    wire N__77835;
    wire N__77830;
    wire N__77827;
    wire N__77824;
    wire N__77821;
    wire N__77818;
    wire N__77813;
    wire N__77810;
    wire N__77799;
    wire N__77796;
    wire N__77795;
    wire N__77794;
    wire N__77791;
    wire N__77788;
    wire N__77787;
    wire N__77784;
    wire N__77783;
    wire N__77782;
    wire N__77781;
    wire N__77780;
    wire N__77779;
    wire N__77774;
    wire N__77771;
    wire N__77768;
    wire N__77767;
    wire N__77764;
    wire N__77763;
    wire N__77762;
    wire N__77761;
    wire N__77760;
    wire N__77759;
    wire N__77756;
    wire N__77755;
    wire N__77752;
    wire N__77751;
    wire N__77748;
    wire N__77747;
    wire N__77744;
    wire N__77743;
    wire N__77740;
    wire N__77739;
    wire N__77738;
    wire N__77737;
    wire N__77736;
    wire N__77731;
    wire N__77728;
    wire N__77725;
    wire N__77720;
    wire N__77715;
    wire N__77710;
    wire N__77705;
    wire N__77704;
    wire N__77703;
    wire N__77700;
    wire N__77699;
    wire N__77698;
    wire N__77695;
    wire N__77688;
    wire N__77687;
    wire N__77684;
    wire N__77683;
    wire N__77682;
    wire N__77681;
    wire N__77678;
    wire N__77675;
    wire N__77670;
    wire N__77667;
    wire N__77662;
    wire N__77653;
    wire N__77650;
    wire N__77647;
    wire N__77644;
    wire N__77639;
    wire N__77634;
    wire N__77631;
    wire N__77628;
    wire N__77621;
    wire N__77608;
    wire N__77599;
    wire N__77586;
    wire N__77585;
    wire N__77582;
    wire N__77579;
    wire N__77578;
    wire N__77575;
    wire N__77574;
    wire N__77573;
    wire N__77572;
    wire N__77571;
    wire N__77570;
    wire N__77567;
    wire N__77564;
    wire N__77561;
    wire N__77558;
    wire N__77555;
    wire N__77550;
    wire N__77549;
    wire N__77548;
    wire N__77547;
    wire N__77546;
    wire N__77543;
    wire N__77538;
    wire N__77531;
    wire N__77528;
    wire N__77527;
    wire N__77524;
    wire N__77521;
    wire N__77520;
    wire N__77517;
    wire N__77514;
    wire N__77511;
    wire N__77510;
    wire N__77507;
    wire N__77504;
    wire N__77501;
    wire N__77500;
    wire N__77499;
    wire N__77498;
    wire N__77495;
    wire N__77492;
    wire N__77489;
    wire N__77486;
    wire N__77483;
    wire N__77480;
    wire N__77477;
    wire N__77474;
    wire N__77467;
    wire N__77460;
    wire N__77459;
    wire N__77456;
    wire N__77453;
    wire N__77450;
    wire N__77445;
    wire N__77438;
    wire N__77435;
    wire N__77432;
    wire N__77429;
    wire N__77412;
    wire N__77411;
    wire N__77410;
    wire N__77407;
    wire N__77406;
    wire N__77405;
    wire N__77404;
    wire N__77403;
    wire N__77402;
    wire N__77401;
    wire N__77398;
    wire N__77395;
    wire N__77394;
    wire N__77393;
    wire N__77392;
    wire N__77387;
    wire N__77386;
    wire N__77383;
    wire N__77380;
    wire N__77377;
    wire N__77372;
    wire N__77369;
    wire N__77366;
    wire N__77363;
    wire N__77360;
    wire N__77357;
    wire N__77354;
    wire N__77351;
    wire N__77348;
    wire N__77345;
    wire N__77342;
    wire N__77339;
    wire N__77334;
    wire N__77331;
    wire N__77328;
    wire N__77323;
    wire N__77320;
    wire N__77315;
    wire N__77310;
    wire N__77301;
    wire N__77292;
    wire N__77289;
    wire N__77286;
    wire N__77283;
    wire N__77280;
    wire N__77279;
    wire N__77276;
    wire N__77273;
    wire N__77270;
    wire N__77267;
    wire N__77264;
    wire N__77263;
    wire N__77262;
    wire N__77259;
    wire N__77258;
    wire N__77255;
    wire N__77252;
    wire N__77249;
    wire N__77246;
    wire N__77243;
    wire N__77240;
    wire N__77237;
    wire N__77234;
    wire N__77233;
    wire N__77232;
    wire N__77227;
    wire N__77220;
    wire N__77215;
    wire N__77212;
    wire N__77205;
    wire N__77204;
    wire N__77201;
    wire N__77198;
    wire N__77195;
    wire N__77192;
    wire N__77189;
    wire N__77186;
    wire N__77185;
    wire N__77182;
    wire N__77179;
    wire N__77176;
    wire N__77175;
    wire N__77172;
    wire N__77167;
    wire N__77166;
    wire N__77163;
    wire N__77158;
    wire N__77155;
    wire N__77152;
    wire N__77145;
    wire N__77142;
    wire N__77139;
    wire N__77138;
    wire N__77135;
    wire N__77132;
    wire N__77129;
    wire N__77126;
    wire N__77125;
    wire N__77120;
    wire N__77119;
    wire N__77118;
    wire N__77115;
    wire N__77112;
    wire N__77109;
    wire N__77106;
    wire N__77103;
    wire N__77094;
    wire N__77091;
    wire N__77090;
    wire N__77087;
    wire N__77084;
    wire N__77081;
    wire N__77078;
    wire N__77075;
    wire N__77072;
    wire N__77071;
    wire N__77068;
    wire N__77067;
    wire N__77064;
    wire N__77061;
    wire N__77060;
    wire N__77057;
    wire N__77054;
    wire N__77049;
    wire N__77046;
    wire N__77039;
    wire N__77034;
    wire N__77031;
    wire N__77030;
    wire N__77029;
    wire N__77026;
    wire N__77025;
    wire N__77024;
    wire N__77023;
    wire N__77022;
    wire N__77019;
    wire N__77018;
    wire N__77015;
    wire N__77014;
    wire N__77013;
    wire N__77012;
    wire N__77009;
    wire N__77006;
    wire N__77005;
    wire N__77004;
    wire N__77003;
    wire N__77002;
    wire N__76999;
    wire N__76994;
    wire N__76991;
    wire N__76990;
    wire N__76987;
    wire N__76986;
    wire N__76985;
    wire N__76984;
    wire N__76981;
    wire N__76980;
    wire N__76979;
    wire N__76976;
    wire N__76971;
    wire N__76968;
    wire N__76965;
    wire N__76962;
    wire N__76961;
    wire N__76960;
    wire N__76959;
    wire N__76956;
    wire N__76955;
    wire N__76954;
    wire N__76953;
    wire N__76950;
    wire N__76947;
    wire N__76946;
    wire N__76945;
    wire N__76944;
    wire N__76943;
    wire N__76942;
    wire N__76941;
    wire N__76934;
    wire N__76931;
    wire N__76926;
    wire N__76923;
    wire N__76920;
    wire N__76917;
    wire N__76914;
    wire N__76913;
    wire N__76910;
    wire N__76907;
    wire N__76904;
    wire N__76897;
    wire N__76886;
    wire N__76885;
    wire N__76884;
    wire N__76879;
    wire N__76876;
    wire N__76873;
    wire N__76870;
    wire N__76869;
    wire N__76868;
    wire N__76865;
    wire N__76864;
    wire N__76863;
    wire N__76860;
    wire N__76857;
    wire N__76854;
    wire N__76853;
    wire N__76850;
    wire N__76841;
    wire N__76840;
    wire N__76837;
    wire N__76832;
    wire N__76829;
    wire N__76818;
    wire N__76813;
    wire N__76808;
    wire N__76805;
    wire N__76802;
    wire N__76799;
    wire N__76796;
    wire N__76793;
    wire N__76790;
    wire N__76789;
    wire N__76788;
    wire N__76785;
    wire N__76780;
    wire N__76773;
    wire N__76770;
    wire N__76767;
    wire N__76756;
    wire N__76753;
    wire N__76750;
    wire N__76747;
    wire N__76742;
    wire N__76737;
    wire N__76732;
    wire N__76727;
    wire N__76724;
    wire N__76721;
    wire N__76716;
    wire N__76711;
    wire N__76706;
    wire N__76701;
    wire N__76696;
    wire N__76693;
    wire N__76690;
    wire N__76687;
    wire N__76684;
    wire N__76681;
    wire N__76676;
    wire N__76673;
    wire N__76670;
    wire N__76659;
    wire N__76658;
    wire N__76657;
    wire N__76656;
    wire N__76655;
    wire N__76652;
    wire N__76643;
    wire N__76642;
    wire N__76641;
    wire N__76640;
    wire N__76639;
    wire N__76638;
    wire N__76637;
    wire N__76632;
    wire N__76631;
    wire N__76630;
    wire N__76629;
    wire N__76628;
    wire N__76625;
    wire N__76624;
    wire N__76619;
    wire N__76618;
    wire N__76617;
    wire N__76616;
    wire N__76615;
    wire N__76612;
    wire N__76611;
    wire N__76606;
    wire N__76605;
    wire N__76602;
    wire N__76597;
    wire N__76594;
    wire N__76591;
    wire N__76588;
    wire N__76585;
    wire N__76582;
    wire N__76581;
    wire N__76578;
    wire N__76573;
    wire N__76572;
    wire N__76569;
    wire N__76566;
    wire N__76563;
    wire N__76560;
    wire N__76559;
    wire N__76558;
    wire N__76557;
    wire N__76554;
    wire N__76553;
    wire N__76552;
    wire N__76551;
    wire N__76550;
    wire N__76549;
    wire N__76548;
    wire N__76547;
    wire N__76546;
    wire N__76545;
    wire N__76544;
    wire N__76541;
    wire N__76536;
    wire N__76535;
    wire N__76526;
    wire N__76523;
    wire N__76518;
    wire N__76515;
    wire N__76514;
    wire N__76513;
    wire N__76510;
    wire N__76507;
    wire N__76504;
    wire N__76501;
    wire N__76496;
    wire N__76493;
    wire N__76490;
    wire N__76487;
    wire N__76484;
    wire N__76473;
    wire N__76466;
    wire N__76461;
    wire N__76458;
    wire N__76455;
    wire N__76450;
    wire N__76447;
    wire N__76444;
    wire N__76441;
    wire N__76430;
    wire N__76423;
    wire N__76414;
    wire N__76395;
    wire N__76392;
    wire N__76391;
    wire N__76386;
    wire N__76383;
    wire N__76382;
    wire N__76379;
    wire N__76376;
    wire N__76373;
    wire N__76372;
    wire N__76369;
    wire N__76366;
    wire N__76363;
    wire N__76362;
    wire N__76359;
    wire N__76354;
    wire N__76351;
    wire N__76344;
    wire N__76341;
    wire N__76338;
    wire N__76337;
    wire N__76334;
    wire N__76331;
    wire N__76326;
    wire N__76323;
    wire N__76322;
    wire N__76321;
    wire N__76320;
    wire N__76319;
    wire N__76318;
    wire N__76315;
    wire N__76312;
    wire N__76311;
    wire N__76310;
    wire N__76305;
    wire N__76302;
    wire N__76301;
    wire N__76300;
    wire N__76299;
    wire N__76298;
    wire N__76295;
    wire N__76292;
    wire N__76287;
    wire N__76286;
    wire N__76283;
    wire N__76282;
    wire N__76281;
    wire N__76280;
    wire N__76279;
    wire N__76276;
    wire N__76273;
    wire N__76272;
    wire N__76271;
    wire N__76270;
    wire N__76269;
    wire N__76268;
    wire N__76267;
    wire N__76264;
    wire N__76261;
    wire N__76258;
    wire N__76255;
    wire N__76248;
    wire N__76243;
    wire N__76242;
    wire N__76241;
    wire N__76238;
    wire N__76235;
    wire N__76230;
    wire N__76227;
    wire N__76224;
    wire N__76221;
    wire N__76218;
    wire N__76215;
    wire N__76212;
    wire N__76209;
    wire N__76208;
    wire N__76205;
    wire N__76200;
    wire N__76197;
    wire N__76194;
    wire N__76191;
    wire N__76188;
    wire N__76185;
    wire N__76182;
    wire N__76171;
    wire N__76162;
    wire N__76157;
    wire N__76154;
    wire N__76149;
    wire N__76142;
    wire N__76139;
    wire N__76136;
    wire N__76129;
    wire N__76126;
    wire N__76121;
    wire N__76116;
    wire N__76113;
    wire N__76108;
    wire N__76101;
    wire N__76098;
    wire N__76097;
    wire N__76096;
    wire N__76095;
    wire N__76094;
    wire N__76093;
    wire N__76086;
    wire N__76083;
    wire N__76078;
    wire N__76075;
    wire N__76068;
    wire N__76067;
    wire N__76066;
    wire N__76063;
    wire N__76062;
    wire N__76061;
    wire N__76060;
    wire N__76055;
    wire N__76054;
    wire N__76051;
    wire N__76048;
    wire N__76043;
    wire N__76040;
    wire N__76037;
    wire N__76026;
    wire N__76023;
    wire N__76020;
    wire N__76017;
    wire N__76014;
    wire N__76011;
    wire N__76010;
    wire N__76009;
    wire N__76006;
    wire N__76005;
    wire N__76002;
    wire N__75999;
    wire N__75998;
    wire N__75997;
    wire N__75996;
    wire N__75995;
    wire N__75990;
    wire N__75985;
    wire N__75984;
    wire N__75981;
    wire N__75974;
    wire N__75969;
    wire N__75968;
    wire N__75965;
    wire N__75964;
    wire N__75963;
    wire N__75962;
    wire N__75959;
    wire N__75956;
    wire N__75953;
    wire N__75950;
    wire N__75947;
    wire N__75944;
    wire N__75939;
    wire N__75936;
    wire N__75933;
    wire N__75930;
    wire N__75925;
    wire N__75916;
    wire N__75909;
    wire N__75908;
    wire N__75905;
    wire N__75904;
    wire N__75901;
    wire N__75900;
    wire N__75897;
    wire N__75896;
    wire N__75893;
    wire N__75892;
    wire N__75887;
    wire N__75884;
    wire N__75883;
    wire N__75880;
    wire N__75879;
    wire N__75876;
    wire N__75873;
    wire N__75870;
    wire N__75867;
    wire N__75864;
    wire N__75859;
    wire N__75856;
    wire N__75853;
    wire N__75850;
    wire N__75843;
    wire N__75840;
    wire N__75831;
    wire N__75830;
    wire N__75829;
    wire N__75828;
    wire N__75825;
    wire N__75824;
    wire N__75823;
    wire N__75822;
    wire N__75821;
    wire N__75818;
    wire N__75813;
    wire N__75812;
    wire N__75811;
    wire N__75808;
    wire N__75805;
    wire N__75802;
    wire N__75797;
    wire N__75794;
    wire N__75791;
    wire N__75786;
    wire N__75783;
    wire N__75780;
    wire N__75775;
    wire N__75768;
    wire N__75759;
    wire N__75756;
    wire N__75753;
    wire N__75752;
    wire N__75751;
    wire N__75750;
    wire N__75749;
    wire N__75748;
    wire N__75745;
    wire N__75744;
    wire N__75743;
    wire N__75742;
    wire N__75741;
    wire N__75740;
    wire N__75739;
    wire N__75738;
    wire N__75735;
    wire N__75734;
    wire N__75733;
    wire N__75732;
    wire N__75729;
    wire N__75726;
    wire N__75725;
    wire N__75722;
    wire N__75719;
    wire N__75718;
    wire N__75717;
    wire N__75714;
    wire N__75709;
    wire N__75706;
    wire N__75705;
    wire N__75704;
    wire N__75703;
    wire N__75702;
    wire N__75701;
    wire N__75698;
    wire N__75697;
    wire N__75694;
    wire N__75691;
    wire N__75690;
    wire N__75687;
    wire N__75682;
    wire N__75677;
    wire N__75670;
    wire N__75669;
    wire N__75664;
    wire N__75659;
    wire N__75656;
    wire N__75653;
    wire N__75650;
    wire N__75645;
    wire N__75642;
    wire N__75639;
    wire N__75636;
    wire N__75631;
    wire N__75628;
    wire N__75623;
    wire N__75620;
    wire N__75613;
    wire N__75610;
    wire N__75607;
    wire N__75604;
    wire N__75597;
    wire N__75594;
    wire N__75585;
    wire N__75580;
    wire N__75573;
    wire N__75568;
    wire N__75565;
    wire N__75558;
    wire N__75555;
    wire N__75546;
    wire N__75543;
    wire N__75540;
    wire N__75537;
    wire N__75536;
    wire N__75535;
    wire N__75534;
    wire N__75533;
    wire N__75532;
    wire N__75529;
    wire N__75528;
    wire N__75525;
    wire N__75522;
    wire N__75519;
    wire N__75518;
    wire N__75515;
    wire N__75512;
    wire N__75509;
    wire N__75508;
    wire N__75505;
    wire N__75500;
    wire N__75495;
    wire N__75492;
    wire N__75489;
    wire N__75488;
    wire N__75485;
    wire N__75482;
    wire N__75481;
    wire N__75478;
    wire N__75477;
    wire N__75476;
    wire N__75475;
    wire N__75474;
    wire N__75465;
    wire N__75462;
    wire N__75459;
    wire N__75456;
    wire N__75453;
    wire N__75450;
    wire N__75445;
    wire N__75442;
    wire N__75439;
    wire N__75434;
    wire N__75429;
    wire N__75426;
    wire N__75423;
    wire N__75420;
    wire N__75417;
    wire N__75410;
    wire N__75403;
    wire N__75400;
    wire N__75397;
    wire N__75390;
    wire N__75387;
    wire N__75384;
    wire N__75381;
    wire N__75378;
    wire N__75375;
    wire N__75372;
    wire N__75369;
    wire N__75368;
    wire N__75367;
    wire N__75366;
    wire N__75363;
    wire N__75360;
    wire N__75357;
    wire N__75356;
    wire N__75353;
    wire N__75348;
    wire N__75345;
    wire N__75344;
    wire N__75341;
    wire N__75338;
    wire N__75333;
    wire N__75332;
    wire N__75331;
    wire N__75330;
    wire N__75329;
    wire N__75326;
    wire N__75323;
    wire N__75318;
    wire N__75315;
    wire N__75312;
    wire N__75309;
    wire N__75306;
    wire N__75305;
    wire N__75302;
    wire N__75301;
    wire N__75294;
    wire N__75291;
    wire N__75290;
    wire N__75289;
    wire N__75284;
    wire N__75281;
    wire N__75278;
    wire N__75275;
    wire N__75272;
    wire N__75269;
    wire N__75266;
    wire N__75263;
    wire N__75260;
    wire N__75255;
    wire N__75250;
    wire N__75247;
    wire N__75240;
    wire N__75237;
    wire N__75234;
    wire N__75225;
    wire N__75222;
    wire N__75219;
    wire N__75216;
    wire N__75213;
    wire N__75210;
    wire N__75207;
    wire N__75204;
    wire N__75201;
    wire N__75198;
    wire N__75197;
    wire N__75194;
    wire N__75193;
    wire N__75192;
    wire N__75189;
    wire N__75186;
    wire N__75185;
    wire N__75184;
    wire N__75181;
    wire N__75178;
    wire N__75175;
    wire N__75172;
    wire N__75167;
    wire N__75164;
    wire N__75161;
    wire N__75158;
    wire N__75153;
    wire N__75150;
    wire N__75147;
    wire N__75138;
    wire N__75135;
    wire N__75134;
    wire N__75131;
    wire N__75130;
    wire N__75129;
    wire N__75128;
    wire N__75125;
    wire N__75122;
    wire N__75119;
    wire N__75118;
    wire N__75113;
    wire N__75110;
    wire N__75107;
    wire N__75102;
    wire N__75099;
    wire N__75096;
    wire N__75091;
    wire N__75088;
    wire N__75081;
    wire N__75078;
    wire N__75075;
    wire N__75074;
    wire N__75073;
    wire N__75070;
    wire N__75069;
    wire N__75068;
    wire N__75065;
    wire N__75062;
    wire N__75059;
    wire N__75054;
    wire N__75051;
    wire N__75050;
    wire N__75047;
    wire N__75042;
    wire N__75039;
    wire N__75036;
    wire N__75027;
    wire N__75024;
    wire N__75023;
    wire N__75020;
    wire N__75017;
    wire N__75016;
    wire N__75015;
    wire N__75014;
    wire N__75011;
    wire N__75008;
    wire N__75007;
    wire N__75004;
    wire N__75001;
    wire N__74998;
    wire N__74995;
    wire N__74992;
    wire N__74989;
    wire N__74986;
    wire N__74981;
    wire N__74978;
    wire N__74967;
    wire N__74964;
    wire N__74961;
    wire N__74958;
    wire N__74955;
    wire N__74952;
    wire N__74949;
    wire N__74948;
    wire N__74945;
    wire N__74940;
    wire N__74937;
    wire N__74934;
    wire N__74931;
    wire N__74930;
    wire N__74929;
    wire N__74928;
    wire N__74927;
    wire N__74926;
    wire N__74925;
    wire N__74924;
    wire N__74923;
    wire N__74922;
    wire N__74921;
    wire N__74918;
    wire N__74915;
    wire N__74912;
    wire N__74907;
    wire N__74906;
    wire N__74905;
    wire N__74904;
    wire N__74901;
    wire N__74896;
    wire N__74889;
    wire N__74886;
    wire N__74885;
    wire N__74884;
    wire N__74883;
    wire N__74880;
    wire N__74875;
    wire N__74872;
    wire N__74869;
    wire N__74868;
    wire N__74865;
    wire N__74858;
    wire N__74855;
    wire N__74848;
    wire N__74845;
    wire N__74844;
    wire N__74843;
    wire N__74842;
    wire N__74841;
    wire N__74838;
    wire N__74835;
    wire N__74832;
    wire N__74829;
    wire N__74826;
    wire N__74823;
    wire N__74820;
    wire N__74817;
    wire N__74814;
    wire N__74811;
    wire N__74804;
    wire N__74795;
    wire N__74792;
    wire N__74785;
    wire N__74772;
    wire N__74769;
    wire N__74768;
    wire N__74767;
    wire N__74764;
    wire N__74761;
    wire N__74758;
    wire N__74757;
    wire N__74756;
    wire N__74751;
    wire N__74750;
    wire N__74747;
    wire N__74742;
    wire N__74739;
    wire N__74736;
    wire N__74735;
    wire N__74734;
    wire N__74729;
    wire N__74726;
    wire N__74723;
    wire N__74720;
    wire N__74717;
    wire N__74714;
    wire N__74703;
    wire N__74700;
    wire N__74699;
    wire N__74694;
    wire N__74691;
    wire N__74688;
    wire N__74685;
    wire N__74682;
    wire N__74679;
    wire N__74676;
    wire N__74673;
    wire N__74670;
    wire N__74667;
    wire N__74664;
    wire N__74661;
    wire N__74658;
    wire N__74657;
    wire N__74656;
    wire N__74655;
    wire N__74652;
    wire N__74649;
    wire N__74646;
    wire N__74643;
    wire N__74642;
    wire N__74637;
    wire N__74634;
    wire N__74631;
    wire N__74630;
    wire N__74629;
    wire N__74628;
    wire N__74625;
    wire N__74624;
    wire N__74621;
    wire N__74616;
    wire N__74613;
    wire N__74608;
    wire N__74603;
    wire N__74592;
    wire N__74591;
    wire N__74590;
    wire N__74587;
    wire N__74584;
    wire N__74583;
    wire N__74582;
    wire N__74579;
    wire N__74576;
    wire N__74575;
    wire N__74574;
    wire N__74571;
    wire N__74566;
    wire N__74561;
    wire N__74558;
    wire N__74557;
    wire N__74554;
    wire N__74549;
    wire N__74548;
    wire N__74547;
    wire N__74544;
    wire N__74541;
    wire N__74538;
    wire N__74533;
    wire N__74528;
    wire N__74525;
    wire N__74514;
    wire N__74513;
    wire N__74510;
    wire N__74509;
    wire N__74506;
    wire N__74503;
    wire N__74502;
    wire N__74499;
    wire N__74496;
    wire N__74493;
    wire N__74490;
    wire N__74489;
    wire N__74486;
    wire N__74483;
    wire N__74482;
    wire N__74481;
    wire N__74480;
    wire N__74479;
    wire N__74476;
    wire N__74473;
    wire N__74470;
    wire N__74467;
    wire N__74464;
    wire N__74461;
    wire N__74458;
    wire N__74455;
    wire N__74452;
    wire N__74445;
    wire N__74442;
    wire N__74439;
    wire N__74424;
    wire N__74421;
    wire N__74420;
    wire N__74419;
    wire N__74418;
    wire N__74413;
    wire N__74410;
    wire N__74409;
    wire N__74408;
    wire N__74405;
    wire N__74404;
    wire N__74403;
    wire N__74402;
    wire N__74399;
    wire N__74394;
    wire N__74391;
    wire N__74388;
    wire N__74387;
    wire N__74384;
    wire N__74383;
    wire N__74382;
    wire N__74381;
    wire N__74376;
    wire N__74371;
    wire N__74368;
    wire N__74365;
    wire N__74362;
    wire N__74359;
    wire N__74356;
    wire N__74351;
    wire N__74348;
    wire N__74345;
    wire N__74342;
    wire N__74339;
    wire N__74322;
    wire N__74319;
    wire N__74316;
    wire N__74313;
    wire N__74310;
    wire N__74307;
    wire N__74304;
    wire N__74301;
    wire N__74298;
    wire N__74295;
    wire N__74292;
    wire N__74289;
    wire N__74286;
    wire N__74283;
    wire N__74280;
    wire N__74277;
    wire N__74274;
    wire N__74271;
    wire N__74268;
    wire N__74265;
    wire N__74262;
    wire N__74259;
    wire N__74256;
    wire N__74253;
    wire N__74250;
    wire N__74247;
    wire N__74244;
    wire N__74241;
    wire N__74238;
    wire N__74235;
    wire N__74232;
    wire N__74229;
    wire N__74226;
    wire N__74223;
    wire N__74220;
    wire N__74217;
    wire N__74214;
    wire N__74211;
    wire N__74208;
    wire N__74205;
    wire N__74202;
    wire N__74199;
    wire N__74196;
    wire N__74193;
    wire N__74190;
    wire N__74189;
    wire N__74188;
    wire N__74185;
    wire N__74182;
    wire N__74181;
    wire N__74178;
    wire N__74177;
    wire N__74176;
    wire N__74173;
    wire N__74170;
    wire N__74167;
    wire N__74166;
    wire N__74165;
    wire N__74164;
    wire N__74161;
    wire N__74156;
    wire N__74153;
    wire N__74152;
    wire N__74149;
    wire N__74146;
    wire N__74139;
    wire N__74134;
    wire N__74131;
    wire N__74128;
    wire N__74123;
    wire N__74118;
    wire N__74109;
    wire N__74106;
    wire N__74103;
    wire N__74100;
    wire N__74097;
    wire N__74094;
    wire N__74093;
    wire N__74092;
    wire N__74089;
    wire N__74084;
    wire N__74079;
    wire N__74076;
    wire N__74073;
    wire N__74072;
    wire N__74071;
    wire N__74068;
    wire N__74067;
    wire N__74064;
    wire N__74063;
    wire N__74060;
    wire N__74057;
    wire N__74056;
    wire N__74053;
    wire N__74050;
    wire N__74049;
    wire N__74048;
    wire N__74045;
    wire N__74042;
    wire N__74039;
    wire N__74038;
    wire N__74035;
    wire N__74030;
    wire N__74025;
    wire N__74022;
    wire N__74019;
    wire N__74016;
    wire N__74013;
    wire N__74006;
    wire N__74001;
    wire N__73998;
    wire N__73989;
    wire N__73986;
    wire N__73983;
    wire N__73980;
    wire N__73977;
    wire N__73974;
    wire N__73973;
    wire N__73970;
    wire N__73967;
    wire N__73962;
    wire N__73959;
    wire N__73956;
    wire N__73953;
    wire N__73950;
    wire N__73947;
    wire N__73944;
    wire N__73941;
    wire N__73940;
    wire N__73935;
    wire N__73932;
    wire N__73929;
    wire N__73926;
    wire N__73923;
    wire N__73920;
    wire N__73917;
    wire N__73914;
    wire N__73911;
    wire N__73908;
    wire N__73905;
    wire N__73902;
    wire N__73899;
    wire N__73896;
    wire N__73893;
    wire N__73890;
    wire N__73887;
    wire N__73884;
    wire N__73881;
    wire N__73878;
    wire N__73877;
    wire N__73874;
    wire N__73873;
    wire N__73872;
    wire N__73869;
    wire N__73868;
    wire N__73867;
    wire N__73864;
    wire N__73861;
    wire N__73858;
    wire N__73855;
    wire N__73850;
    wire N__73847;
    wire N__73844;
    wire N__73839;
    wire N__73836;
    wire N__73833;
    wire N__73830;
    wire N__73825;
    wire N__73818;
    wire N__73815;
    wire N__73812;
    wire N__73809;
    wire N__73806;
    wire N__73803;
    wire N__73800;
    wire N__73797;
    wire N__73794;
    wire N__73791;
    wire N__73788;
    wire N__73785;
    wire N__73782;
    wire N__73779;
    wire N__73776;
    wire N__73773;
    wire N__73770;
    wire N__73767;
    wire N__73764;
    wire N__73761;
    wire N__73758;
    wire N__73755;
    wire N__73752;
    wire N__73749;
    wire N__73746;
    wire N__73743;
    wire N__73740;
    wire N__73737;
    wire N__73734;
    wire N__73731;
    wire N__73728;
    wire N__73725;
    wire N__73722;
    wire N__73721;
    wire N__73718;
    wire N__73715;
    wire N__73710;
    wire N__73707;
    wire N__73704;
    wire N__73701;
    wire N__73698;
    wire N__73695;
    wire N__73692;
    wire N__73691;
    wire N__73688;
    wire N__73685;
    wire N__73682;
    wire N__73679;
    wire N__73674;
    wire N__73671;
    wire N__73668;
    wire N__73665;
    wire N__73662;
    wire N__73659;
    wire N__73656;
    wire N__73655;
    wire N__73652;
    wire N__73651;
    wire N__73650;
    wire N__73647;
    wire N__73646;
    wire N__73643;
    wire N__73640;
    wire N__73639;
    wire N__73638;
    wire N__73635;
    wire N__73632;
    wire N__73629;
    wire N__73628;
    wire N__73627;
    wire N__73626;
    wire N__73623;
    wire N__73620;
    wire N__73617;
    wire N__73614;
    wire N__73611;
    wire N__73606;
    wire N__73605;
    wire N__73602;
    wire N__73599;
    wire N__73596;
    wire N__73591;
    wire N__73590;
    wire N__73585;
    wire N__73580;
    wire N__73579;
    wire N__73576;
    wire N__73573;
    wire N__73570;
    wire N__73567;
    wire N__73564;
    wire N__73563;
    wire N__73560;
    wire N__73555;
    wire N__73552;
    wire N__73547;
    wire N__73540;
    wire N__73537;
    wire N__73534;
    wire N__73529;
    wire N__73522;
    wire N__73515;
    wire N__73514;
    wire N__73513;
    wire N__73510;
    wire N__73505;
    wire N__73500;
    wire N__73499;
    wire N__73494;
    wire N__73491;
    wire N__73488;
    wire N__73485;
    wire N__73482;
    wire N__73481;
    wire N__73478;
    wire N__73475;
    wire N__73470;
    wire N__73467;
    wire N__73466;
    wire N__73465;
    wire N__73462;
    wire N__73459;
    wire N__73456;
    wire N__73449;
    wire N__73446;
    wire N__73443;
    wire N__73440;
    wire N__73437;
    wire N__73434;
    wire N__73431;
    wire N__73430;
    wire N__73427;
    wire N__73424;
    wire N__73419;
    wire N__73416;
    wire N__73413;
    wire N__73412;
    wire N__73411;
    wire N__73408;
    wire N__73403;
    wire N__73398;
    wire N__73395;
    wire N__73392;
    wire N__73389;
    wire N__73386;
    wire N__73385;
    wire N__73382;
    wire N__73379;
    wire N__73374;
    wire N__73373;
    wire N__73372;
    wire N__73367;
    wire N__73364;
    wire N__73359;
    wire N__73356;
    wire N__73353;
    wire N__73350;
    wire N__73349;
    wire N__73346;
    wire N__73343;
    wire N__73342;
    wire N__73339;
    wire N__73336;
    wire N__73333;
    wire N__73326;
    wire N__73325;
    wire N__73322;
    wire N__73319;
    wire N__73314;
    wire N__73313;
    wire N__73310;
    wire N__73307;
    wire N__73302;
    wire N__73299;
    wire N__73296;
    wire N__73293;
    wire N__73290;
    wire N__73289;
    wire N__73286;
    wire N__73285;
    wire N__73282;
    wire N__73279;
    wire N__73276;
    wire N__73273;
    wire N__73270;
    wire N__73267;
    wire N__73264;
    wire N__73257;
    wire N__73254;
    wire N__73253;
    wire N__73250;
    wire N__73247;
    wire N__73242;
    wire N__73239;
    wire N__73236;
    wire N__73233;
    wire N__73230;
    wire N__73229;
    wire N__73226;
    wire N__73223;
    wire N__73218;
    wire N__73215;
    wire N__73212;
    wire N__73211;
    wire N__73210;
    wire N__73209;
    wire N__73208;
    wire N__73207;
    wire N__73206;
    wire N__73205;
    wire N__73204;
    wire N__73201;
    wire N__73198;
    wire N__73195;
    wire N__73194;
    wire N__73191;
    wire N__73190;
    wire N__73187;
    wire N__73186;
    wire N__73183;
    wire N__73182;
    wire N__73179;
    wire N__73176;
    wire N__73167;
    wire N__73162;
    wire N__73157;
    wire N__73154;
    wire N__73149;
    wire N__73144;
    wire N__73141;
    wire N__73136;
    wire N__73131;
    wire N__73128;
    wire N__73125;
    wire N__73120;
    wire N__73113;
    wire N__73112;
    wire N__73107;
    wire N__73104;
    wire N__73103;
    wire N__73100;
    wire N__73097;
    wire N__73094;
    wire N__73091;
    wire N__73088;
    wire N__73085;
    wire N__73080;
    wire N__73077;
    wire N__73074;
    wire N__73071;
    wire N__73068;
    wire N__73065;
    wire N__73062;
    wire N__73059;
    wire N__73058;
    wire N__73055;
    wire N__73052;
    wire N__73049;
    wire N__73044;
    wire N__73043;
    wire N__73040;
    wire N__73037;
    wire N__73034;
    wire N__73031;
    wire N__73030;
    wire N__73027;
    wire N__73024;
    wire N__73021;
    wire N__73014;
    wire N__73013;
    wire N__73008;
    wire N__73005;
    wire N__73002;
    wire N__73001;
    wire N__72998;
    wire N__72995;
    wire N__72992;
    wire N__72989;
    wire N__72984;
    wire N__72981;
    wire N__72978;
    wire N__72975;
    wire N__72972;
    wire N__72969;
    wire N__72966;
    wire N__72963;
    wire N__72962;
    wire N__72959;
    wire N__72956;
    wire N__72951;
    wire N__72950;
    wire N__72945;
    wire N__72942;
    wire N__72939;
    wire N__72936;
    wire N__72933;
    wire N__72932;
    wire N__72931;
    wire N__72928;
    wire N__72923;
    wire N__72920;
    wire N__72917;
    wire N__72912;
    wire N__72909;
    wire N__72906;
    wire N__72903;
    wire N__72900;
    wire N__72899;
    wire N__72896;
    wire N__72893;
    wire N__72892;
    wire N__72889;
    wire N__72886;
    wire N__72883;
    wire N__72880;
    wire N__72877;
    wire N__72870;
    wire N__72867;
    wire N__72866;
    wire N__72863;
    wire N__72860;
    wire N__72855;
    wire N__72852;
    wire N__72849;
    wire N__72848;
    wire N__72845;
    wire N__72842;
    wire N__72837;
    wire N__72834;
    wire N__72831;
    wire N__72828;
    wire N__72827;
    wire N__72826;
    wire N__72823;
    wire N__72820;
    wire N__72817;
    wire N__72814;
    wire N__72811;
    wire N__72808;
    wire N__72805;
    wire N__72802;
    wire N__72795;
    wire N__72792;
    wire N__72789;
    wire N__72788;
    wire N__72785;
    wire N__72782;
    wire N__72777;
    wire N__72774;
    wire N__72771;
    wire N__72768;
    wire N__72765;
    wire N__72762;
    wire N__72759;
    wire N__72756;
    wire N__72753;
    wire N__72750;
    wire N__72747;
    wire N__72744;
    wire N__72741;
    wire N__72738;
    wire N__72735;
    wire N__72732;
    wire N__72729;
    wire N__72726;
    wire N__72723;
    wire N__72720;
    wire N__72719;
    wire N__72716;
    wire N__72713;
    wire N__72710;
    wire N__72707;
    wire N__72704;
    wire N__72699;
    wire N__72696;
    wire N__72693;
    wire N__72692;
    wire N__72689;
    wire N__72686;
    wire N__72685;
    wire N__72680;
    wire N__72677;
    wire N__72674;
    wire N__72669;
    wire N__72666;
    wire N__72663;
    wire N__72660;
    wire N__72657;
    wire N__72656;
    wire N__72655;
    wire N__72654;
    wire N__72651;
    wire N__72648;
    wire N__72645;
    wire N__72644;
    wire N__72643;
    wire N__72642;
    wire N__72641;
    wire N__72638;
    wire N__72637;
    wire N__72624;
    wire N__72621;
    wire N__72620;
    wire N__72619;
    wire N__72618;
    wire N__72615;
    wire N__72614;
    wire N__72613;
    wire N__72610;
    wire N__72607;
    wire N__72604;
    wire N__72601;
    wire N__72596;
    wire N__72593;
    wire N__72588;
    wire N__72587;
    wire N__72584;
    wire N__72581;
    wire N__72570;
    wire N__72567;
    wire N__72562;
    wire N__72559;
    wire N__72552;
    wire N__72549;
    wire N__72548;
    wire N__72545;
    wire N__72544;
    wire N__72541;
    wire N__72538;
    wire N__72533;
    wire N__72530;
    wire N__72527;
    wire N__72522;
    wire N__72521;
    wire N__72520;
    wire N__72519;
    wire N__72510;
    wire N__72507;
    wire N__72504;
    wire N__72501;
    wire N__72498;
    wire N__72495;
    wire N__72492;
    wire N__72489;
    wire N__72486;
    wire N__72485;
    wire N__72482;
    wire N__72481;
    wire N__72478;
    wire N__72475;
    wire N__72472;
    wire N__72469;
    wire N__72466;
    wire N__72463;
    wire N__72460;
    wire N__72453;
    wire N__72450;
    wire N__72447;
    wire N__72444;
    wire N__72441;
    wire N__72438;
    wire N__72435;
    wire N__72432;
    wire N__72429;
    wire N__72426;
    wire N__72423;
    wire N__72422;
    wire N__72419;
    wire N__72418;
    wire N__72417;
    wire N__72416;
    wire N__72415;
    wire N__72414;
    wire N__72413;
    wire N__72412;
    wire N__72409;
    wire N__72408;
    wire N__72407;
    wire N__72406;
    wire N__72403;
    wire N__72400;
    wire N__72397;
    wire N__72394;
    wire N__72391;
    wire N__72390;
    wire N__72387;
    wire N__72384;
    wire N__72381;
    wire N__72378;
    wire N__72375;
    wire N__72372;
    wire N__72369;
    wire N__72360;
    wire N__72357;
    wire N__72354;
    wire N__72353;
    wire N__72350;
    wire N__72347;
    wire N__72342;
    wire N__72339;
    wire N__72336;
    wire N__72331;
    wire N__72326;
    wire N__72323;
    wire N__72320;
    wire N__72317;
    wire N__72314;
    wire N__72311;
    wire N__72308;
    wire N__72303;
    wire N__72300;
    wire N__72297;
    wire N__72292;
    wire N__72289;
    wire N__72284;
    wire N__72273;
    wire N__72270;
    wire N__72267;
    wire N__72264;
    wire N__72263;
    wire N__72262;
    wire N__72259;
    wire N__72254;
    wire N__72251;
    wire N__72248;
    wire N__72245;
    wire N__72242;
    wire N__72237;
    wire N__72236;
    wire N__72233;
    wire N__72230;
    wire N__72227;
    wire N__72224;
    wire N__72223;
    wire N__72218;
    wire N__72215;
    wire N__72210;
    wire N__72207;
    wire N__72204;
    wire N__72203;
    wire N__72200;
    wire N__72197;
    wire N__72192;
    wire N__72189;
    wire N__72186;
    wire N__72185;
    wire N__72182;
    wire N__72179;
    wire N__72174;
    wire N__72171;
    wire N__72168;
    wire N__72167;
    wire N__72166;
    wire N__72161;
    wire N__72158;
    wire N__72153;
    wire N__72152;
    wire N__72149;
    wire N__72146;
    wire N__72143;
    wire N__72140;
    wire N__72137;
    wire N__72134;
    wire N__72133;
    wire N__72132;
    wire N__72131;
    wire N__72130;
    wire N__72127;
    wire N__72124;
    wire N__72121;
    wire N__72120;
    wire N__72117;
    wire N__72112;
    wire N__72111;
    wire N__72110;
    wire N__72107;
    wire N__72102;
    wire N__72099;
    wire N__72094;
    wire N__72093;
    wire N__72088;
    wire N__72083;
    wire N__72078;
    wire N__72075;
    wire N__72072;
    wire N__72063;
    wire N__72062;
    wire N__72061;
    wire N__72058;
    wire N__72057;
    wire N__72054;
    wire N__72053;
    wire N__72052;
    wire N__72051;
    wire N__72050;
    wire N__72047;
    wire N__72046;
    wire N__72045;
    wire N__72044;
    wire N__72041;
    wire N__72040;
    wire N__72039;
    wire N__72038;
    wire N__72037;
    wire N__72036;
    wire N__72033;
    wire N__72032;
    wire N__72027;
    wire N__72022;
    wire N__72017;
    wire N__72012;
    wire N__72009;
    wire N__72008;
    wire N__72005;
    wire N__72002;
    wire N__71997;
    wire N__71992;
    wire N__71989;
    wire N__71988;
    wire N__71987;
    wire N__71984;
    wire N__71981;
    wire N__71978;
    wire N__71975;
    wire N__71974;
    wire N__71971;
    wire N__71970;
    wire N__71969;
    wire N__71968;
    wire N__71967;
    wire N__71966;
    wire N__71963;
    wire N__71960;
    wire N__71953;
    wire N__71950;
    wire N__71947;
    wire N__71944;
    wire N__71939;
    wire N__71936;
    wire N__71931;
    wire N__71928;
    wire N__71925;
    wire N__71922;
    wire N__71917;
    wire N__71912;
    wire N__71903;
    wire N__71896;
    wire N__71891;
    wire N__71874;
    wire N__71871;
    wire N__71868;
    wire N__71865;
    wire N__71862;
    wire N__71859;
    wire N__71856;
    wire N__71853;
    wire N__71850;
    wire N__71847;
    wire N__71844;
    wire N__71841;
    wire N__71838;
    wire N__71837;
    wire N__71834;
    wire N__71833;
    wire N__71830;
    wire N__71827;
    wire N__71824;
    wire N__71821;
    wire N__71818;
    wire N__71815;
    wire N__71810;
    wire N__71805;
    wire N__71804;
    wire N__71801;
    wire N__71798;
    wire N__71797;
    wire N__71794;
    wire N__71791;
    wire N__71788;
    wire N__71783;
    wire N__71780;
    wire N__71777;
    wire N__71772;
    wire N__71771;
    wire N__71768;
    wire N__71767;
    wire N__71764;
    wire N__71761;
    wire N__71758;
    wire N__71755;
    wire N__71752;
    wire N__71749;
    wire N__71744;
    wire N__71741;
    wire N__71738;
    wire N__71733;
    wire N__71732;
    wire N__71727;
    wire N__71726;
    wire N__71723;
    wire N__71720;
    wire N__71717;
    wire N__71712;
    wire N__71711;
    wire N__71710;
    wire N__71709;
    wire N__71708;
    wire N__71705;
    wire N__71702;
    wire N__71701;
    wire N__71694;
    wire N__71689;
    wire N__71686;
    wire N__71683;
    wire N__71678;
    wire N__71675;
    wire N__71670;
    wire N__71669;
    wire N__71666;
    wire N__71663;
    wire N__71662;
    wire N__71659;
    wire N__71656;
    wire N__71653;
    wire N__71650;
    wire N__71647;
    wire N__71644;
    wire N__71641;
    wire N__71634;
    wire N__71631;
    wire N__71630;
    wire N__71627;
    wire N__71624;
    wire N__71623;
    wire N__71620;
    wire N__71617;
    wire N__71614;
    wire N__71611;
    wire N__71608;
    wire N__71605;
    wire N__71602;
    wire N__71595;
    wire N__71592;
    wire N__71591;
    wire N__71590;
    wire N__71587;
    wire N__71584;
    wire N__71581;
    wire N__71578;
    wire N__71573;
    wire N__71570;
    wire N__71567;
    wire N__71562;
    wire N__71561;
    wire N__71560;
    wire N__71559;
    wire N__71558;
    wire N__71557;
    wire N__71556;
    wire N__71553;
    wire N__71552;
    wire N__71551;
    wire N__71550;
    wire N__71549;
    wire N__71548;
    wire N__71547;
    wire N__71546;
    wire N__71545;
    wire N__71544;
    wire N__71537;
    wire N__71532;
    wire N__71531;
    wire N__71530;
    wire N__71527;
    wire N__71526;
    wire N__71525;
    wire N__71520;
    wire N__71519;
    wire N__71518;
    wire N__71517;
    wire N__71516;
    wire N__71513;
    wire N__71510;
    wire N__71509;
    wire N__71506;
    wire N__71503;
    wire N__71502;
    wire N__71501;
    wire N__71498;
    wire N__71495;
    wire N__71490;
    wire N__71485;
    wire N__71482;
    wire N__71481;
    wire N__71480;
    wire N__71477;
    wire N__71474;
    wire N__71469;
    wire N__71466;
    wire N__71461;
    wire N__71460;
    wire N__71455;
    wire N__71450;
    wire N__71447;
    wire N__71444;
    wire N__71441;
    wire N__71438;
    wire N__71435;
    wire N__71428;
    wire N__71425;
    wire N__71418;
    wire N__71415;
    wire N__71412;
    wire N__71407;
    wire N__71404;
    wire N__71401;
    wire N__71396;
    wire N__71393;
    wire N__71390;
    wire N__71387;
    wire N__71380;
    wire N__71375;
    wire N__71368;
    wire N__71363;
    wire N__71358;
    wire N__71355;
    wire N__71350;
    wire N__71345;
    wire N__71340;
    wire N__71331;
    wire N__71328;
    wire N__71325;
    wire N__71322;
    wire N__71319;
    wire N__71316;
    wire N__71313;
    wire N__71310;
    wire N__71307;
    wire N__71306;
    wire N__71305;
    wire N__71304;
    wire N__71301;
    wire N__71298;
    wire N__71293;
    wire N__71286;
    wire N__71283;
    wire N__71282;
    wire N__71281;
    wire N__71278;
    wire N__71275;
    wire N__71272;
    wire N__71271;
    wire N__71266;
    wire N__71265;
    wire N__71262;
    wire N__71259;
    wire N__71256;
    wire N__71253;
    wire N__71246;
    wire N__71243;
    wire N__71238;
    wire N__71235;
    wire N__71232;
    wire N__71229;
    wire N__71226;
    wire N__71223;
    wire N__71220;
    wire N__71219;
    wire N__71218;
    wire N__71211;
    wire N__71208;
    wire N__71205;
    wire N__71202;
    wire N__71199;
    wire N__71198;
    wire N__71195;
    wire N__71192;
    wire N__71189;
    wire N__71188;
    wire N__71185;
    wire N__71184;
    wire N__71183;
    wire N__71180;
    wire N__71179;
    wire N__71176;
    wire N__71175;
    wire N__71174;
    wire N__71171;
    wire N__71170;
    wire N__71169;
    wire N__71168;
    wire N__71167;
    wire N__71162;
    wire N__71159;
    wire N__71156;
    wire N__71153;
    wire N__71148;
    wire N__71145;
    wire N__71140;
    wire N__71137;
    wire N__71134;
    wire N__71133;
    wire N__71132;
    wire N__71131;
    wire N__71130;
    wire N__71129;
    wire N__71128;
    wire N__71125;
    wire N__71124;
    wire N__71123;
    wire N__71122;
    wire N__71113;
    wire N__71110;
    wire N__71103;
    wire N__71098;
    wire N__71089;
    wire N__71086;
    wire N__71079;
    wire N__71076;
    wire N__71071;
    wire N__71066;
    wire N__71055;
    wire N__71052;
    wire N__71049;
    wire N__71046;
    wire N__71043;
    wire N__71040;
    wire N__71037;
    wire N__71036;
    wire N__71033;
    wire N__71030;
    wire N__71025;
    wire N__71022;
    wire N__71021;
    wire N__71020;
    wire N__71017;
    wire N__71016;
    wire N__71013;
    wire N__71010;
    wire N__71007;
    wire N__71004;
    wire N__71001;
    wire N__70998;
    wire N__70995;
    wire N__70992;
    wire N__70989;
    wire N__70980;
    wire N__70979;
    wire N__70978;
    wire N__70977;
    wire N__70974;
    wire N__70973;
    wire N__70970;
    wire N__70969;
    wire N__70968;
    wire N__70965;
    wire N__70964;
    wire N__70961;
    wire N__70958;
    wire N__70957;
    wire N__70954;
    wire N__70951;
    wire N__70946;
    wire N__70943;
    wire N__70940;
    wire N__70937;
    wire N__70934;
    wire N__70929;
    wire N__70928;
    wire N__70923;
    wire N__70920;
    wire N__70915;
    wire N__70910;
    wire N__70907;
    wire N__70904;
    wire N__70903;
    wire N__70902;
    wire N__70899;
    wire N__70894;
    wire N__70891;
    wire N__70888;
    wire N__70885;
    wire N__70882;
    wire N__70869;
    wire N__70868;
    wire N__70865;
    wire N__70862;
    wire N__70859;
    wire N__70858;
    wire N__70857;
    wire N__70854;
    wire N__70851;
    wire N__70848;
    wire N__70845;
    wire N__70836;
    wire N__70833;
    wire N__70830;
    wire N__70827;
    wire N__70824;
    wire N__70821;
    wire N__70818;
    wire N__70815;
    wire N__70812;
    wire N__70809;
    wire N__70806;
    wire N__70803;
    wire N__70800;
    wire N__70797;
    wire N__70794;
    wire N__70791;
    wire N__70788;
    wire N__70785;
    wire N__70782;
    wire N__70779;
    wire N__70776;
    wire N__70773;
    wire N__70770;
    wire N__70767;
    wire N__70764;
    wire N__70761;
    wire N__70758;
    wire N__70755;
    wire N__70752;
    wire N__70749;
    wire N__70746;
    wire N__70743;
    wire N__70740;
    wire N__70737;
    wire N__70734;
    wire N__70731;
    wire N__70728;
    wire N__70725;
    wire N__70722;
    wire N__70719;
    wire N__70716;
    wire N__70713;
    wire N__70710;
    wire N__70709;
    wire N__70704;
    wire N__70703;
    wire N__70700;
    wire N__70697;
    wire N__70694;
    wire N__70691;
    wire N__70686;
    wire N__70683;
    wire N__70680;
    wire N__70677;
    wire N__70676;
    wire N__70675;
    wire N__70672;
    wire N__70669;
    wire N__70666;
    wire N__70663;
    wire N__70660;
    wire N__70657;
    wire N__70652;
    wire N__70649;
    wire N__70646;
    wire N__70643;
    wire N__70638;
    wire N__70635;
    wire N__70634;
    wire N__70633;
    wire N__70630;
    wire N__70625;
    wire N__70622;
    wire N__70619;
    wire N__70616;
    wire N__70613;
    wire N__70610;
    wire N__70607;
    wire N__70602;
    wire N__70601;
    wire N__70596;
    wire N__70593;
    wire N__70590;
    wire N__70587;
    wire N__70584;
    wire N__70581;
    wire N__70580;
    wire N__70579;
    wire N__70576;
    wire N__70573;
    wire N__70572;
    wire N__70569;
    wire N__70566;
    wire N__70563;
    wire N__70560;
    wire N__70557;
    wire N__70548;
    wire N__70545;
    wire N__70542;
    wire N__70539;
    wire N__70536;
    wire N__70535;
    wire N__70532;
    wire N__70529;
    wire N__70524;
    wire N__70521;
    wire N__70518;
    wire N__70515;
    wire N__70512;
    wire N__70509;
    wire N__70508;
    wire N__70505;
    wire N__70502;
    wire N__70499;
    wire N__70494;
    wire N__70491;
    wire N__70490;
    wire N__70487;
    wire N__70484;
    wire N__70483;
    wire N__70482;
    wire N__70479;
    wire N__70476;
    wire N__70473;
    wire N__70472;
    wire N__70471;
    wire N__70470;
    wire N__70469;
    wire N__70468;
    wire N__70467;
    wire N__70464;
    wire N__70457;
    wire N__70454;
    wire N__70453;
    wire N__70450;
    wire N__70447;
    wire N__70444;
    wire N__70441;
    wire N__70438;
    wire N__70435;
    wire N__70432;
    wire N__70429;
    wire N__70428;
    wire N__70427;
    wire N__70424;
    wire N__70421;
    wire N__70416;
    wire N__70413;
    wire N__70410;
    wire N__70407;
    wire N__70402;
    wire N__70399;
    wire N__70396;
    wire N__70393;
    wire N__70390;
    wire N__70387;
    wire N__70384;
    wire N__70377;
    wire N__70362;
    wire N__70359;
    wire N__70358;
    wire N__70357;
    wire N__70356;
    wire N__70355;
    wire N__70354;
    wire N__70353;
    wire N__70352;
    wire N__70351;
    wire N__70350;
    wire N__70349;
    wire N__70348;
    wire N__70347;
    wire N__70346;
    wire N__70343;
    wire N__70314;
    wire N__70311;
    wire N__70308;
    wire N__70307;
    wire N__70302;
    wire N__70299;
    wire N__70296;
    wire N__70293;
    wire N__70290;
    wire N__70289;
    wire N__70286;
    wire N__70283;
    wire N__70278;
    wire N__70275;
    wire N__70272;
    wire N__70271;
    wire N__70270;
    wire N__70263;
    wire N__70260;
    wire N__70257;
    wire N__70254;
    wire N__70251;
    wire N__70248;
    wire N__70245;
    wire N__70242;
    wire N__70239;
    wire N__70236;
    wire N__70233;
    wire N__70230;
    wire N__70227;
    wire N__70224;
    wire N__70221;
    wire N__70218;
    wire N__70215;
    wire N__70212;
    wire N__70209;
    wire N__70206;
    wire N__70203;
    wire N__70202;
    wire N__70199;
    wire N__70196;
    wire N__70193;
    wire N__70190;
    wire N__70185;
    wire N__70182;
    wire N__70179;
    wire N__70176;
    wire N__70173;
    wire N__70170;
    wire N__70167;
    wire N__70164;
    wire N__70161;
    wire N__70158;
    wire N__70155;
    wire N__70152;
    wire N__70149;
    wire N__70148;
    wire N__70147;
    wire N__70144;
    wire N__70139;
    wire N__70134;
    wire N__70133;
    wire N__70128;
    wire N__70125;
    wire N__70122;
    wire N__70119;
    wire N__70116;
    wire N__70113;
    wire N__70110;
    wire N__70107;
    wire N__70104;
    wire N__70101;
    wire N__70098;
    wire N__70095;
    wire N__70092;
    wire N__70091;
    wire N__70090;
    wire N__70087;
    wire N__70084;
    wire N__70081;
    wire N__70074;
    wire N__70073;
    wire N__70072;
    wire N__70065;
    wire N__70062;
    wire N__70059;
    wire N__70056;
    wire N__70053;
    wire N__70050;
    wire N__70047;
    wire N__70044;
    wire N__70041;
    wire N__70038;
    wire N__70035;
    wire N__70032;
    wire N__70029;
    wire N__70026;
    wire N__70023;
    wire N__70020;
    wire N__70017;
    wire N__70014;
    wire N__70011;
    wire N__70010;
    wire N__70007;
    wire N__70006;
    wire N__70005;
    wire N__70002;
    wire N__70001;
    wire N__70000;
    wire N__69999;
    wire N__69998;
    wire N__69997;
    wire N__69996;
    wire N__69995;
    wire N__69994;
    wire N__69993;
    wire N__69992;
    wire N__69991;
    wire N__69990;
    wire N__69989;
    wire N__69988;
    wire N__69985;
    wire N__69980;
    wire N__69973;
    wire N__69956;
    wire N__69951;
    wire N__69946;
    wire N__69943;
    wire N__69938;
    wire N__69935;
    wire N__69930;
    wire N__69925;
    wire N__69922;
    wire N__69919;
    wire N__69916;
    wire N__69909;
    wire N__69908;
    wire N__69905;
    wire N__69902;
    wire N__69901;
    wire N__69900;
    wire N__69899;
    wire N__69898;
    wire N__69897;
    wire N__69896;
    wire N__69895;
    wire N__69894;
    wire N__69893;
    wire N__69892;
    wire N__69891;
    wire N__69888;
    wire N__69885;
    wire N__69858;
    wire N__69855;
    wire N__69852;
    wire N__69849;
    wire N__69846;
    wire N__69843;
    wire N__69840;
    wire N__69837;
    wire N__69836;
    wire N__69833;
    wire N__69830;
    wire N__69827;
    wire N__69826;
    wire N__69823;
    wire N__69820;
    wire N__69817;
    wire N__69814;
    wire N__69807;
    wire N__69804;
    wire N__69801;
    wire N__69798;
    wire N__69795;
    wire N__69792;
    wire N__69789;
    wire N__69788;
    wire N__69787;
    wire N__69784;
    wire N__69779;
    wire N__69774;
    wire N__69771;
    wire N__69768;
    wire N__69765;
    wire N__69762;
    wire N__69759;
    wire N__69756;
    wire N__69753;
    wire N__69750;
    wire N__69747;
    wire N__69744;
    wire N__69741;
    wire N__69738;
    wire N__69735;
    wire N__69732;
    wire N__69729;
    wire N__69726;
    wire N__69723;
    wire N__69720;
    wire N__69717;
    wire N__69714;
    wire N__69711;
    wire N__69708;
    wire N__69705;
    wire N__69702;
    wire N__69699;
    wire N__69696;
    wire N__69693;
    wire N__69690;
    wire N__69687;
    wire N__69684;
    wire N__69681;
    wire N__69678;
    wire N__69675;
    wire N__69672;
    wire N__69669;
    wire N__69666;
    wire N__69663;
    wire N__69660;
    wire N__69657;
    wire N__69654;
    wire N__69651;
    wire N__69648;
    wire N__69645;
    wire N__69642;
    wire N__69639;
    wire N__69636;
    wire N__69633;
    wire N__69630;
    wire N__69627;
    wire N__69624;
    wire N__69621;
    wire N__69618;
    wire N__69615;
    wire N__69612;
    wire N__69609;
    wire N__69606;
    wire N__69603;
    wire N__69600;
    wire N__69597;
    wire N__69594;
    wire N__69591;
    wire N__69588;
    wire N__69585;
    wire N__69582;
    wire N__69579;
    wire N__69576;
    wire N__69573;
    wire N__69570;
    wire N__69567;
    wire N__69564;
    wire N__69561;
    wire N__69558;
    wire N__69555;
    wire N__69552;
    wire N__69549;
    wire N__69546;
    wire N__69543;
    wire N__69540;
    wire N__69537;
    wire N__69534;
    wire N__69531;
    wire N__69528;
    wire N__69525;
    wire N__69522;
    wire N__69519;
    wire N__69516;
    wire N__69513;
    wire N__69510;
    wire N__69507;
    wire N__69504;
    wire N__69501;
    wire N__69500;
    wire N__69499;
    wire N__69498;
    wire N__69497;
    wire N__69494;
    wire N__69489;
    wire N__69484;
    wire N__69479;
    wire N__69476;
    wire N__69473;
    wire N__69470;
    wire N__69465;
    wire N__69462;
    wire N__69459;
    wire N__69456;
    wire N__69453;
    wire N__69450;
    wire N__69447;
    wire N__69444;
    wire N__69441;
    wire N__69438;
    wire N__69435;
    wire N__69432;
    wire N__69429;
    wire N__69426;
    wire N__69423;
    wire N__69420;
    wire N__69417;
    wire N__69416;
    wire N__69413;
    wire N__69412;
    wire N__69411;
    wire N__69408;
    wire N__69405;
    wire N__69402;
    wire N__69399;
    wire N__69396;
    wire N__69389;
    wire N__69386;
    wire N__69383;
    wire N__69378;
    wire N__69375;
    wire N__69374;
    wire N__69373;
    wire N__69370;
    wire N__69367;
    wire N__69366;
    wire N__69363;
    wire N__69358;
    wire N__69355;
    wire N__69348;
    wire N__69345;
    wire N__69342;
    wire N__69339;
    wire N__69336;
    wire N__69333;
    wire N__69330;
    wire N__69327;
    wire N__69324;
    wire N__69321;
    wire N__69318;
    wire N__69315;
    wire N__69312;
    wire N__69311;
    wire N__69308;
    wire N__69305;
    wire N__69302;
    wire N__69297;
    wire N__69294;
    wire N__69291;
    wire N__69288;
    wire N__69285;
    wire N__69284;
    wire N__69281;
    wire N__69278;
    wire N__69275;
    wire N__69272;
    wire N__69269;
    wire N__69266;
    wire N__69261;
    wire N__69258;
    wire N__69255;
    wire N__69252;
    wire N__69251;
    wire N__69248;
    wire N__69245;
    wire N__69240;
    wire N__69237;
    wire N__69236;
    wire N__69235;
    wire N__69232;
    wire N__69229;
    wire N__69226;
    wire N__69223;
    wire N__69218;
    wire N__69213;
    wire N__69210;
    wire N__69209;
    wire N__69208;
    wire N__69201;
    wire N__69198;
    wire N__69195;
    wire N__69194;
    wire N__69191;
    wire N__69188;
    wire N__69185;
    wire N__69184;
    wire N__69181;
    wire N__69178;
    wire N__69175;
    wire N__69172;
    wire N__69167;
    wire N__69164;
    wire N__69161;
    wire N__69156;
    wire N__69153;
    wire N__69150;
    wire N__69147;
    wire N__69146;
    wire N__69145;
    wire N__69142;
    wire N__69139;
    wire N__69136;
    wire N__69131;
    wire N__69128;
    wire N__69125;
    wire N__69120;
    wire N__69117;
    wire N__69116;
    wire N__69115;
    wire N__69110;
    wire N__69107;
    wire N__69104;
    wire N__69101;
    wire N__69098;
    wire N__69093;
    wire N__69090;
    wire N__69089;
    wire N__69086;
    wire N__69085;
    wire N__69082;
    wire N__69079;
    wire N__69076;
    wire N__69073;
    wire N__69070;
    wire N__69067;
    wire N__69064;
    wire N__69061;
    wire N__69058;
    wire N__69055;
    wire N__69048;
    wire N__69045;
    wire N__69044;
    wire N__69039;
    wire N__69036;
    wire N__69035;
    wire N__69030;
    wire N__69027;
    wire N__69024;
    wire N__69023;
    wire N__69018;
    wire N__69015;
    wire N__69014;
    wire N__69011;
    wire N__69008;
    wire N__69005;
    wire N__69002;
    wire N__68999;
    wire N__68994;
    wire N__68991;
    wire N__68990;
    wire N__68989;
    wire N__68986;
    wire N__68983;
    wire N__68980;
    wire N__68973;
    wire N__68970;
    wire N__68967;
    wire N__68964;
    wire N__68961;
    wire N__68960;
    wire N__68957;
    wire N__68954;
    wire N__68949;
    wire N__68946;
    wire N__68943;
    wire N__68940;
    wire N__68939;
    wire N__68936;
    wire N__68933;
    wire N__68928;
    wire N__68925;
    wire N__68924;
    wire N__68923;
    wire N__68920;
    wire N__68915;
    wire N__68910;
    wire N__68907;
    wire N__68904;
    wire N__68903;
    wire N__68902;
    wire N__68901;
    wire N__68896;
    wire N__68891;
    wire N__68888;
    wire N__68887;
    wire N__68884;
    wire N__68881;
    wire N__68878;
    wire N__68875;
    wire N__68870;
    wire N__68867;
    wire N__68864;
    wire N__68859;
    wire N__68856;
    wire N__68853;
    wire N__68850;
    wire N__68847;
    wire N__68844;
    wire N__68843;
    wire N__68840;
    wire N__68837;
    wire N__68836;
    wire N__68831;
    wire N__68828;
    wire N__68825;
    wire N__68820;
    wire N__68819;
    wire N__68816;
    wire N__68815;
    wire N__68814;
    wire N__68813;
    wire N__68808;
    wire N__68805;
    wire N__68800;
    wire N__68795;
    wire N__68792;
    wire N__68789;
    wire N__68786;
    wire N__68783;
    wire N__68778;
    wire N__68775;
    wire N__68772;
    wire N__68769;
    wire N__68768;
    wire N__68767;
    wire N__68766;
    wire N__68763;
    wire N__68762;
    wire N__68759;
    wire N__68758;
    wire N__68755;
    wire N__68752;
    wire N__68751;
    wire N__68748;
    wire N__68745;
    wire N__68744;
    wire N__68741;
    wire N__68738;
    wire N__68735;
    wire N__68732;
    wire N__68729;
    wire N__68724;
    wire N__68721;
    wire N__68716;
    wire N__68711;
    wire N__68708;
    wire N__68703;
    wire N__68700;
    wire N__68697;
    wire N__68694;
    wire N__68691;
    wire N__68686;
    wire N__68681;
    wire N__68676;
    wire N__68675;
    wire N__68674;
    wire N__68671;
    wire N__68670;
    wire N__68667;
    wire N__68664;
    wire N__68661;
    wire N__68660;
    wire N__68657;
    wire N__68654;
    wire N__68651;
    wire N__68648;
    wire N__68645;
    wire N__68642;
    wire N__68637;
    wire N__68632;
    wire N__68629;
    wire N__68626;
    wire N__68625;
    wire N__68620;
    wire N__68617;
    wire N__68614;
    wire N__68607;
    wire N__68604;
    wire N__68601;
    wire N__68598;
    wire N__68595;
    wire N__68594;
    wire N__68591;
    wire N__68588;
    wire N__68585;
    wire N__68584;
    wire N__68581;
    wire N__68578;
    wire N__68575;
    wire N__68572;
    wire N__68569;
    wire N__68562;
    wire N__68559;
    wire N__68556;
    wire N__68555;
    wire N__68554;
    wire N__68551;
    wire N__68548;
    wire N__68545;
    wire N__68538;
    wire N__68535;
    wire N__68532;
    wire N__68529;
    wire N__68526;
    wire N__68523;
    wire N__68520;
    wire N__68517;
    wire N__68516;
    wire N__68513;
    wire N__68510;
    wire N__68507;
    wire N__68506;
    wire N__68501;
    wire N__68498;
    wire N__68493;
    wire N__68490;
    wire N__68487;
    wire N__68484;
    wire N__68481;
    wire N__68480;
    wire N__68479;
    wire N__68476;
    wire N__68473;
    wire N__68470;
    wire N__68467;
    wire N__68464;
    wire N__68457;
    wire N__68456;
    wire N__68455;
    wire N__68452;
    wire N__68449;
    wire N__68446;
    wire N__68439;
    wire N__68436;
    wire N__68435;
    wire N__68434;
    wire N__68431;
    wire N__68428;
    wire N__68425;
    wire N__68422;
    wire N__68419;
    wire N__68412;
    wire N__68411;
    wire N__68410;
    wire N__68407;
    wire N__68404;
    wire N__68401;
    wire N__68394;
    wire N__68391;
    wire N__68388;
    wire N__68385;
    wire N__68382;
    wire N__68379;
    wire N__68376;
    wire N__68373;
    wire N__68370;
    wire N__68367;
    wire N__68366;
    wire N__68365;
    wire N__68362;
    wire N__68359;
    wire N__68356;
    wire N__68353;
    wire N__68348;
    wire N__68345;
    wire N__68342;
    wire N__68337;
    wire N__68336;
    wire N__68333;
    wire N__68330;
    wire N__68327;
    wire N__68322;
    wire N__68319;
    wire N__68318;
    wire N__68317;
    wire N__68314;
    wire N__68309;
    wire N__68304;
    wire N__68301;
    wire N__68298;
    wire N__68295;
    wire N__68294;
    wire N__68291;
    wire N__68290;
    wire N__68287;
    wire N__68284;
    wire N__68281;
    wire N__68280;
    wire N__68277;
    wire N__68274;
    wire N__68271;
    wire N__68268;
    wire N__68265;
    wire N__68260;
    wire N__68253;
    wire N__68250;
    wire N__68249;
    wire N__68246;
    wire N__68243;
    wire N__68240;
    wire N__68237;
    wire N__68234;
    wire N__68231;
    wire N__68226;
    wire N__68223;
    wire N__68220;
    wire N__68217;
    wire N__68214;
    wire N__68211;
    wire N__68208;
    wire N__68205;
    wire N__68202;
    wire N__68199;
    wire N__68196;
    wire N__68193;
    wire N__68190;
    wire N__68187;
    wire N__68184;
    wire N__68181;
    wire N__68178;
    wire N__68175;
    wire N__68172;
    wire N__68171;
    wire N__68170;
    wire N__68167;
    wire N__68164;
    wire N__68161;
    wire N__68158;
    wire N__68155;
    wire N__68152;
    wire N__68149;
    wire N__68146;
    wire N__68139;
    wire N__68136;
    wire N__68133;
    wire N__68130;
    wire N__68127;
    wire N__68124;
    wire N__68121;
    wire N__68118;
    wire N__68115;
    wire N__68112;
    wire N__68109;
    wire N__68106;
    wire N__68103;
    wire N__68100;
    wire N__68097;
    wire N__68096;
    wire N__68091;
    wire N__68088;
    wire N__68085;
    wire N__68082;
    wire N__68079;
    wire N__68076;
    wire N__68073;
    wire N__68070;
    wire N__68067;
    wire N__68064;
    wire N__68063;
    wire N__68060;
    wire N__68057;
    wire N__68052;
    wire N__68049;
    wire N__68046;
    wire N__68043;
    wire N__68040;
    wire N__68037;
    wire N__68034;
    wire N__68031;
    wire N__68028;
    wire N__68025;
    wire N__68022;
    wire N__68019;
    wire N__68016;
    wire N__68013;
    wire N__68010;
    wire N__68007;
    wire N__68004;
    wire N__68001;
    wire N__67998;
    wire N__67995;
    wire N__67992;
    wire N__67989;
    wire N__67988;
    wire N__67983;
    wire N__67980;
    wire N__67977;
    wire N__67974;
    wire N__67971;
    wire N__67968;
    wire N__67965;
    wire N__67962;
    wire N__67959;
    wire N__67956;
    wire N__67953;
    wire N__67950;
    wire N__67947;
    wire N__67944;
    wire N__67941;
    wire N__67938;
    wire N__67935;
    wire N__67932;
    wire N__67929;
    wire N__67928;
    wire N__67925;
    wire N__67922;
    wire N__67917;
    wire N__67914;
    wire N__67911;
    wire N__67908;
    wire N__67905;
    wire N__67902;
    wire N__67899;
    wire N__67896;
    wire N__67893;
    wire N__67890;
    wire N__67887;
    wire N__67884;
    wire N__67881;
    wire N__67878;
    wire N__67875;
    wire N__67872;
    wire N__67869;
    wire N__67866;
    wire N__67863;
    wire N__67860;
    wire N__67857;
    wire N__67854;
    wire N__67851;
    wire N__67850;
    wire N__67847;
    wire N__67846;
    wire N__67845;
    wire N__67842;
    wire N__67839;
    wire N__67838;
    wire N__67835;
    wire N__67832;
    wire N__67829;
    wire N__67826;
    wire N__67823;
    wire N__67816;
    wire N__67813;
    wire N__67806;
    wire N__67805;
    wire N__67802;
    wire N__67799;
    wire N__67796;
    wire N__67793;
    wire N__67790;
    wire N__67789;
    wire N__67788;
    wire N__67785;
    wire N__67784;
    wire N__67781;
    wire N__67778;
    wire N__67775;
    wire N__67772;
    wire N__67769;
    wire N__67762;
    wire N__67755;
    wire N__67754;
    wire N__67751;
    wire N__67748;
    wire N__67747;
    wire N__67746;
    wire N__67743;
    wire N__67740;
    wire N__67739;
    wire N__67736;
    wire N__67733;
    wire N__67730;
    wire N__67727;
    wire N__67726;
    wire N__67723;
    wire N__67718;
    wire N__67715;
    wire N__67712;
    wire N__67709;
    wire N__67706;
    wire N__67703;
    wire N__67700;
    wire N__67697;
    wire N__67686;
    wire N__67683;
    wire N__67682;
    wire N__67679;
    wire N__67676;
    wire N__67673;
    wire N__67670;
    wire N__67669;
    wire N__67668;
    wire N__67667;
    wire N__67664;
    wire N__67663;
    wire N__67662;
    wire N__67659;
    wire N__67656;
    wire N__67651;
    wire N__67648;
    wire N__67645;
    wire N__67642;
    wire N__67639;
    wire N__67638;
    wire N__67635;
    wire N__67632;
    wire N__67629;
    wire N__67622;
    wire N__67619;
    wire N__67616;
    wire N__67609;
    wire N__67602;
    wire N__67599;
    wire N__67596;
    wire N__67593;
    wire N__67590;
    wire N__67587;
    wire N__67586;
    wire N__67583;
    wire N__67580;
    wire N__67579;
    wire N__67574;
    wire N__67571;
    wire N__67570;
    wire N__67569;
    wire N__67566;
    wire N__67563;
    wire N__67558;
    wire N__67555;
    wire N__67550;
    wire N__67547;
    wire N__67544;
    wire N__67539;
    wire N__67536;
    wire N__67533;
    wire N__67532;
    wire N__67529;
    wire N__67526;
    wire N__67523;
    wire N__67520;
    wire N__67519;
    wire N__67516;
    wire N__67513;
    wire N__67510;
    wire N__67507;
    wire N__67502;
    wire N__67497;
    wire N__67494;
    wire N__67491;
    wire N__67488;
    wire N__67487;
    wire N__67484;
    wire N__67481;
    wire N__67478;
    wire N__67473;
    wire N__67470;
    wire N__67467;
    wire N__67464;
    wire N__67461;
    wire N__67458;
    wire N__67455;
    wire N__67452;
    wire N__67449;
    wire N__67446;
    wire N__67443;
    wire N__67440;
    wire N__67437;
    wire N__67434;
    wire N__67431;
    wire N__67430;
    wire N__67427;
    wire N__67424;
    wire N__67421;
    wire N__67416;
    wire N__67415;
    wire N__67412;
    wire N__67409;
    wire N__67406;
    wire N__67405;
    wire N__67404;
    wire N__67401;
    wire N__67398;
    wire N__67397;
    wire N__67392;
    wire N__67391;
    wire N__67390;
    wire N__67387;
    wire N__67384;
    wire N__67381;
    wire N__67380;
    wire N__67377;
    wire N__67374;
    wire N__67371;
    wire N__67368;
    wire N__67365;
    wire N__67360;
    wire N__67357;
    wire N__67350;
    wire N__67347;
    wire N__67338;
    wire N__67335;
    wire N__67334;
    wire N__67331;
    wire N__67330;
    wire N__67327;
    wire N__67324;
    wire N__67321;
    wire N__67320;
    wire N__67317;
    wire N__67314;
    wire N__67313;
    wire N__67308;
    wire N__67307;
    wire N__67306;
    wire N__67305;
    wire N__67302;
    wire N__67299;
    wire N__67296;
    wire N__67293;
    wire N__67290;
    wire N__67287;
    wire N__67284;
    wire N__67281;
    wire N__67278;
    wire N__67273;
    wire N__67262;
    wire N__67257;
    wire N__67254;
    wire N__67253;
    wire N__67250;
    wire N__67247;
    wire N__67244;
    wire N__67241;
    wire N__67238;
    wire N__67237;
    wire N__67234;
    wire N__67233;
    wire N__67230;
    wire N__67227;
    wire N__67224;
    wire N__67221;
    wire N__67216;
    wire N__67215;
    wire N__67214;
    wire N__67209;
    wire N__67206;
    wire N__67201;
    wire N__67194;
    wire N__67191;
    wire N__67188;
    wire N__67185;
    wire N__67184;
    wire N__67183;
    wire N__67180;
    wire N__67179;
    wire N__67176;
    wire N__67173;
    wire N__67170;
    wire N__67167;
    wire N__67166;
    wire N__67165;
    wire N__67164;
    wire N__67163;
    wire N__67160;
    wire N__67157;
    wire N__67154;
    wire N__67151;
    wire N__67146;
    wire N__67141;
    wire N__67138;
    wire N__67133;
    wire N__67122;
    wire N__67119;
    wire N__67116;
    wire N__67115;
    wire N__67112;
    wire N__67109;
    wire N__67108;
    wire N__67107;
    wire N__67104;
    wire N__67101;
    wire N__67098;
    wire N__67095;
    wire N__67092;
    wire N__67087;
    wire N__67084;
    wire N__67081;
    wire N__67078;
    wire N__67071;
    wire N__67068;
    wire N__67067;
    wire N__67066;
    wire N__67065;
    wire N__67062;
    wire N__67055;
    wire N__67050;
    wire N__67047;
    wire N__67044;
    wire N__67043;
    wire N__67040;
    wire N__67037;
    wire N__67034;
    wire N__67029;
    wire N__67026;
    wire N__67023;
    wire N__67020;
    wire N__67019;
    wire N__67016;
    wire N__67013;
    wire N__67008;
    wire N__67005;
    wire N__67002;
    wire N__66999;
    wire N__66996;
    wire N__66993;
    wire N__66990;
    wire N__66987;
    wire N__66984;
    wire N__66981;
    wire N__66978;
    wire N__66975;
    wire N__66972;
    wire N__66969;
    wire N__66966;
    wire N__66963;
    wire N__66960;
    wire N__66957;
    wire N__66954;
    wire N__66951;
    wire N__66948;
    wire N__66945;
    wire N__66942;
    wire N__66939;
    wire N__66936;
    wire N__66933;
    wire N__66930;
    wire N__66927;
    wire N__66926;
    wire N__66923;
    wire N__66920;
    wire N__66917;
    wire N__66912;
    wire N__66909;
    wire N__66908;
    wire N__66903;
    wire N__66900;
    wire N__66897;
    wire N__66894;
    wire N__66891;
    wire N__66888;
    wire N__66885;
    wire N__66882;
    wire N__66879;
    wire N__66876;
    wire N__66873;
    wire N__66870;
    wire N__66867;
    wire N__66864;
    wire N__66861;
    wire N__66858;
    wire N__66855;
    wire N__66852;
    wire N__66849;
    wire N__66846;
    wire N__66843;
    wire N__66842;
    wire N__66841;
    wire N__66838;
    wire N__66833;
    wire N__66830;
    wire N__66827;
    wire N__66822;
    wire N__66819;
    wire N__66818;
    wire N__66813;
    wire N__66810;
    wire N__66807;
    wire N__66806;
    wire N__66805;
    wire N__66804;
    wire N__66803;
    wire N__66802;
    wire N__66801;
    wire N__66800;
    wire N__66797;
    wire N__66796;
    wire N__66793;
    wire N__66792;
    wire N__66789;
    wire N__66788;
    wire N__66785;
    wire N__66784;
    wire N__66781;
    wire N__66780;
    wire N__66777;
    wire N__66776;
    wire N__66775;
    wire N__66772;
    wire N__66771;
    wire N__66760;
    wire N__66743;
    wire N__66736;
    wire N__66729;
    wire N__66726;
    wire N__66723;
    wire N__66722;
    wire N__66721;
    wire N__66718;
    wire N__66715;
    wire N__66712;
    wire N__66709;
    wire N__66706;
    wire N__66699;
    wire N__66698;
    wire N__66695;
    wire N__66690;
    wire N__66687;
    wire N__66684;
    wire N__66681;
    wire N__66678;
    wire N__66675;
    wire N__66672;
    wire N__66669;
    wire N__66666;
    wire N__66663;
    wire N__66660;
    wire N__66657;
    wire N__66654;
    wire N__66651;
    wire N__66648;
    wire N__66645;
    wire N__66642;
    wire N__66639;
    wire N__66636;
    wire N__66633;
    wire N__66630;
    wire N__66627;
    wire N__66624;
    wire N__66621;
    wire N__66618;
    wire N__66615;
    wire N__66612;
    wire N__66609;
    wire N__66606;
    wire N__66603;
    wire N__66600;
    wire N__66597;
    wire N__66594;
    wire N__66591;
    wire N__66588;
    wire N__66585;
    wire N__66582;
    wire N__66579;
    wire N__66576;
    wire N__66573;
    wire N__66570;
    wire N__66567;
    wire N__66564;
    wire N__66561;
    wire N__66558;
    wire N__66555;
    wire N__66552;
    wire N__66549;
    wire N__66546;
    wire N__66543;
    wire N__66540;
    wire N__66537;
    wire N__66534;
    wire N__66531;
    wire N__66528;
    wire N__66525;
    wire N__66522;
    wire N__66519;
    wire N__66516;
    wire N__66513;
    wire N__66510;
    wire N__66507;
    wire N__66506;
    wire N__66505;
    wire N__66502;
    wire N__66497;
    wire N__66494;
    wire N__66491;
    wire N__66488;
    wire N__66485;
    wire N__66480;
    wire N__66477;
    wire N__66474;
    wire N__66471;
    wire N__66468;
    wire N__66467;
    wire N__66466;
    wire N__66463;
    wire N__66460;
    wire N__66457;
    wire N__66454;
    wire N__66449;
    wire N__66446;
    wire N__66443;
    wire N__66438;
    wire N__66435;
    wire N__66432;
    wire N__66429;
    wire N__66426;
    wire N__66425;
    wire N__66424;
    wire N__66419;
    wire N__66416;
    wire N__66413;
    wire N__66410;
    wire N__66407;
    wire N__66402;
    wire N__66399;
    wire N__66396;
    wire N__66393;
    wire N__66390;
    wire N__66387;
    wire N__66384;
    wire N__66381;
    wire N__66378;
    wire N__66375;
    wire N__66372;
    wire N__66369;
    wire N__66366;
    wire N__66363;
    wire N__66360;
    wire N__66357;
    wire N__66354;
    wire N__66351;
    wire N__66348;
    wire N__66345;
    wire N__66342;
    wire N__66339;
    wire N__66336;
    wire N__66333;
    wire N__66330;
    wire N__66327;
    wire N__66324;
    wire N__66323;
    wire N__66320;
    wire N__66317;
    wire N__66312;
    wire N__66311;
    wire N__66308;
    wire N__66307;
    wire N__66304;
    wire N__66299;
    wire N__66296;
    wire N__66291;
    wire N__66290;
    wire N__66289;
    wire N__66288;
    wire N__66287;
    wire N__66286;
    wire N__66281;
    wire N__66276;
    wire N__66271;
    wire N__66266;
    wire N__66261;
    wire N__66258;
    wire N__66255;
    wire N__66254;
    wire N__66251;
    wire N__66248;
    wire N__66243;
    wire N__66240;
    wire N__66239;
    wire N__66236;
    wire N__66233;
    wire N__66230;
    wire N__66227;
    wire N__66222;
    wire N__66219;
    wire N__66216;
    wire N__66213;
    wire N__66210;
    wire N__66207;
    wire N__66204;
    wire N__66201;
    wire N__66198;
    wire N__66195;
    wire N__66192;
    wire N__66189;
    wire N__66186;
    wire N__66183;
    wire N__66180;
    wire N__66177;
    wire N__66174;
    wire N__66171;
    wire N__66168;
    wire N__66165;
    wire N__66162;
    wire N__66159;
    wire N__66156;
    wire N__66153;
    wire N__66150;
    wire N__66147;
    wire N__66144;
    wire N__66141;
    wire N__66138;
    wire N__66135;
    wire N__66132;
    wire N__66129;
    wire N__66126;
    wire N__66125;
    wire N__66124;
    wire N__66119;
    wire N__66116;
    wire N__66113;
    wire N__66108;
    wire N__66107;
    wire N__66104;
    wire N__66101;
    wire N__66100;
    wire N__66097;
    wire N__66094;
    wire N__66093;
    wire N__66090;
    wire N__66085;
    wire N__66082;
    wire N__66079;
    wire N__66074;
    wire N__66071;
    wire N__66068;
    wire N__66063;
    wire N__66060;
    wire N__66057;
    wire N__66054;
    wire N__66051;
    wire N__66048;
    wire N__66045;
    wire N__66044;
    wire N__66043;
    wire N__66040;
    wire N__66039;
    wire N__66038;
    wire N__66037;
    wire N__66034;
    wire N__66031;
    wire N__66028;
    wire N__66025;
    wire N__66022;
    wire N__66019;
    wire N__66016;
    wire N__66013;
    wire N__66008;
    wire N__66005;
    wire N__66004;
    wire N__66001;
    wire N__65998;
    wire N__65995;
    wire N__65994;
    wire N__65991;
    wire N__65988;
    wire N__65987;
    wire N__65984;
    wire N__65979;
    wire N__65976;
    wire N__65973;
    wire N__65970;
    wire N__65967;
    wire N__65964;
    wire N__65961;
    wire N__65958;
    wire N__65951;
    wire N__65944;
    wire N__65943;
    wire N__65936;
    wire N__65933;
    wire N__65928;
    wire N__65927;
    wire N__65926;
    wire N__65925;
    wire N__65924;
    wire N__65923;
    wire N__65920;
    wire N__65909;
    wire N__65904;
    wire N__65901;
    wire N__65898;
    wire N__65895;
    wire N__65894;
    wire N__65893;
    wire N__65892;
    wire N__65891;
    wire N__65890;
    wire N__65889;
    wire N__65886;
    wire N__65885;
    wire N__65884;
    wire N__65883;
    wire N__65882;
    wire N__65881;
    wire N__65880;
    wire N__65879;
    wire N__65876;
    wire N__65865;
    wire N__65858;
    wire N__65847;
    wire N__65838;
    wire N__65835;
    wire N__65832;
    wire N__65829;
    wire N__65828;
    wire N__65823;
    wire N__65820;
    wire N__65819;
    wire N__65816;
    wire N__65813;
    wire N__65810;
    wire N__65805;
    wire N__65804;
    wire N__65801;
    wire N__65798;
    wire N__65795;
    wire N__65794;
    wire N__65791;
    wire N__65788;
    wire N__65785;
    wire N__65782;
    wire N__65775;
    wire N__65774;
    wire N__65769;
    wire N__65766;
    wire N__65763;
    wire N__65760;
    wire N__65759;
    wire N__65758;
    wire N__65755;
    wire N__65750;
    wire N__65745;
    wire N__65744;
    wire N__65743;
    wire N__65740;
    wire N__65735;
    wire N__65730;
    wire N__65727;
    wire N__65724;
    wire N__65721;
    wire N__65718;
    wire N__65715;
    wire N__65714;
    wire N__65711;
    wire N__65708;
    wire N__65703;
    wire N__65702;
    wire N__65699;
    wire N__65696;
    wire N__65691;
    wire N__65688;
    wire N__65685;
    wire N__65682;
    wire N__65679;
    wire N__65676;
    wire N__65673;
    wire N__65672;
    wire N__65667;
    wire N__65664;
    wire N__65663;
    wire N__65658;
    wire N__65655;
    wire N__65654;
    wire N__65651;
    wire N__65648;
    wire N__65645;
    wire N__65640;
    wire N__65637;
    wire N__65634;
    wire N__65631;
    wire N__65628;
    wire N__65625;
    wire N__65622;
    wire N__65619;
    wire N__65618;
    wire N__65615;
    wire N__65612;
    wire N__65607;
    wire N__65606;
    wire N__65603;
    wire N__65600;
    wire N__65595;
    wire N__65592;
    wire N__65591;
    wire N__65588;
    wire N__65585;
    wire N__65580;
    wire N__65577;
    wire N__65576;
    wire N__65575;
    wire N__65572;
    wire N__65569;
    wire N__65566;
    wire N__65563;
    wire N__65556;
    wire N__65553;
    wire N__65552;
    wire N__65551;
    wire N__65548;
    wire N__65545;
    wire N__65542;
    wire N__65539;
    wire N__65532;
    wire N__65529;
    wire N__65526;
    wire N__65523;
    wire N__65520;
    wire N__65517;
    wire N__65514;
    wire N__65511;
    wire N__65510;
    wire N__65509;
    wire N__65508;
    wire N__65505;
    wire N__65502;
    wire N__65497;
    wire N__65494;
    wire N__65487;
    wire N__65486;
    wire N__65483;
    wire N__65480;
    wire N__65479;
    wire N__65476;
    wire N__65473;
    wire N__65470;
    wire N__65467;
    wire N__65462;
    wire N__65457;
    wire N__65456;
    wire N__65455;
    wire N__65454;
    wire N__65451;
    wire N__65450;
    wire N__65449;
    wire N__65446;
    wire N__65443;
    wire N__65440;
    wire N__65439;
    wire N__65438;
    wire N__65437;
    wire N__65436;
    wire N__65433;
    wire N__65432;
    wire N__65415;
    wire N__65412;
    wire N__65409;
    wire N__65408;
    wire N__65407;
    wire N__65404;
    wire N__65403;
    wire N__65402;
    wire N__65401;
    wire N__65400;
    wire N__65399;
    wire N__65398;
    wire N__65397;
    wire N__65396;
    wire N__65393;
    wire N__65390;
    wire N__65387;
    wire N__65372;
    wire N__65365;
    wire N__65362;
    wire N__65359;
    wire N__65356;
    wire N__65351;
    wire N__65348;
    wire N__65347;
    wire N__65344;
    wire N__65341;
    wire N__65340;
    wire N__65333;
    wire N__65330;
    wire N__65327;
    wire N__65324;
    wire N__65321;
    wire N__65318;
    wire N__65307;
    wire N__65306;
    wire N__65305;
    wire N__65304;
    wire N__65303;
    wire N__65300;
    wire N__65299;
    wire N__65298;
    wire N__65297;
    wire N__65296;
    wire N__65295;
    wire N__65292;
    wire N__65291;
    wire N__65290;
    wire N__65289;
    wire N__65288;
    wire N__65287;
    wire N__65286;
    wire N__65285;
    wire N__65284;
    wire N__65283;
    wire N__65280;
    wire N__65279;
    wire N__65278;
    wire N__65277;
    wire N__65274;
    wire N__65273;
    wire N__65272;
    wire N__65271;
    wire N__65268;
    wire N__65267;
    wire N__65266;
    wire N__65265;
    wire N__65264;
    wire N__65261;
    wire N__65258;
    wire N__65255;
    wire N__65252;
    wire N__65249;
    wire N__65248;
    wire N__65247;
    wire N__65244;
    wire N__65243;
    wire N__65240;
    wire N__65237;
    wire N__65234;
    wire N__65231;
    wire N__65228;
    wire N__65225;
    wire N__65224;
    wire N__65223;
    wire N__65222;
    wire N__65219;
    wire N__65218;
    wire N__65217;
    wire N__65214;
    wire N__65213;
    wire N__65210;
    wire N__65197;
    wire N__65194;
    wire N__65191;
    wire N__65190;
    wire N__65189;
    wire N__65188;
    wire N__65187;
    wire N__65184;
    wire N__65183;
    wire N__65182;
    wire N__65177;
    wire N__65174;
    wire N__65173;
    wire N__65172;
    wire N__65169;
    wire N__65168;
    wire N__65167;
    wire N__65164;
    wire N__65161;
    wire N__65156;
    wire N__65149;
    wire N__65142;
    wire N__65139;
    wire N__65134;
    wire N__65121;
    wire N__65108;
    wire N__65105;
    wire N__65100;
    wire N__65099;
    wire N__65096;
    wire N__65093;
    wire N__65082;
    wire N__65081;
    wire N__65078;
    wire N__65069;
    wire N__65062;
    wire N__65055;
    wire N__65054;
    wire N__65051;
    wire N__65048;
    wire N__65045;
    wire N__65036;
    wire N__65029;
    wire N__65026;
    wire N__65023;
    wire N__65014;
    wire N__65011;
    wire N__65008;
    wire N__65001;
    wire N__64998;
    wire N__64991;
    wire N__64988;
    wire N__64985;
    wire N__64976;
    wire N__64971;
    wire N__64968;
    wire N__64965;
    wire N__64962;
    wire N__64959;
    wire N__64956;
    wire N__64953;
    wire N__64950;
    wire N__64947;
    wire N__64946;
    wire N__64945;
    wire N__64942;
    wire N__64939;
    wire N__64936;
    wire N__64931;
    wire N__64926;
    wire N__64923;
    wire N__64920;
    wire N__64917;
    wire N__64916;
    wire N__64915;
    wire N__64912;
    wire N__64909;
    wire N__64906;
    wire N__64901;
    wire N__64896;
    wire N__64893;
    wire N__64890;
    wire N__64889;
    wire N__64886;
    wire N__64883;
    wire N__64882;
    wire N__64879;
    wire N__64876;
    wire N__64873;
    wire N__64868;
    wire N__64863;
    wire N__64860;
    wire N__64857;
    wire N__64854;
    wire N__64851;
    wire N__64850;
    wire N__64847;
    wire N__64844;
    wire N__64843;
    wire N__64838;
    wire N__64835;
    wire N__64832;
    wire N__64827;
    wire N__64824;
    wire N__64823;
    wire N__64822;
    wire N__64819;
    wire N__64816;
    wire N__64813;
    wire N__64806;
    wire N__64803;
    wire N__64802;
    wire N__64801;
    wire N__64798;
    wire N__64795;
    wire N__64792;
    wire N__64785;
    wire N__64782;
    wire N__64781;
    wire N__64780;
    wire N__64777;
    wire N__64774;
    wire N__64771;
    wire N__64768;
    wire N__64761;
    wire N__64758;
    wire N__64757;
    wire N__64754;
    wire N__64753;
    wire N__64750;
    wire N__64747;
    wire N__64744;
    wire N__64737;
    wire N__64734;
    wire N__64731;
    wire N__64728;
    wire N__64725;
    wire N__64722;
    wire N__64719;
    wire N__64716;
    wire N__64713;
    wire N__64710;
    wire N__64707;
    wire N__64704;
    wire N__64701;
    wire N__64698;
    wire N__64695;
    wire N__64692;
    wire N__64689;
    wire N__64686;
    wire N__64683;
    wire N__64680;
    wire N__64677;
    wire N__64674;
    wire N__64673;
    wire N__64670;
    wire N__64669;
    wire N__64666;
    wire N__64663;
    wire N__64658;
    wire N__64655;
    wire N__64654;
    wire N__64651;
    wire N__64648;
    wire N__64645;
    wire N__64642;
    wire N__64635;
    wire N__64634;
    wire N__64631;
    wire N__64628;
    wire N__64625;
    wire N__64622;
    wire N__64619;
    wire N__64618;
    wire N__64615;
    wire N__64612;
    wire N__64609;
    wire N__64602;
    wire N__64601;
    wire N__64600;
    wire N__64599;
    wire N__64598;
    wire N__64597;
    wire N__64596;
    wire N__64595;
    wire N__64592;
    wire N__64591;
    wire N__64590;
    wire N__64587;
    wire N__64586;
    wire N__64585;
    wire N__64584;
    wire N__64583;
    wire N__64582;
    wire N__64577;
    wire N__64576;
    wire N__64573;
    wire N__64570;
    wire N__64565;
    wire N__64562;
    wire N__64557;
    wire N__64552;
    wire N__64549;
    wire N__64548;
    wire N__64547;
    wire N__64546;
    wire N__64543;
    wire N__64538;
    wire N__64535;
    wire N__64532;
    wire N__64527;
    wire N__64524;
    wire N__64521;
    wire N__64520;
    wire N__64517;
    wire N__64514;
    wire N__64505;
    wire N__64504;
    wire N__64495;
    wire N__64488;
    wire N__64487;
    wire N__64484;
    wire N__64479;
    wire N__64476;
    wire N__64473;
    wire N__64468;
    wire N__64463;
    wire N__64458;
    wire N__64449;
    wire N__64448;
    wire N__64445;
    wire N__64444;
    wire N__64443;
    wire N__64442;
    wire N__64441;
    wire N__64438;
    wire N__64437;
    wire N__64436;
    wire N__64435;
    wire N__64432;
    wire N__64431;
    wire N__64428;
    wire N__64423;
    wire N__64420;
    wire N__64411;
    wire N__64408;
    wire N__64405;
    wire N__64402;
    wire N__64399;
    wire N__64398;
    wire N__64397;
    wire N__64396;
    wire N__64395;
    wire N__64392;
    wire N__64391;
    wire N__64390;
    wire N__64389;
    wire N__64388;
    wire N__64377;
    wire N__64374;
    wire N__64371;
    wire N__64366;
    wire N__64363;
    wire N__64358;
    wire N__64353;
    wire N__64350;
    wire N__64347;
    wire N__64332;
    wire N__64329;
    wire N__64326;
    wire N__64323;
    wire N__64320;
    wire N__64317;
    wire N__64314;
    wire N__64311;
    wire N__64308;
    wire N__64305;
    wire N__64304;
    wire N__64303;
    wire N__64302;
    wire N__64299;
    wire N__64296;
    wire N__64295;
    wire N__64294;
    wire N__64293;
    wire N__64292;
    wire N__64291;
    wire N__64290;
    wire N__64289;
    wire N__64288;
    wire N__64287;
    wire N__64286;
    wire N__64281;
    wire N__64278;
    wire N__64275;
    wire N__64274;
    wire N__64273;
    wire N__64272;
    wire N__64271;
    wire N__64270;
    wire N__64269;
    wire N__64268;
    wire N__64267;
    wire N__64266;
    wire N__64265;
    wire N__64264;
    wire N__64263;
    wire N__64262;
    wire N__64261;
    wire N__64260;
    wire N__64259;
    wire N__64258;
    wire N__64257;
    wire N__64256;
    wire N__64255;
    wire N__64248;
    wire N__64243;
    wire N__64240;
    wire N__64239;
    wire N__64234;
    wire N__64233;
    wire N__64232;
    wire N__64231;
    wire N__64230;
    wire N__64225;
    wire N__64218;
    wire N__64211;
    wire N__64206;
    wire N__64201;
    wire N__64192;
    wire N__64185;
    wire N__64176;
    wire N__64173;
    wire N__64172;
    wire N__64169;
    wire N__64168;
    wire N__64167;
    wire N__64166;
    wire N__64165;
    wire N__64164;
    wire N__64161;
    wire N__64158;
    wire N__64155;
    wire N__64152;
    wire N__64149;
    wire N__64148;
    wire N__64147;
    wire N__64146;
    wire N__64137;
    wire N__64128;
    wire N__64123;
    wire N__64116;
    wire N__64113;
    wire N__64110;
    wire N__64105;
    wire N__64104;
    wire N__64103;
    wire N__64102;
    wire N__64101;
    wire N__64094;
    wire N__64091;
    wire N__64082;
    wire N__64079;
    wire N__64074;
    wire N__64067;
    wire N__64064;
    wire N__64057;
    wire N__64050;
    wire N__64047;
    wire N__64026;
    wire N__64023;
    wire N__64020;
    wire N__64019;
    wire N__64016;
    wire N__64015;
    wire N__64012;
    wire N__64009;
    wire N__64006;
    wire N__63999;
    wire N__63996;
    wire N__63993;
    wire N__63992;
    wire N__63989;
    wire N__63988;
    wire N__63985;
    wire N__63982;
    wire N__63979;
    wire N__63972;
    wire N__63969;
    wire N__63966;
    wire N__63963;
    wire N__63960;
    wire N__63957;
    wire N__63954;
    wire N__63951;
    wire N__63948;
    wire N__63945;
    wire N__63942;
    wire N__63939;
    wire N__63936;
    wire N__63935;
    wire N__63932;
    wire N__63929;
    wire N__63928;
    wire N__63925;
    wire N__63922;
    wire N__63919;
    wire N__63912;
    wire N__63909;
    wire N__63908;
    wire N__63907;
    wire N__63904;
    wire N__63903;
    wire N__63900;
    wire N__63897;
    wire N__63894;
    wire N__63891;
    wire N__63888;
    wire N__63885;
    wire N__63882;
    wire N__63879;
    wire N__63874;
    wire N__63869;
    wire N__63864;
    wire N__63861;
    wire N__63860;
    wire N__63859;
    wire N__63858;
    wire N__63857;
    wire N__63854;
    wire N__63851;
    wire N__63848;
    wire N__63847;
    wire N__63844;
    wire N__63841;
    wire N__63836;
    wire N__63833;
    wire N__63830;
    wire N__63827;
    wire N__63824;
    wire N__63819;
    wire N__63816;
    wire N__63807;
    wire N__63806;
    wire N__63805;
    wire N__63804;
    wire N__63803;
    wire N__63798;
    wire N__63797;
    wire N__63796;
    wire N__63795;
    wire N__63794;
    wire N__63793;
    wire N__63790;
    wire N__63789;
    wire N__63788;
    wire N__63783;
    wire N__63780;
    wire N__63779;
    wire N__63776;
    wire N__63771;
    wire N__63766;
    wire N__63763;
    wire N__63758;
    wire N__63757;
    wire N__63756;
    wire N__63753;
    wire N__63750;
    wire N__63747;
    wire N__63742;
    wire N__63741;
    wire N__63738;
    wire N__63733;
    wire N__63730;
    wire N__63727;
    wire N__63722;
    wire N__63717;
    wire N__63714;
    wire N__63709;
    wire N__63706;
    wire N__63693;
    wire N__63690;
    wire N__63689;
    wire N__63686;
    wire N__63683;
    wire N__63682;
    wire N__63679;
    wire N__63676;
    wire N__63675;
    wire N__63672;
    wire N__63669;
    wire N__63666;
    wire N__63663;
    wire N__63660;
    wire N__63657;
    wire N__63652;
    wire N__63645;
    wire N__63644;
    wire N__63641;
    wire N__63638;
    wire N__63635;
    wire N__63632;
    wire N__63629;
    wire N__63626;
    wire N__63621;
    wire N__63618;
    wire N__63617;
    wire N__63614;
    wire N__63613;
    wire N__63610;
    wire N__63607;
    wire N__63602;
    wire N__63597;
    wire N__63594;
    wire N__63593;
    wire N__63592;
    wire N__63591;
    wire N__63590;
    wire N__63589;
    wire N__63588;
    wire N__63585;
    wire N__63584;
    wire N__63581;
    wire N__63576;
    wire N__63573;
    wire N__63568;
    wire N__63565;
    wire N__63562;
    wire N__63559;
    wire N__63556;
    wire N__63555;
    wire N__63552;
    wire N__63549;
    wire N__63546;
    wire N__63545;
    wire N__63544;
    wire N__63539;
    wire N__63536;
    wire N__63533;
    wire N__63526;
    wire N__63521;
    wire N__63510;
    wire N__63507;
    wire N__63504;
    wire N__63501;
    wire N__63500;
    wire N__63499;
    wire N__63498;
    wire N__63495;
    wire N__63492;
    wire N__63489;
    wire N__63486;
    wire N__63483;
    wire N__63478;
    wire N__63475;
    wire N__63470;
    wire N__63465;
    wire N__63462;
    wire N__63461;
    wire N__63460;
    wire N__63459;
    wire N__63458;
    wire N__63457;
    wire N__63456;
    wire N__63451;
    wire N__63450;
    wire N__63449;
    wire N__63442;
    wire N__63441;
    wire N__63440;
    wire N__63439;
    wire N__63438;
    wire N__63435;
    wire N__63432;
    wire N__63431;
    wire N__63430;
    wire N__63427;
    wire N__63424;
    wire N__63423;
    wire N__63422;
    wire N__63419;
    wire N__63416;
    wire N__63407;
    wire N__63406;
    wire N__63405;
    wire N__63404;
    wire N__63403;
    wire N__63400;
    wire N__63397;
    wire N__63392;
    wire N__63391;
    wire N__63390;
    wire N__63389;
    wire N__63388;
    wire N__63385;
    wire N__63382;
    wire N__63381;
    wire N__63376;
    wire N__63371;
    wire N__63368;
    wire N__63363;
    wire N__63360;
    wire N__63359;
    wire N__63356;
    wire N__63355;
    wire N__63354;
    wire N__63349;
    wire N__63346;
    wire N__63341;
    wire N__63338;
    wire N__63335;
    wire N__63330;
    wire N__63327;
    wire N__63320;
    wire N__63317;
    wire N__63306;
    wire N__63299;
    wire N__63282;
    wire N__63279;
    wire N__63276;
    wire N__63273;
    wire N__63270;
    wire N__63267;
    wire N__63264;
    wire N__63261;
    wire N__63258;
    wire N__63255;
    wire N__63252;
    wire N__63249;
    wire N__63246;
    wire N__63243;
    wire N__63240;
    wire N__63237;
    wire N__63236;
    wire N__63235;
    wire N__63232;
    wire N__63231;
    wire N__63228;
    wire N__63225;
    wire N__63222;
    wire N__63217;
    wire N__63214;
    wire N__63209;
    wire N__63204;
    wire N__63201;
    wire N__63198;
    wire N__63195;
    wire N__63192;
    wire N__63189;
    wire N__63186;
    wire N__63183;
    wire N__63180;
    wire N__63177;
    wire N__63174;
    wire N__63171;
    wire N__63168;
    wire N__63165;
    wire N__63162;
    wire N__63161;
    wire N__63158;
    wire N__63155;
    wire N__63150;
    wire N__63149;
    wire N__63148;
    wire N__63145;
    wire N__63142;
    wire N__63141;
    wire N__63138;
    wire N__63135;
    wire N__63130;
    wire N__63123;
    wire N__63120;
    wire N__63119;
    wire N__63116;
    wire N__63113;
    wire N__63110;
    wire N__63105;
    wire N__63102;
    wire N__63101;
    wire N__63098;
    wire N__63097;
    wire N__63096;
    wire N__63093;
    wire N__63090;
    wire N__63085;
    wire N__63078;
    wire N__63077;
    wire N__63076;
    wire N__63073;
    wire N__63068;
    wire N__63063;
    wire N__63060;
    wire N__63057;
    wire N__63054;
    wire N__63051;
    wire N__63048;
    wire N__63045;
    wire N__63042;
    wire N__63039;
    wire N__63036;
    wire N__63033;
    wire N__63030;
    wire N__63027;
    wire N__63024;
    wire N__63023;
    wire N__63020;
    wire N__63017;
    wire N__63012;
    wire N__63009;
    wire N__63006;
    wire N__63003;
    wire N__63000;
    wire N__62997;
    wire N__62996;
    wire N__62993;
    wire N__62990;
    wire N__62987;
    wire N__62986;
    wire N__62983;
    wire N__62980;
    wire N__62977;
    wire N__62976;
    wire N__62973;
    wire N__62970;
    wire N__62969;
    wire N__62968;
    wire N__62965;
    wire N__62962;
    wire N__62959;
    wire N__62956;
    wire N__62951;
    wire N__62948;
    wire N__62943;
    wire N__62940;
    wire N__62931;
    wire N__62928;
    wire N__62925;
    wire N__62924;
    wire N__62921;
    wire N__62918;
    wire N__62913;
    wire N__62910;
    wire N__62907;
    wire N__62904;
    wire N__62901;
    wire N__62900;
    wire N__62899;
    wire N__62898;
    wire N__62895;
    wire N__62888;
    wire N__62883;
    wire N__62880;
    wire N__62879;
    wire N__62876;
    wire N__62873;
    wire N__62870;
    wire N__62867;
    wire N__62862;
    wire N__62859;
    wire N__62858;
    wire N__62855;
    wire N__62852;
    wire N__62847;
    wire N__62844;
    wire N__62841;
    wire N__62838;
    wire N__62835;
    wire N__62832;
    wire N__62829;
    wire N__62828;
    wire N__62827;
    wire N__62824;
    wire N__62823;
    wire N__62822;
    wire N__62817;
    wire N__62814;
    wire N__62809;
    wire N__62806;
    wire N__62801;
    wire N__62798;
    wire N__62795;
    wire N__62790;
    wire N__62787;
    wire N__62786;
    wire N__62783;
    wire N__62782;
    wire N__62779;
    wire N__62776;
    wire N__62773;
    wire N__62766;
    wire N__62763;
    wire N__62760;
    wire N__62757;
    wire N__62754;
    wire N__62751;
    wire N__62748;
    wire N__62745;
    wire N__62742;
    wire N__62739;
    wire N__62736;
    wire N__62733;
    wire N__62730;
    wire N__62727;
    wire N__62724;
    wire N__62721;
    wire N__62718;
    wire N__62715;
    wire N__62712;
    wire N__62709;
    wire N__62706;
    wire N__62703;
    wire N__62700;
    wire N__62697;
    wire N__62694;
    wire N__62691;
    wire N__62688;
    wire N__62685;
    wire N__62682;
    wire N__62679;
    wire N__62676;
    wire N__62673;
    wire N__62670;
    wire N__62667;
    wire N__62664;
    wire N__62661;
    wire N__62658;
    wire N__62655;
    wire N__62652;
    wire N__62649;
    wire N__62646;
    wire N__62643;
    wire N__62640;
    wire N__62637;
    wire N__62634;
    wire N__62631;
    wire N__62628;
    wire N__62625;
    wire N__62622;
    wire N__62619;
    wire N__62616;
    wire N__62613;
    wire N__62610;
    wire N__62607;
    wire N__62604;
    wire N__62603;
    wire N__62600;
    wire N__62597;
    wire N__62592;
    wire N__62589;
    wire N__62586;
    wire N__62583;
    wire N__62580;
    wire N__62577;
    wire N__62574;
    wire N__62571;
    wire N__62568;
    wire N__62567;
    wire N__62566;
    wire N__62561;
    wire N__62558;
    wire N__62555;
    wire N__62554;
    wire N__62553;
    wire N__62552;
    wire N__62547;
    wire N__62540;
    wire N__62535;
    wire N__62534;
    wire N__62533;
    wire N__62532;
    wire N__62529;
    wire N__62526;
    wire N__62521;
    wire N__62514;
    wire N__62511;
    wire N__62510;
    wire N__62507;
    wire N__62504;
    wire N__62499;
    wire N__62496;
    wire N__62495;
    wire N__62492;
    wire N__62489;
    wire N__62486;
    wire N__62483;
    wire N__62478;
    wire N__62477;
    wire N__62474;
    wire N__62471;
    wire N__62466;
    wire N__62463;
    wire N__62460;
    wire N__62457;
    wire N__62456;
    wire N__62455;
    wire N__62454;
    wire N__62451;
    wire N__62446;
    wire N__62443;
    wire N__62436;
    wire N__62433;
    wire N__62432;
    wire N__62431;
    wire N__62430;
    wire N__62429;
    wire N__62426;
    wire N__62423;
    wire N__62420;
    wire N__62415;
    wire N__62406;
    wire N__62403;
    wire N__62400;
    wire N__62399;
    wire N__62396;
    wire N__62393;
    wire N__62388;
    wire N__62387;
    wire N__62382;
    wire N__62379;
    wire N__62378;
    wire N__62375;
    wire N__62372;
    wire N__62367;
    wire N__62364;
    wire N__62361;
    wire N__62358;
    wire N__62355;
    wire N__62352;
    wire N__62351;
    wire N__62350;
    wire N__62347;
    wire N__62342;
    wire N__62337;
    wire N__62334;
    wire N__62331;
    wire N__62328;
    wire N__62325;
    wire N__62322;
    wire N__62319;
    wire N__62318;
    wire N__62317;
    wire N__62314;
    wire N__62311;
    wire N__62308;
    wire N__62307;
    wire N__62304;
    wire N__62301;
    wire N__62296;
    wire N__62289;
    wire N__62286;
    wire N__62283;
    wire N__62282;
    wire N__62281;
    wire N__62278;
    wire N__62275;
    wire N__62272;
    wire N__62265;
    wire N__62264;
    wire N__62263;
    wire N__62260;
    wire N__62257;
    wire N__62254;
    wire N__62247;
    wire N__62246;
    wire N__62243;
    wire N__62240;
    wire N__62235;
    wire N__62232;
    wire N__62229;
    wire N__62226;
    wire N__62225;
    wire N__62222;
    wire N__62219;
    wire N__62214;
    wire N__62211;
    wire N__62208;
    wire N__62207;
    wire N__62206;
    wire N__62205;
    wire N__62204;
    wire N__62201;
    wire N__62198;
    wire N__62197;
    wire N__62194;
    wire N__62191;
    wire N__62190;
    wire N__62187;
    wire N__62186;
    wire N__62185;
    wire N__62182;
    wire N__62171;
    wire N__62166;
    wire N__62163;
    wire N__62160;
    wire N__62157;
    wire N__62154;
    wire N__62145;
    wire N__62142;
    wire N__62141;
    wire N__62138;
    wire N__62137;
    wire N__62136;
    wire N__62135;
    wire N__62134;
    wire N__62133;
    wire N__62132;
    wire N__62131;
    wire N__62130;
    wire N__62127;
    wire N__62124;
    wire N__62113;
    wire N__62108;
    wire N__62103;
    wire N__62100;
    wire N__62097;
    wire N__62094;
    wire N__62085;
    wire N__62084;
    wire N__62081;
    wire N__62078;
    wire N__62075;
    wire N__62074;
    wire N__62073;
    wire N__62072;
    wire N__62071;
    wire N__62070;
    wire N__62065;
    wire N__62054;
    wire N__62053;
    wire N__62048;
    wire N__62047;
    wire N__62046;
    wire N__62045;
    wire N__62042;
    wire N__62039;
    wire N__62032;
    wire N__62025;
    wire N__62022;
    wire N__62019;
    wire N__62016;
    wire N__62013;
    wire N__62010;
    wire N__62007;
    wire N__62006;
    wire N__62005;
    wire N__62002;
    wire N__61997;
    wire N__61992;
    wire N__61989;
    wire N__61986;
    wire N__61983;
    wire N__61980;
    wire N__61977;
    wire N__61974;
    wire N__61971;
    wire N__61968;
    wire N__61965;
    wire N__61962;
    wire N__61959;
    wire N__61956;
    wire N__61953;
    wire N__61950;
    wire N__61947;
    wire N__61944;
    wire N__61941;
    wire N__61938;
    wire N__61935;
    wire N__61934;
    wire N__61931;
    wire N__61928;
    wire N__61925;
    wire N__61920;
    wire N__61917;
    wire N__61916;
    wire N__61913;
    wire N__61910;
    wire N__61907;
    wire N__61904;
    wire N__61901;
    wire N__61898;
    wire N__61893;
    wire N__61892;
    wire N__61891;
    wire N__61890;
    wire N__61889;
    wire N__61884;
    wire N__61879;
    wire N__61876;
    wire N__61869;
    wire N__61866;
    wire N__61863;
    wire N__61860;
    wire N__61857;
    wire N__61854;
    wire N__61853;
    wire N__61852;
    wire N__61851;
    wire N__61850;
    wire N__61849;
    wire N__61848;
    wire N__61841;
    wire N__61840;
    wire N__61837;
    wire N__61836;
    wire N__61829;
    wire N__61826;
    wire N__61823;
    wire N__61818;
    wire N__61809;
    wire N__61808;
    wire N__61805;
    wire N__61802;
    wire N__61799;
    wire N__61796;
    wire N__61795;
    wire N__61790;
    wire N__61787;
    wire N__61784;
    wire N__61779;
    wire N__61776;
    wire N__61773;
    wire N__61770;
    wire N__61767;
    wire N__61766;
    wire N__61763;
    wire N__61762;
    wire N__61759;
    wire N__61756;
    wire N__61753;
    wire N__61750;
    wire N__61747;
    wire N__61744;
    wire N__61741;
    wire N__61738;
    wire N__61731;
    wire N__61730;
    wire N__61727;
    wire N__61724;
    wire N__61723;
    wire N__61720;
    wire N__61717;
    wire N__61714;
    wire N__61711;
    wire N__61708;
    wire N__61701;
    wire N__61698;
    wire N__61695;
    wire N__61694;
    wire N__61691;
    wire N__61690;
    wire N__61689;
    wire N__61686;
    wire N__61683;
    wire N__61680;
    wire N__61675;
    wire N__61672;
    wire N__61669;
    wire N__61666;
    wire N__61663;
    wire N__61660;
    wire N__61657;
    wire N__61650;
    wire N__61647;
    wire N__61644;
    wire N__61641;
    wire N__61640;
    wire N__61639;
    wire N__61638;
    wire N__61637;
    wire N__61634;
    wire N__61633;
    wire N__61632;
    wire N__61631;
    wire N__61630;
    wire N__61629;
    wire N__61628;
    wire N__61627;
    wire N__61626;
    wire N__61625;
    wire N__61620;
    wire N__61619;
    wire N__61618;
    wire N__61615;
    wire N__61612;
    wire N__61605;
    wire N__61604;
    wire N__61601;
    wire N__61596;
    wire N__61593;
    wire N__61590;
    wire N__61585;
    wire N__61582;
    wire N__61581;
    wire N__61580;
    wire N__61575;
    wire N__61572;
    wire N__61567;
    wire N__61566;
    wire N__61565;
    wire N__61562;
    wire N__61559;
    wire N__61556;
    wire N__61553;
    wire N__61550;
    wire N__61547;
    wire N__61544;
    wire N__61539;
    wire N__61536;
    wire N__61531;
    wire N__61528;
    wire N__61525;
    wire N__61518;
    wire N__61509;
    wire N__61504;
    wire N__61501;
    wire N__61488;
    wire N__61487;
    wire N__61486;
    wire N__61483;
    wire N__61480;
    wire N__61477;
    wire N__61474;
    wire N__61471;
    wire N__61468;
    wire N__61463;
    wire N__61458;
    wire N__61457;
    wire N__61456;
    wire N__61453;
    wire N__61452;
    wire N__61451;
    wire N__61450;
    wire N__61449;
    wire N__61448;
    wire N__61447;
    wire N__61444;
    wire N__61443;
    wire N__61440;
    wire N__61437;
    wire N__61434;
    wire N__61431;
    wire N__61430;
    wire N__61427;
    wire N__61424;
    wire N__61421;
    wire N__61420;
    wire N__61419;
    wire N__61418;
    wire N__61417;
    wire N__61414;
    wire N__61407;
    wire N__61404;
    wire N__61397;
    wire N__61396;
    wire N__61395;
    wire N__61394;
    wire N__61389;
    wire N__61384;
    wire N__61379;
    wire N__61376;
    wire N__61373;
    wire N__61370;
    wire N__61365;
    wire N__61362;
    wire N__61357;
    wire N__61352;
    wire N__61349;
    wire N__61346;
    wire N__61341;
    wire N__61338;
    wire N__61335;
    wire N__61332;
    wire N__61329;
    wire N__61326;
    wire N__61319;
    wire N__61308;
    wire N__61307;
    wire N__61304;
    wire N__61303;
    wire N__61300;
    wire N__61297;
    wire N__61294;
    wire N__61291;
    wire N__61286;
    wire N__61281;
    wire N__61278;
    wire N__61275;
    wire N__61272;
    wire N__61269;
    wire N__61266;
    wire N__61263;
    wire N__61260;
    wire N__61257;
    wire N__61254;
    wire N__61251;
    wire N__61248;
    wire N__61245;
    wire N__61242;
    wire N__61239;
    wire N__61238;
    wire N__61233;
    wire N__61230;
    wire N__61227;
    wire N__61224;
    wire N__61221;
    wire N__61218;
    wire N__61217;
    wire N__61214;
    wire N__61211;
    wire N__61208;
    wire N__61205;
    wire N__61204;
    wire N__61203;
    wire N__61202;
    wire N__61199;
    wire N__61196;
    wire N__61193;
    wire N__61188;
    wire N__61179;
    wire N__61178;
    wire N__61173;
    wire N__61170;
    wire N__61167;
    wire N__61164;
    wire N__61163;
    wire N__61162;
    wire N__61161;
    wire N__61156;
    wire N__61153;
    wire N__61150;
    wire N__61147;
    wire N__61144;
    wire N__61141;
    wire N__61138;
    wire N__61137;
    wire N__61136;
    wire N__61135;
    wire N__61130;
    wire N__61127;
    wire N__61124;
    wire N__61119;
    wire N__61110;
    wire N__61109;
    wire N__61106;
    wire N__61105;
    wire N__61102;
    wire N__61099;
    wire N__61096;
    wire N__61093;
    wire N__61086;
    wire N__61083;
    wire N__61080;
    wire N__61077;
    wire N__61074;
    wire N__61071;
    wire N__61068;
    wire N__61065;
    wire N__61064;
    wire N__61061;
    wire N__61058;
    wire N__61057;
    wire N__61056;
    wire N__61055;
    wire N__61054;
    wire N__61053;
    wire N__61052;
    wire N__61047;
    wire N__61044;
    wire N__61043;
    wire N__61042;
    wire N__61041;
    wire N__61034;
    wire N__61029;
    wire N__61026;
    wire N__61023;
    wire N__61020;
    wire N__61019;
    wire N__61016;
    wire N__61015;
    wire N__61014;
    wire N__61011;
    wire N__61008;
    wire N__61001;
    wire N__60996;
    wire N__60991;
    wire N__60988;
    wire N__60987;
    wire N__60986;
    wire N__60985;
    wire N__60978;
    wire N__60975;
    wire N__60972;
    wire N__60969;
    wire N__60964;
    wire N__60961;
    wire N__60958;
    wire N__60953;
    wire N__60942;
    wire N__60941;
    wire N__60940;
    wire N__60939;
    wire N__60938;
    wire N__60935;
    wire N__60934;
    wire N__60933;
    wire N__60932;
    wire N__60931;
    wire N__60926;
    wire N__60925;
    wire N__60924;
    wire N__60923;
    wire N__60918;
    wire N__60909;
    wire N__60908;
    wire N__60907;
    wire N__60906;
    wire N__60905;
    wire N__60904;
    wire N__60901;
    wire N__60898;
    wire N__60897;
    wire N__60894;
    wire N__60891;
    wire N__60888;
    wire N__60885;
    wire N__60882;
    wire N__60881;
    wire N__60880;
    wire N__60879;
    wire N__60876;
    wire N__60869;
    wire N__60866;
    wire N__60861;
    wire N__60860;
    wire N__60859;
    wire N__60856;
    wire N__60853;
    wire N__60848;
    wire N__60843;
    wire N__60836;
    wire N__60833;
    wire N__60830;
    wire N__60825;
    wire N__60820;
    wire N__60801;
    wire N__60798;
    wire N__60795;
    wire N__60794;
    wire N__60791;
    wire N__60790;
    wire N__60787;
    wire N__60784;
    wire N__60781;
    wire N__60778;
    wire N__60775;
    wire N__60768;
    wire N__60765;
    wire N__60762;
    wire N__60759;
    wire N__60758;
    wire N__60757;
    wire N__60754;
    wire N__60751;
    wire N__60748;
    wire N__60745;
    wire N__60742;
    wire N__60739;
    wire N__60736;
    wire N__60733;
    wire N__60728;
    wire N__60723;
    wire N__60720;
    wire N__60717;
    wire N__60716;
    wire N__60713;
    wire N__60710;
    wire N__60707;
    wire N__60704;
    wire N__60703;
    wire N__60700;
    wire N__60697;
    wire N__60694;
    wire N__60689;
    wire N__60684;
    wire N__60683;
    wire N__60682;
    wire N__60679;
    wire N__60676;
    wire N__60673;
    wire N__60670;
    wire N__60667;
    wire N__60664;
    wire N__60661;
    wire N__60658;
    wire N__60651;
    wire N__60648;
    wire N__60645;
    wire N__60642;
    wire N__60639;
    wire N__60636;
    wire N__60633;
    wire N__60630;
    wire N__60627;
    wire N__60624;
    wire N__60621;
    wire N__60618;
    wire N__60615;
    wire N__60612;
    wire N__60609;
    wire N__60608;
    wire N__60605;
    wire N__60602;
    wire N__60601;
    wire N__60598;
    wire N__60595;
    wire N__60592;
    wire N__60585;
    wire N__60582;
    wire N__60579;
    wire N__60578;
    wire N__60577;
    wire N__60576;
    wire N__60573;
    wire N__60570;
    wire N__60567;
    wire N__60564;
    wire N__60561;
    wire N__60556;
    wire N__60553;
    wire N__60548;
    wire N__60543;
    wire N__60540;
    wire N__60537;
    wire N__60534;
    wire N__60531;
    wire N__60528;
    wire N__60525;
    wire N__60522;
    wire N__60519;
    wire N__60516;
    wire N__60513;
    wire N__60510;
    wire N__60507;
    wire N__60504;
    wire N__60501;
    wire N__60498;
    wire N__60495;
    wire N__60492;
    wire N__60489;
    wire N__60486;
    wire N__60483;
    wire N__60480;
    wire N__60477;
    wire N__60474;
    wire N__60471;
    wire N__60468;
    wire N__60465;
    wire N__60462;
    wire N__60459;
    wire N__60456;
    wire N__60455;
    wire N__60452;
    wire N__60449;
    wire N__60444;
    wire N__60441;
    wire N__60438;
    wire N__60435;
    wire N__60432;
    wire N__60429;
    wire N__60426;
    wire N__60423;
    wire N__60420;
    wire N__60417;
    wire N__60414;
    wire N__60411;
    wire N__60408;
    wire N__60405;
    wire N__60402;
    wire N__60399;
    wire N__60396;
    wire N__60393;
    wire N__60390;
    wire N__60387;
    wire N__60384;
    wire N__60381;
    wire N__60378;
    wire N__60375;
    wire N__60372;
    wire N__60371;
    wire N__60368;
    wire N__60367;
    wire N__60364;
    wire N__60361;
    wire N__60358;
    wire N__60355;
    wire N__60350;
    wire N__60345;
    wire N__60342;
    wire N__60339;
    wire N__60336;
    wire N__60333;
    wire N__60330;
    wire N__60327;
    wire N__60324;
    wire N__60321;
    wire N__60318;
    wire N__60315;
    wire N__60312;
    wire N__60309;
    wire N__60306;
    wire N__60303;
    wire N__60300;
    wire N__60299;
    wire N__60296;
    wire N__60293;
    wire N__60292;
    wire N__60287;
    wire N__60284;
    wire N__60281;
    wire N__60276;
    wire N__60273;
    wire N__60270;
    wire N__60267;
    wire N__60264;
    wire N__60261;
    wire N__60258;
    wire N__60255;
    wire N__60252;
    wire N__60249;
    wire N__60246;
    wire N__60243;
    wire N__60240;
    wire N__60239;
    wire N__60236;
    wire N__60235;
    wire N__60232;
    wire N__60231;
    wire N__60228;
    wire N__60223;
    wire N__60220;
    wire N__60215;
    wire N__60210;
    wire N__60207;
    wire N__60204;
    wire N__60203;
    wire N__60198;
    wire N__60197;
    wire N__60196;
    wire N__60195;
    wire N__60192;
    wire N__60189;
    wire N__60186;
    wire N__60185;
    wire N__60184;
    wire N__60181;
    wire N__60178;
    wire N__60175;
    wire N__60172;
    wire N__60169;
    wire N__60166;
    wire N__60165;
    wire N__60162;
    wire N__60157;
    wire N__60154;
    wire N__60151;
    wire N__60146;
    wire N__60141;
    wire N__60136;
    wire N__60129;
    wire N__60128;
    wire N__60125;
    wire N__60122;
    wire N__60121;
    wire N__60120;
    wire N__60119;
    wire N__60118;
    wire N__60117;
    wire N__60116;
    wire N__60115;
    wire N__60114;
    wire N__60113;
    wire N__60112;
    wire N__60109;
    wire N__60094;
    wire N__60093;
    wire N__60090;
    wire N__60087;
    wire N__60082;
    wire N__60081;
    wire N__60076;
    wire N__60073;
    wire N__60070;
    wire N__60067;
    wire N__60064;
    wire N__60061;
    wire N__60060;
    wire N__60057;
    wire N__60054;
    wire N__60051;
    wire N__60048;
    wire N__60045;
    wire N__60042;
    wire N__60039;
    wire N__60036;
    wire N__60033;
    wire N__60024;
    wire N__60019;
    wire N__60014;
    wire N__60009;
    wire N__60006;
    wire N__60005;
    wire N__60002;
    wire N__59999;
    wire N__59996;
    wire N__59993;
    wire N__59990;
    wire N__59987;
    wire N__59984;
    wire N__59981;
    wire N__59978;
    wire N__59973;
    wire N__59970;
    wire N__59967;
    wire N__59964;
    wire N__59961;
    wire N__59958;
    wire N__59955;
    wire N__59954;
    wire N__59953;
    wire N__59952;
    wire N__59951;
    wire N__59950;
    wire N__59949;
    wire N__59946;
    wire N__59941;
    wire N__59936;
    wire N__59933;
    wire N__59930;
    wire N__59925;
    wire N__59922;
    wire N__59921;
    wire N__59920;
    wire N__59917;
    wire N__59916;
    wire N__59909;
    wire N__59908;
    wire N__59907;
    wire N__59904;
    wire N__59901;
    wire N__59898;
    wire N__59895;
    wire N__59892;
    wire N__59887;
    wire N__59874;
    wire N__59871;
    wire N__59868;
    wire N__59865;
    wire N__59864;
    wire N__59863;
    wire N__59860;
    wire N__59859;
    wire N__59856;
    wire N__59853;
    wire N__59850;
    wire N__59849;
    wire N__59848;
    wire N__59845;
    wire N__59844;
    wire N__59839;
    wire N__59836;
    wire N__59835;
    wire N__59832;
    wire N__59827;
    wire N__59824;
    wire N__59821;
    wire N__59818;
    wire N__59815;
    wire N__59802;
    wire N__59799;
    wire N__59796;
    wire N__59793;
    wire N__59790;
    wire N__59787;
    wire N__59784;
    wire N__59781;
    wire N__59778;
    wire N__59775;
    wire N__59772;
    wire N__59769;
    wire N__59766;
    wire N__59763;
    wire N__59760;
    wire N__59757;
    wire N__59754;
    wire N__59753;
    wire N__59750;
    wire N__59747;
    wire N__59744;
    wire N__59741;
    wire N__59736;
    wire N__59733;
    wire N__59730;
    wire N__59727;
    wire N__59724;
    wire N__59721;
    wire N__59718;
    wire N__59717;
    wire N__59716;
    wire N__59715;
    wire N__59712;
    wire N__59709;
    wire N__59706;
    wire N__59701;
    wire N__59698;
    wire N__59695;
    wire N__59692;
    wire N__59687;
    wire N__59684;
    wire N__59679;
    wire N__59676;
    wire N__59673;
    wire N__59670;
    wire N__59667;
    wire N__59666;
    wire N__59663;
    wire N__59662;
    wire N__59661;
    wire N__59658;
    wire N__59655;
    wire N__59652;
    wire N__59647;
    wire N__59640;
    wire N__59637;
    wire N__59634;
    wire N__59631;
    wire N__59628;
    wire N__59625;
    wire N__59622;
    wire N__59619;
    wire N__59618;
    wire N__59615;
    wire N__59612;
    wire N__59609;
    wire N__59604;
    wire N__59601;
    wire N__59598;
    wire N__59595;
    wire N__59592;
    wire N__59589;
    wire N__59586;
    wire N__59583;
    wire N__59580;
    wire N__59577;
    wire N__59574;
    wire N__59571;
    wire N__59568;
    wire N__59565;
    wire N__59562;
    wire N__59559;
    wire N__59556;
    wire N__59553;
    wire N__59550;
    wire N__59547;
    wire N__59544;
    wire N__59541;
    wire N__59538;
    wire N__59535;
    wire N__59532;
    wire N__59529;
    wire N__59526;
    wire N__59523;
    wire N__59520;
    wire N__59517;
    wire N__59514;
    wire N__59513;
    wire N__59510;
    wire N__59507;
    wire N__59504;
    wire N__59501;
    wire N__59496;
    wire N__59493;
    wire N__59490;
    wire N__59487;
    wire N__59484;
    wire N__59481;
    wire N__59478;
    wire N__59475;
    wire N__59472;
    wire N__59469;
    wire N__59466;
    wire N__59463;
    wire N__59462;
    wire N__59459;
    wire N__59456;
    wire N__59455;
    wire N__59452;
    wire N__59449;
    wire N__59446;
    wire N__59441;
    wire N__59438;
    wire N__59437;
    wire N__59436;
    wire N__59435;
    wire N__59432;
    wire N__59429;
    wire N__59426;
    wire N__59423;
    wire N__59420;
    wire N__59409;
    wire N__59406;
    wire N__59403;
    wire N__59400;
    wire N__59397;
    wire N__59394;
    wire N__59391;
    wire N__59388;
    wire N__59385;
    wire N__59382;
    wire N__59379;
    wire N__59376;
    wire N__59373;
    wire N__59370;
    wire N__59367;
    wire N__59364;
    wire N__59361;
    wire N__59358;
    wire N__59355;
    wire N__59352;
    wire N__59349;
    wire N__59346;
    wire N__59343;
    wire N__59340;
    wire N__59337;
    wire N__59334;
    wire N__59333;
    wire N__59332;
    wire N__59329;
    wire N__59326;
    wire N__59323;
    wire N__59320;
    wire N__59319;
    wire N__59318;
    wire N__59315;
    wire N__59312;
    wire N__59309;
    wire N__59304;
    wire N__59303;
    wire N__59302;
    wire N__59297;
    wire N__59292;
    wire N__59287;
    wire N__59286;
    wire N__59281;
    wire N__59278;
    wire N__59275;
    wire N__59274;
    wire N__59271;
    wire N__59266;
    wire N__59263;
    wire N__59256;
    wire N__59253;
    wire N__59250;
    wire N__59247;
    wire N__59246;
    wire N__59243;
    wire N__59240;
    wire N__59235;
    wire N__59232;
    wire N__59229;
    wire N__59226;
    wire N__59223;
    wire N__59220;
    wire N__59217;
    wire N__59214;
    wire N__59211;
    wire N__59208;
    wire N__59205;
    wire N__59204;
    wire N__59201;
    wire N__59198;
    wire N__59197;
    wire N__59196;
    wire N__59195;
    wire N__59192;
    wire N__59189;
    wire N__59186;
    wire N__59183;
    wire N__59182;
    wire N__59179;
    wire N__59176;
    wire N__59173;
    wire N__59168;
    wire N__59167;
    wire N__59166;
    wire N__59163;
    wire N__59160;
    wire N__59157;
    wire N__59154;
    wire N__59151;
    wire N__59148;
    wire N__59147;
    wire N__59144;
    wire N__59139;
    wire N__59136;
    wire N__59131;
    wire N__59128;
    wire N__59125;
    wire N__59112;
    wire N__59109;
    wire N__59106;
    wire N__59105;
    wire N__59104;
    wire N__59101;
    wire N__59098;
    wire N__59095;
    wire N__59094;
    wire N__59093;
    wire N__59090;
    wire N__59087;
    wire N__59084;
    wire N__59081;
    wire N__59078;
    wire N__59075;
    wire N__59072;
    wire N__59067;
    wire N__59064;
    wire N__59063;
    wire N__59056;
    wire N__59053;
    wire N__59050;
    wire N__59049;
    wire N__59046;
    wire N__59041;
    wire N__59038;
    wire N__59031;
    wire N__59028;
    wire N__59025;
    wire N__59024;
    wire N__59023;
    wire N__59020;
    wire N__59017;
    wire N__59016;
    wire N__59013;
    wire N__59012;
    wire N__59009;
    wire N__59006;
    wire N__59003;
    wire N__59000;
    wire N__58997;
    wire N__58994;
    wire N__58991;
    wire N__58988;
    wire N__58983;
    wire N__58982;
    wire N__58975;
    wire N__58972;
    wire N__58969;
    wire N__58968;
    wire N__58967;
    wire N__58966;
    wire N__58963;
    wire N__58958;
    wire N__58955;
    wire N__58950;
    wire N__58941;
    wire N__58938;
    wire N__58935;
    wire N__58934;
    wire N__58931;
    wire N__58930;
    wire N__58929;
    wire N__58928;
    wire N__58925;
    wire N__58922;
    wire N__58919;
    wire N__58918;
    wire N__58915;
    wire N__58912;
    wire N__58909;
    wire N__58906;
    wire N__58903;
    wire N__58900;
    wire N__58897;
    wire N__58894;
    wire N__58891;
    wire N__58888;
    wire N__58885;
    wire N__58878;
    wire N__58877;
    wire N__58876;
    wire N__58875;
    wire N__58870;
    wire N__58865;
    wire N__58862;
    wire N__58857;
    wire N__58848;
    wire N__58845;
    wire N__58842;
    wire N__58841;
    wire N__58838;
    wire N__58835;
    wire N__58834;
    wire N__58833;
    wire N__58830;
    wire N__58829;
    wire N__58826;
    wire N__58825;
    wire N__58822;
    wire N__58819;
    wire N__58816;
    wire N__58813;
    wire N__58810;
    wire N__58807;
    wire N__58804;
    wire N__58801;
    wire N__58796;
    wire N__58791;
    wire N__58790;
    wire N__58787;
    wire N__58784;
    wire N__58781;
    wire N__58778;
    wire N__58775;
    wire N__58764;
    wire N__58761;
    wire N__58758;
    wire N__58757;
    wire N__58754;
    wire N__58753;
    wire N__58752;
    wire N__58749;
    wire N__58746;
    wire N__58743;
    wire N__58742;
    wire N__58739;
    wire N__58738;
    wire N__58735;
    wire N__58732;
    wire N__58729;
    wire N__58726;
    wire N__58725;
    wire N__58722;
    wire N__58719;
    wire N__58716;
    wire N__58713;
    wire N__58708;
    wire N__58705;
    wire N__58702;
    wire N__58699;
    wire N__58698;
    wire N__58697;
    wire N__58694;
    wire N__58689;
    wire N__58686;
    wire N__58681;
    wire N__58676;
    wire N__58665;
    wire N__58662;
    wire N__58659;
    wire N__58658;
    wire N__58655;
    wire N__58652;
    wire N__58651;
    wire N__58648;
    wire N__58645;
    wire N__58644;
    wire N__58643;
    wire N__58640;
    wire N__58635;
    wire N__58634;
    wire N__58631;
    wire N__58628;
    wire N__58627;
    wire N__58624;
    wire N__58621;
    wire N__58618;
    wire N__58615;
    wire N__58612;
    wire N__58609;
    wire N__58606;
    wire N__58603;
    wire N__58596;
    wire N__58593;
    wire N__58584;
    wire N__58581;
    wire N__58578;
    wire N__58575;
    wire N__58572;
    wire N__58569;
    wire N__58566;
    wire N__58563;
    wire N__58560;
    wire N__58557;
    wire N__58554;
    wire N__58551;
    wire N__58548;
    wire N__58545;
    wire N__58542;
    wire N__58539;
    wire N__58536;
    wire N__58533;
    wire N__58532;
    wire N__58529;
    wire N__58526;
    wire N__58523;
    wire N__58518;
    wire N__58515;
    wire N__58512;
    wire N__58511;
    wire N__58508;
    wire N__58505;
    wire N__58500;
    wire N__58497;
    wire N__58494;
    wire N__58491;
    wire N__58488;
    wire N__58485;
    wire N__58482;
    wire N__58479;
    wire N__58476;
    wire N__58473;
    wire N__58470;
    wire N__58467;
    wire N__58464;
    wire N__58461;
    wire N__58458;
    wire N__58455;
    wire N__58452;
    wire N__58449;
    wire N__58446;
    wire N__58443;
    wire N__58440;
    wire N__58437;
    wire N__58434;
    wire N__58431;
    wire N__58428;
    wire N__58425;
    wire N__58424;
    wire N__58421;
    wire N__58418;
    wire N__58413;
    wire N__58410;
    wire N__58407;
    wire N__58404;
    wire N__58401;
    wire N__58398;
    wire N__58395;
    wire N__58394;
    wire N__58389;
    wire N__58386;
    wire N__58383;
    wire N__58380;
    wire N__58379;
    wire N__58378;
    wire N__58371;
    wire N__58368;
    wire N__58365;
    wire N__58362;
    wire N__58359;
    wire N__58356;
    wire N__58353;
    wire N__58350;
    wire N__58347;
    wire N__58344;
    wire N__58341;
    wire N__58338;
    wire N__58335;
    wire N__58332;
    wire N__58329;
    wire N__58328;
    wire N__58325;
    wire N__58322;
    wire N__58317;
    wire N__58314;
    wire N__58311;
    wire N__58310;
    wire N__58307;
    wire N__58304;
    wire N__58301;
    wire N__58298;
    wire N__58293;
    wire N__58292;
    wire N__58291;
    wire N__58288;
    wire N__58285;
    wire N__58282;
    wire N__58281;
    wire N__58278;
    wire N__58275;
    wire N__58272;
    wire N__58269;
    wire N__58266;
    wire N__58261;
    wire N__58258;
    wire N__58251;
    wire N__58248;
    wire N__58247;
    wire N__58246;
    wire N__58245;
    wire N__58242;
    wire N__58239;
    wire N__58236;
    wire N__58233;
    wire N__58230;
    wire N__58227;
    wire N__58224;
    wire N__58221;
    wire N__58218;
    wire N__58215;
    wire N__58206;
    wire N__58203;
    wire N__58202;
    wire N__58199;
    wire N__58196;
    wire N__58193;
    wire N__58188;
    wire N__58185;
    wire N__58182;
    wire N__58181;
    wire N__58178;
    wire N__58175;
    wire N__58172;
    wire N__58169;
    wire N__58166;
    wire N__58161;
    wire N__58158;
    wire N__58157;
    wire N__58156;
    wire N__58153;
    wire N__58152;
    wire N__58151;
    wire N__58148;
    wire N__58145;
    wire N__58136;
    wire N__58131;
    wire N__58128;
    wire N__58125;
    wire N__58122;
    wire N__58121;
    wire N__58120;
    wire N__58119;
    wire N__58118;
    wire N__58115;
    wire N__58112;
    wire N__58111;
    wire N__58110;
    wire N__58109;
    wire N__58108;
    wire N__58107;
    wire N__58104;
    wire N__58103;
    wire N__58102;
    wire N__58097;
    wire N__58092;
    wire N__58075;
    wire N__58068;
    wire N__58067;
    wire N__58064;
    wire N__58061;
    wire N__58060;
    wire N__58057;
    wire N__58054;
    wire N__58051;
    wire N__58046;
    wire N__58043;
    wire N__58040;
    wire N__58035;
    wire N__58034;
    wire N__58029;
    wire N__58028;
    wire N__58025;
    wire N__58022;
    wire N__58019;
    wire N__58014;
    wire N__58013;
    wire N__58012;
    wire N__58011;
    wire N__58010;
    wire N__58009;
    wire N__58006;
    wire N__58005;
    wire N__58004;
    wire N__58001;
    wire N__57998;
    wire N__57995;
    wire N__57994;
    wire N__57991;
    wire N__57990;
    wire N__57987;
    wire N__57984;
    wire N__57983;
    wire N__57982;
    wire N__57979;
    wire N__57978;
    wire N__57975;
    wire N__57970;
    wire N__57967;
    wire N__57964;
    wire N__57963;
    wire N__57960;
    wire N__57957;
    wire N__57952;
    wire N__57949;
    wire N__57946;
    wire N__57943;
    wire N__57940;
    wire N__57931;
    wire N__57928;
    wire N__57909;
    wire N__57906;
    wire N__57905;
    wire N__57904;
    wire N__57901;
    wire N__57896;
    wire N__57893;
    wire N__57888;
    wire N__57885;
    wire N__57882;
    wire N__57879;
    wire N__57876;
    wire N__57873;
    wire N__57870;
    wire N__57869;
    wire N__57866;
    wire N__57863;
    wire N__57862;
    wire N__57859;
    wire N__57856;
    wire N__57853;
    wire N__57848;
    wire N__57843;
    wire N__57840;
    wire N__57837;
    wire N__57834;
    wire N__57831;
    wire N__57828;
    wire N__57825;
    wire N__57824;
    wire N__57821;
    wire N__57818;
    wire N__57813;
    wire N__57810;
    wire N__57807;
    wire N__57804;
    wire N__57801;
    wire N__57798;
    wire N__57795;
    wire N__57794;
    wire N__57791;
    wire N__57788;
    wire N__57785;
    wire N__57782;
    wire N__57781;
    wire N__57778;
    wire N__57775;
    wire N__57772;
    wire N__57767;
    wire N__57762;
    wire N__57759;
    wire N__57758;
    wire N__57755;
    wire N__57752;
    wire N__57749;
    wire N__57746;
    wire N__57741;
    wire N__57738;
    wire N__57735;
    wire N__57732;
    wire N__57729;
    wire N__57726;
    wire N__57723;
    wire N__57720;
    wire N__57717;
    wire N__57714;
    wire N__57711;
    wire N__57710;
    wire N__57707;
    wire N__57704;
    wire N__57703;
    wire N__57702;
    wire N__57699;
    wire N__57696;
    wire N__57691;
    wire N__57690;
    wire N__57689;
    wire N__57682;
    wire N__57681;
    wire N__57680;
    wire N__57679;
    wire N__57676;
    wire N__57673;
    wire N__57670;
    wire N__57667;
    wire N__57662;
    wire N__57657;
    wire N__57648;
    wire N__57647;
    wire N__57644;
    wire N__57641;
    wire N__57638;
    wire N__57635;
    wire N__57632;
    wire N__57629;
    wire N__57626;
    wire N__57625;
    wire N__57624;
    wire N__57621;
    wire N__57618;
    wire N__57613;
    wire N__57606;
    wire N__57603;
    wire N__57602;
    wire N__57601;
    wire N__57598;
    wire N__57597;
    wire N__57594;
    wire N__57593;
    wire N__57590;
    wire N__57587;
    wire N__57580;
    wire N__57573;
    wire N__57572;
    wire N__57569;
    wire N__57566;
    wire N__57563;
    wire N__57560;
    wire N__57557;
    wire N__57554;
    wire N__57551;
    wire N__57548;
    wire N__57545;
    wire N__57540;
    wire N__57537;
    wire N__57536;
    wire N__57533;
    wire N__57530;
    wire N__57527;
    wire N__57524;
    wire N__57521;
    wire N__57518;
    wire N__57513;
    wire N__57510;
    wire N__57509;
    wire N__57506;
    wire N__57505;
    wire N__57502;
    wire N__57499;
    wire N__57494;
    wire N__57493;
    wire N__57488;
    wire N__57485;
    wire N__57482;
    wire N__57477;
    wire N__57474;
    wire N__57471;
    wire N__57470;
    wire N__57467;
    wire N__57464;
    wire N__57461;
    wire N__57458;
    wire N__57453;
    wire N__57450;
    wire N__57449;
    wire N__57446;
    wire N__57443;
    wire N__57440;
    wire N__57437;
    wire N__57436;
    wire N__57431;
    wire N__57428;
    wire N__57425;
    wire N__57422;
    wire N__57417;
    wire N__57416;
    wire N__57413;
    wire N__57410;
    wire N__57407;
    wire N__57406;
    wire N__57403;
    wire N__57400;
    wire N__57397;
    wire N__57392;
    wire N__57389;
    wire N__57386;
    wire N__57383;
    wire N__57378;
    wire N__57377;
    wire N__57374;
    wire N__57371;
    wire N__57368;
    wire N__57365;
    wire N__57362;
    wire N__57361;
    wire N__57356;
    wire N__57353;
    wire N__57350;
    wire N__57345;
    wire N__57342;
    wire N__57339;
    wire N__57336;
    wire N__57333;
    wire N__57332;
    wire N__57331;
    wire N__57330;
    wire N__57327;
    wire N__57324;
    wire N__57321;
    wire N__57318;
    wire N__57315;
    wire N__57312;
    wire N__57309;
    wire N__57306;
    wire N__57301;
    wire N__57298;
    wire N__57295;
    wire N__57288;
    wire N__57285;
    wire N__57282;
    wire N__57279;
    wire N__57276;
    wire N__57273;
    wire N__57270;
    wire N__57267;
    wire N__57266;
    wire N__57263;
    wire N__57262;
    wire N__57261;
    wire N__57258;
    wire N__57257;
    wire N__57256;
    wire N__57255;
    wire N__57254;
    wire N__57253;
    wire N__57250;
    wire N__57247;
    wire N__57244;
    wire N__57239;
    wire N__57234;
    wire N__57229;
    wire N__57216;
    wire N__57213;
    wire N__57212;
    wire N__57211;
    wire N__57210;
    wire N__57209;
    wire N__57206;
    wire N__57203;
    wire N__57200;
    wire N__57195;
    wire N__57186;
    wire N__57185;
    wire N__57184;
    wire N__57183;
    wire N__57182;
    wire N__57179;
    wire N__57176;
    wire N__57173;
    wire N__57170;
    wire N__57167;
    wire N__57166;
    wire N__57163;
    wire N__57160;
    wire N__57159;
    wire N__57158;
    wire N__57157;
    wire N__57156;
    wire N__57155;
    wire N__57152;
    wire N__57151;
    wire N__57148;
    wire N__57145;
    wire N__57144;
    wire N__57141;
    wire N__57136;
    wire N__57133;
    wire N__57128;
    wire N__57125;
    wire N__57124;
    wire N__57123;
    wire N__57122;
    wire N__57119;
    wire N__57116;
    wire N__57113;
    wire N__57108;
    wire N__57105;
    wire N__57100;
    wire N__57093;
    wire N__57086;
    wire N__57069;
    wire N__57068;
    wire N__57067;
    wire N__57066;
    wire N__57063;
    wire N__57060;
    wire N__57059;
    wire N__57058;
    wire N__57057;
    wire N__57056;
    wire N__57053;
    wire N__57052;
    wire N__57051;
    wire N__57048;
    wire N__57043;
    wire N__57040;
    wire N__57039;
    wire N__57034;
    wire N__57031;
    wire N__57028;
    wire N__57027;
    wire N__57026;
    wire N__57025;
    wire N__57022;
    wire N__57019;
    wire N__57016;
    wire N__57011;
    wire N__57010;
    wire N__57009;
    wire N__57006;
    wire N__56999;
    wire N__56994;
    wire N__56991;
    wire N__56988;
    wire N__56981;
    wire N__56978;
    wire N__56975;
    wire N__56958;
    wire N__56955;
    wire N__56952;
    wire N__56949;
    wire N__56948;
    wire N__56947;
    wire N__56946;
    wire N__56945;
    wire N__56944;
    wire N__56941;
    wire N__56940;
    wire N__56939;
    wire N__56938;
    wire N__56937;
    wire N__56936;
    wire N__56935;
    wire N__56932;
    wire N__56929;
    wire N__56928;
    wire N__56925;
    wire N__56924;
    wire N__56921;
    wire N__56918;
    wire N__56915;
    wire N__56912;
    wire N__56909;
    wire N__56904;
    wire N__56899;
    wire N__56894;
    wire N__56891;
    wire N__56888;
    wire N__56885;
    wire N__56882;
    wire N__56879;
    wire N__56876;
    wire N__56871;
    wire N__56868;
    wire N__56865;
    wire N__56864;
    wire N__56863;
    wire N__56856;
    wire N__56853;
    wire N__56846;
    wire N__56839;
    wire N__56834;
    wire N__56829;
    wire N__56820;
    wire N__56817;
    wire N__56816;
    wire N__56813;
    wire N__56810;
    wire N__56807;
    wire N__56804;
    wire N__56803;
    wire N__56798;
    wire N__56795;
    wire N__56792;
    wire N__56787;
    wire N__56784;
    wire N__56781;
    wire N__56780;
    wire N__56779;
    wire N__56776;
    wire N__56773;
    wire N__56770;
    wire N__56765;
    wire N__56762;
    wire N__56759;
    wire N__56754;
    wire N__56751;
    wire N__56748;
    wire N__56745;
    wire N__56742;
    wire N__56739;
    wire N__56736;
    wire N__56733;
    wire N__56730;
    wire N__56727;
    wire N__56724;
    wire N__56721;
    wire N__56720;
    wire N__56719;
    wire N__56716;
    wire N__56715;
    wire N__56710;
    wire N__56707;
    wire N__56704;
    wire N__56701;
    wire N__56698;
    wire N__56695;
    wire N__56692;
    wire N__56685;
    wire N__56682;
    wire N__56679;
    wire N__56676;
    wire N__56673;
    wire N__56670;
    wire N__56667;
    wire N__56666;
    wire N__56663;
    wire N__56660;
    wire N__56657;
    wire N__56654;
    wire N__56653;
    wire N__56652;
    wire N__56647;
    wire N__56644;
    wire N__56641;
    wire N__56640;
    wire N__56639;
    wire N__56638;
    wire N__56637;
    wire N__56636;
    wire N__56635;
    wire N__56634;
    wire N__56633;
    wire N__56632;
    wire N__56631;
    wire N__56630;
    wire N__56623;
    wire N__56620;
    wire N__56617;
    wire N__56614;
    wire N__56611;
    wire N__56608;
    wire N__56605;
    wire N__56602;
    wire N__56599;
    wire N__56596;
    wire N__56595;
    wire N__56594;
    wire N__56591;
    wire N__56588;
    wire N__56581;
    wire N__56580;
    wire N__56577;
    wire N__56576;
    wire N__56575;
    wire N__56570;
    wire N__56559;
    wire N__56554;
    wire N__56553;
    wire N__56552;
    wire N__56551;
    wire N__56550;
    wire N__56549;
    wire N__56548;
    wire N__56547;
    wire N__56546;
    wire N__56543;
    wire N__56540;
    wire N__56539;
    wire N__56536;
    wire N__56535;
    wire N__56532;
    wire N__56529;
    wire N__56528;
    wire N__56525;
    wire N__56524;
    wire N__56523;
    wire N__56520;
    wire N__56515;
    wire N__56514;
    wire N__56511;
    wire N__56508;
    wire N__56507;
    wire N__56506;
    wire N__56503;
    wire N__56500;
    wire N__56497;
    wire N__56494;
    wire N__56491;
    wire N__56488;
    wire N__56485;
    wire N__56484;
    wire N__56483;
    wire N__56480;
    wire N__56477;
    wire N__56474;
    wire N__56471;
    wire N__56466;
    wire N__56463;
    wire N__56460;
    wire N__56459;
    wire N__56456;
    wire N__56453;
    wire N__56448;
    wire N__56441;
    wire N__56438;
    wire N__56435;
    wire N__56432;
    wire N__56429;
    wire N__56426;
    wire N__56421;
    wire N__56418;
    wire N__56415;
    wire N__56412;
    wire N__56409;
    wire N__56406;
    wire N__56403;
    wire N__56400;
    wire N__56397;
    wire N__56392;
    wire N__56389;
    wire N__56382;
    wire N__56377;
    wire N__56374;
    wire N__56371;
    wire N__56362;
    wire N__56359;
    wire N__56354;
    wire N__56351;
    wire N__56348;
    wire N__56339;
    wire N__56334;
    wire N__56329;
    wire N__56326;
    wire N__56323;
    wire N__56316;
    wire N__56309;
    wire N__56306;
    wire N__56295;
    wire N__56292;
    wire N__56291;
    wire N__56288;
    wire N__56285;
    wire N__56280;
    wire N__56279;
    wire N__56276;
    wire N__56273;
    wire N__56270;
    wire N__56265;
    wire N__56264;
    wire N__56261;
    wire N__56256;
    wire N__56253;
    wire N__56252;
    wire N__56251;
    wire N__56248;
    wire N__56245;
    wire N__56242;
    wire N__56239;
    wire N__56236;
    wire N__56233;
    wire N__56230;
    wire N__56227;
    wire N__56220;
    wire N__56219;
    wire N__56214;
    wire N__56211;
    wire N__56210;
    wire N__56205;
    wire N__56202;
    wire N__56199;
    wire N__56198;
    wire N__56195;
    wire N__56192;
    wire N__56189;
    wire N__56184;
    wire N__56183;
    wire N__56178;
    wire N__56175;
    wire N__56174;
    wire N__56173;
    wire N__56170;
    wire N__56165;
    wire N__56162;
    wire N__56159;
    wire N__56154;
    wire N__56153;
    wire N__56150;
    wire N__56145;
    wire N__56142;
    wire N__56139;
    wire N__56136;
    wire N__56133;
    wire N__56130;
    wire N__56129;
    wire N__56126;
    wire N__56123;
    wire N__56118;
    wire N__56117;
    wire N__56114;
    wire N__56111;
    wire N__56108;
    wire N__56105;
    wire N__56100;
    wire N__56097;
    wire N__56094;
    wire N__56093;
    wire N__56088;
    wire N__56087;
    wire N__56086;
    wire N__56085;
    wire N__56084;
    wire N__56083;
    wire N__56082;
    wire N__56081;
    wire N__56080;
    wire N__56079;
    wire N__56078;
    wire N__56077;
    wire N__56076;
    wire N__56075;
    wire N__56072;
    wire N__56043;
    wire N__56040;
    wire N__56037;
    wire N__56034;
    wire N__56031;
    wire N__56030;
    wire N__56027;
    wire N__56024;
    wire N__56021;
    wire N__56020;
    wire N__56019;
    wire N__56018;
    wire N__56015;
    wire N__56012;
    wire N__56009;
    wire N__56004;
    wire N__55999;
    wire N__55996;
    wire N__55989;
    wire N__55986;
    wire N__55983;
    wire N__55980;
    wire N__55977;
    wire N__55974;
    wire N__55971;
    wire N__55968;
    wire N__55965;
    wire N__55962;
    wire N__55959;
    wire N__55956;
    wire N__55955;
    wire N__55954;
    wire N__55953;
    wire N__55952;
    wire N__55951;
    wire N__55948;
    wire N__55945;
    wire N__55944;
    wire N__55943;
    wire N__55942;
    wire N__55941;
    wire N__55940;
    wire N__55939;
    wire N__55938;
    wire N__55937;
    wire N__55936;
    wire N__55933;
    wire N__55930;
    wire N__55927;
    wire N__55924;
    wire N__55909;
    wire N__55908;
    wire N__55905;
    wire N__55902;
    wire N__55899;
    wire N__55896;
    wire N__55895;
    wire N__55894;
    wire N__55891;
    wire N__55886;
    wire N__55883;
    wire N__55880;
    wire N__55877;
    wire N__55876;
    wire N__55873;
    wire N__55862;
    wire N__55859;
    wire N__55854;
    wire N__55851;
    wire N__55846;
    wire N__55841;
    wire N__55834;
    wire N__55827;
    wire N__55824;
    wire N__55823;
    wire N__55822;
    wire N__55819;
    wire N__55814;
    wire N__55809;
    wire N__55808;
    wire N__55807;
    wire N__55806;
    wire N__55805;
    wire N__55804;
    wire N__55803;
    wire N__55800;
    wire N__55797;
    wire N__55792;
    wire N__55791;
    wire N__55788;
    wire N__55787;
    wire N__55784;
    wire N__55783;
    wire N__55782;
    wire N__55781;
    wire N__55780;
    wire N__55777;
    wire N__55776;
    wire N__55775;
    wire N__55774;
    wire N__55773;
    wire N__55770;
    wire N__55765;
    wire N__55752;
    wire N__55737;
    wire N__55728;
    wire N__55725;
    wire N__55724;
    wire N__55721;
    wire N__55718;
    wire N__55713;
    wire N__55712;
    wire N__55709;
    wire N__55706;
    wire N__55703;
    wire N__55698;
    wire N__55695;
    wire N__55694;
    wire N__55689;
    wire N__55686;
    wire N__55685;
    wire N__55682;
    wire N__55679;
    wire N__55676;
    wire N__55671;
    wire N__55668;
    wire N__55665;
    wire N__55664;
    wire N__55659;
    wire N__55656;
    wire N__55655;
    wire N__55652;
    wire N__55649;
    wire N__55646;
    wire N__55641;
    wire N__55638;
    wire N__55635;
    wire N__55634;
    wire N__55629;
    wire N__55626;
    wire N__55625;
    wire N__55622;
    wire N__55619;
    wire N__55616;
    wire N__55611;
    wire N__55608;
    wire N__55605;
    wire N__55604;
    wire N__55603;
    wire N__55600;
    wire N__55599;
    wire N__55596;
    wire N__55595;
    wire N__55594;
    wire N__55593;
    wire N__55592;
    wire N__55591;
    wire N__55590;
    wire N__55579;
    wire N__55576;
    wire N__55575;
    wire N__55572;
    wire N__55571;
    wire N__55568;
    wire N__55567;
    wire N__55564;
    wire N__55563;
    wire N__55562;
    wire N__55559;
    wire N__55558;
    wire N__55555;
    wire N__55538;
    wire N__55531;
    wire N__55524;
    wire N__55521;
    wire N__55520;
    wire N__55515;
    wire N__55512;
    wire N__55511;
    wire N__55508;
    wire N__55505;
    wire N__55502;
    wire N__55497;
    wire N__55496;
    wire N__55493;
    wire N__55492;
    wire N__55489;
    wire N__55486;
    wire N__55481;
    wire N__55478;
    wire N__55475;
    wire N__55472;
    wire N__55469;
    wire N__55464;
    wire N__55461;
    wire N__55460;
    wire N__55459;
    wire N__55458;
    wire N__55455;
    wire N__55452;
    wire N__55449;
    wire N__55446;
    wire N__55441;
    wire N__55438;
    wire N__55435;
    wire N__55432;
    wire N__55429;
    wire N__55422;
    wire N__55419;
    wire N__55418;
    wire N__55415;
    wire N__55414;
    wire N__55411;
    wire N__55408;
    wire N__55405;
    wire N__55402;
    wire N__55399;
    wire N__55396;
    wire N__55391;
    wire N__55388;
    wire N__55383;
    wire N__55380;
    wire N__55379;
    wire N__55378;
    wire N__55375;
    wire N__55370;
    wire N__55367;
    wire N__55364;
    wire N__55361;
    wire N__55358;
    wire N__55353;
    wire N__55350;
    wire N__55347;
    wire N__55346;
    wire N__55345;
    wire N__55342;
    wire N__55339;
    wire N__55336;
    wire N__55331;
    wire N__55326;
    wire N__55323;
    wire N__55320;
    wire N__55319;
    wire N__55316;
    wire N__55313;
    wire N__55312;
    wire N__55309;
    wire N__55306;
    wire N__55303;
    wire N__55298;
    wire N__55295;
    wire N__55290;
    wire N__55287;
    wire N__55286;
    wire N__55283;
    wire N__55282;
    wire N__55279;
    wire N__55276;
    wire N__55273;
    wire N__55270;
    wire N__55267;
    wire N__55264;
    wire N__55257;
    wire N__55254;
    wire N__55251;
    wire N__55250;
    wire N__55245;
    wire N__55242;
    wire N__55241;
    wire N__55238;
    wire N__55235;
    wire N__55232;
    wire N__55227;
    wire N__55224;
    wire N__55221;
    wire N__55218;
    wire N__55215;
    wire N__55212;
    wire N__55211;
    wire N__55208;
    wire N__55205;
    wire N__55202;
    wire N__55197;
    wire N__55196;
    wire N__55195;
    wire N__55194;
    wire N__55191;
    wire N__55186;
    wire N__55183;
    wire N__55178;
    wire N__55175;
    wire N__55172;
    wire N__55169;
    wire N__55166;
    wire N__55161;
    wire N__55158;
    wire N__55155;
    wire N__55152;
    wire N__55151;
    wire N__55150;
    wire N__55145;
    wire N__55142;
    wire N__55139;
    wire N__55136;
    wire N__55133;
    wire N__55128;
    wire N__55125;
    wire N__55122;
    wire N__55119;
    wire N__55116;
    wire N__55115;
    wire N__55114;
    wire N__55111;
    wire N__55106;
    wire N__55103;
    wire N__55100;
    wire N__55095;
    wire N__55092;
    wire N__55089;
    wire N__55086;
    wire N__55083;
    wire N__55082;
    wire N__55077;
    wire N__55076;
    wire N__55073;
    wire N__55070;
    wire N__55067;
    wire N__55064;
    wire N__55061;
    wire N__55056;
    wire N__55053;
    wire N__55050;
    wire N__55047;
    wire N__55044;
    wire N__55043;
    wire N__55042;
    wire N__55039;
    wire N__55034;
    wire N__55031;
    wire N__55028;
    wire N__55025;
    wire N__55022;
    wire N__55017;
    wire N__55014;
    wire N__55011;
    wire N__55008;
    wire N__55007;
    wire N__55006;
    wire N__55001;
    wire N__54998;
    wire N__54995;
    wire N__54992;
    wire N__54989;
    wire N__54984;
    wire N__54981;
    wire N__54978;
    wire N__54975;
    wire N__54972;
    wire N__54971;
    wire N__54968;
    wire N__54965;
    wire N__54964;
    wire N__54963;
    wire N__54960;
    wire N__54957;
    wire N__54952;
    wire N__54945;
    wire N__54942;
    wire N__54939;
    wire N__54936;
    wire N__54933;
    wire N__54932;
    wire N__54931;
    wire N__54926;
    wire N__54923;
    wire N__54920;
    wire N__54915;
    wire N__54912;
    wire N__54909;
    wire N__54906;
    wire N__54903;
    wire N__54900;
    wire N__54897;
    wire N__54894;
    wire N__54893;
    wire N__54890;
    wire N__54887;
    wire N__54882;
    wire N__54879;
    wire N__54876;
    wire N__54873;
    wire N__54870;
    wire N__54867;
    wire N__54864;
    wire N__54863;
    wire N__54860;
    wire N__54855;
    wire N__54852;
    wire N__54849;
    wire N__54846;
    wire N__54845;
    wire N__54842;
    wire N__54839;
    wire N__54836;
    wire N__54833;
    wire N__54830;
    wire N__54827;
    wire N__54824;
    wire N__54819;
    wire N__54816;
    wire N__54813;
    wire N__54810;
    wire N__54809;
    wire N__54808;
    wire N__54805;
    wire N__54802;
    wire N__54799;
    wire N__54796;
    wire N__54793;
    wire N__54790;
    wire N__54787;
    wire N__54784;
    wire N__54779;
    wire N__54774;
    wire N__54771;
    wire N__54768;
    wire N__54765;
    wire N__54762;
    wire N__54761;
    wire N__54758;
    wire N__54757;
    wire N__54754;
    wire N__54751;
    wire N__54748;
    wire N__54745;
    wire N__54742;
    wire N__54739;
    wire N__54736;
    wire N__54733;
    wire N__54726;
    wire N__54723;
    wire N__54720;
    wire N__54717;
    wire N__54716;
    wire N__54715;
    wire N__54712;
    wire N__54707;
    wire N__54704;
    wire N__54701;
    wire N__54696;
    wire N__54693;
    wire N__54690;
    wire N__54687;
    wire N__54684;
    wire N__54683;
    wire N__54682;
    wire N__54677;
    wire N__54674;
    wire N__54671;
    wire N__54668;
    wire N__54665;
    wire N__54662;
    wire N__54659;
    wire N__54654;
    wire N__54651;
    wire N__54648;
    wire N__54645;
    wire N__54642;
    wire N__54639;
    wire N__54636;
    wire N__54633;
    wire N__54630;
    wire N__54627;
    wire N__54624;
    wire N__54621;
    wire N__54618;
    wire N__54615;
    wire N__54612;
    wire N__54609;
    wire N__54606;
    wire N__54603;
    wire N__54600;
    wire N__54597;
    wire N__54594;
    wire N__54591;
    wire N__54588;
    wire N__54585;
    wire N__54582;
    wire N__54579;
    wire N__54576;
    wire N__54573;
    wire N__54570;
    wire N__54567;
    wire N__54564;
    wire N__54561;
    wire N__54558;
    wire N__54555;
    wire N__54552;
    wire N__54549;
    wire N__54546;
    wire N__54543;
    wire N__54540;
    wire N__54537;
    wire N__54534;
    wire N__54531;
    wire N__54528;
    wire N__54525;
    wire N__54522;
    wire N__54519;
    wire N__54516;
    wire N__54513;
    wire N__54510;
    wire N__54507;
    wire N__54506;
    wire N__54505;
    wire N__54502;
    wire N__54499;
    wire N__54496;
    wire N__54493;
    wire N__54490;
    wire N__54483;
    wire N__54480;
    wire N__54477;
    wire N__54476;
    wire N__54473;
    wire N__54470;
    wire N__54467;
    wire N__54462;
    wire N__54461;
    wire N__54458;
    wire N__54455;
    wire N__54452;
    wire N__54447;
    wire N__54444;
    wire N__54441;
    wire N__54438;
    wire N__54435;
    wire N__54432;
    wire N__54429;
    wire N__54426;
    wire N__54423;
    wire N__54420;
    wire N__54417;
    wire N__54414;
    wire N__54411;
    wire N__54408;
    wire N__54405;
    wire N__54402;
    wire N__54399;
    wire N__54396;
    wire N__54393;
    wire N__54390;
    wire N__54387;
    wire N__54384;
    wire N__54381;
    wire N__54378;
    wire N__54377;
    wire N__54374;
    wire N__54371;
    wire N__54368;
    wire N__54365;
    wire N__54362;
    wire N__54359;
    wire N__54356;
    wire N__54353;
    wire N__54348;
    wire N__54347;
    wire N__54344;
    wire N__54341;
    wire N__54338;
    wire N__54335;
    wire N__54330;
    wire N__54327;
    wire N__54324;
    wire N__54321;
    wire N__54318;
    wire N__54315;
    wire N__54312;
    wire N__54309;
    wire N__54306;
    wire N__54303;
    wire N__54302;
    wire N__54301;
    wire N__54298;
    wire N__54295;
    wire N__54292;
    wire N__54291;
    wire N__54286;
    wire N__54283;
    wire N__54280;
    wire N__54277;
    wire N__54270;
    wire N__54269;
    wire N__54268;
    wire N__54265;
    wire N__54262;
    wire N__54259;
    wire N__54256;
    wire N__54255;
    wire N__54252;
    wire N__54249;
    wire N__54246;
    wire N__54243;
    wire N__54240;
    wire N__54237;
    wire N__54232;
    wire N__54227;
    wire N__54224;
    wire N__54219;
    wire N__54216;
    wire N__54213;
    wire N__54210;
    wire N__54207;
    wire N__54204;
    wire N__54201;
    wire N__54198;
    wire N__54195;
    wire N__54194;
    wire N__54191;
    wire N__54188;
    wire N__54185;
    wire N__54182;
    wire N__54179;
    wire N__54176;
    wire N__54173;
    wire N__54170;
    wire N__54165;
    wire N__54162;
    wire N__54159;
    wire N__54156;
    wire N__54153;
    wire N__54150;
    wire N__54147;
    wire N__54144;
    wire N__54141;
    wire N__54138;
    wire N__54135;
    wire N__54132;
    wire N__54129;
    wire N__54126;
    wire N__54125;
    wire N__54122;
    wire N__54119;
    wire N__54116;
    wire N__54113;
    wire N__54110;
    wire N__54107;
    wire N__54102;
    wire N__54099;
    wire N__54096;
    wire N__54093;
    wire N__54092;
    wire N__54087;
    wire N__54084;
    wire N__54081;
    wire N__54078;
    wire N__54075;
    wire N__54072;
    wire N__54069;
    wire N__54066;
    wire N__54063;
    wire N__54060;
    wire N__54057;
    wire N__54054;
    wire N__54051;
    wire N__54048;
    wire N__54045;
    wire N__54042;
    wire N__54041;
    wire N__54036;
    wire N__54033;
    wire N__54030;
    wire N__54027;
    wire N__54026;
    wire N__54023;
    wire N__54020;
    wire N__54019;
    wire N__54016;
    wire N__54011;
    wire N__54008;
    wire N__54003;
    wire N__54000;
    wire N__53999;
    wire N__53998;
    wire N__53993;
    wire N__53990;
    wire N__53985;
    wire N__53982;
    wire N__53979;
    wire N__53978;
    wire N__53975;
    wire N__53972;
    wire N__53969;
    wire N__53966;
    wire N__53965;
    wire N__53964;
    wire N__53963;
    wire N__53958;
    wire N__53955;
    wire N__53950;
    wire N__53947;
    wire N__53944;
    wire N__53939;
    wire N__53934;
    wire N__53931;
    wire N__53930;
    wire N__53927;
    wire N__53924;
    wire N__53921;
    wire N__53918;
    wire N__53913;
    wire N__53910;
    wire N__53907;
    wire N__53904;
    wire N__53901;
    wire N__53898;
    wire N__53897;
    wire N__53894;
    wire N__53891;
    wire N__53886;
    wire N__53883;
    wire N__53880;
    wire N__53877;
    wire N__53874;
    wire N__53871;
    wire N__53870;
    wire N__53867;
    wire N__53864;
    wire N__53861;
    wire N__53856;
    wire N__53855;
    wire N__53852;
    wire N__53849;
    wire N__53846;
    wire N__53843;
    wire N__53840;
    wire N__53837;
    wire N__53832;
    wire N__53829;
    wire N__53828;
    wire N__53825;
    wire N__53822;
    wire N__53819;
    wire N__53816;
    wire N__53811;
    wire N__53810;
    wire N__53807;
    wire N__53804;
    wire N__53801;
    wire N__53798;
    wire N__53793;
    wire N__53790;
    wire N__53787;
    wire N__53786;
    wire N__53783;
    wire N__53780;
    wire N__53775;
    wire N__53772;
    wire N__53769;
    wire N__53768;
    wire N__53765;
    wire N__53762;
    wire N__53759;
    wire N__53756;
    wire N__53753;
    wire N__53748;
    wire N__53745;
    wire N__53744;
    wire N__53741;
    wire N__53738;
    wire N__53733;
    wire N__53730;
    wire N__53727;
    wire N__53726;
    wire N__53723;
    wire N__53720;
    wire N__53715;
    wire N__53712;
    wire N__53709;
    wire N__53708;
    wire N__53705;
    wire N__53702;
    wire N__53699;
    wire N__53696;
    wire N__53691;
    wire N__53688;
    wire N__53685;
    wire N__53682;
    wire N__53679;
    wire N__53678;
    wire N__53675;
    wire N__53672;
    wire N__53671;
    wire N__53668;
    wire N__53665;
    wire N__53662;
    wire N__53657;
    wire N__53652;
    wire N__53651;
    wire N__53648;
    wire N__53647;
    wire N__53644;
    wire N__53641;
    wire N__53638;
    wire N__53635;
    wire N__53632;
    wire N__53625;
    wire N__53622;
    wire N__53619;
    wire N__53618;
    wire N__53615;
    wire N__53612;
    wire N__53611;
    wire N__53608;
    wire N__53605;
    wire N__53602;
    wire N__53597;
    wire N__53592;
    wire N__53589;
    wire N__53586;
    wire N__53583;
    wire N__53580;
    wire N__53579;
    wire N__53578;
    wire N__53575;
    wire N__53572;
    wire N__53569;
    wire N__53564;
    wire N__53559;
    wire N__53556;
    wire N__53555;
    wire N__53552;
    wire N__53549;
    wire N__53544;
    wire N__53543;
    wire N__53538;
    wire N__53535;
    wire N__53534;
    wire N__53531;
    wire N__53528;
    wire N__53525;
    wire N__53522;
    wire N__53519;
    wire N__53516;
    wire N__53511;
    wire N__53510;
    wire N__53507;
    wire N__53504;
    wire N__53501;
    wire N__53496;
    wire N__53493;
    wire N__53490;
    wire N__53487;
    wire N__53484;
    wire N__53481;
    wire N__53478;
    wire N__53475;
    wire N__53472;
    wire N__53469;
    wire N__53466;
    wire N__53463;
    wire N__53460;
    wire N__53457;
    wire N__53454;
    wire N__53451;
    wire N__53448;
    wire N__53445;
    wire N__53444;
    wire N__53441;
    wire N__53438;
    wire N__53437;
    wire N__53434;
    wire N__53431;
    wire N__53428;
    wire N__53425;
    wire N__53422;
    wire N__53415;
    wire N__53412;
    wire N__53409;
    wire N__53406;
    wire N__53403;
    wire N__53400;
    wire N__53397;
    wire N__53394;
    wire N__53391;
    wire N__53390;
    wire N__53385;
    wire N__53382;
    wire N__53381;
    wire N__53378;
    wire N__53373;
    wire N__53372;
    wire N__53369;
    wire N__53368;
    wire N__53365;
    wire N__53362;
    wire N__53359;
    wire N__53352;
    wire N__53349;
    wire N__53346;
    wire N__53343;
    wire N__53340;
    wire N__53339;
    wire N__53336;
    wire N__53333;
    wire N__53332;
    wire N__53329;
    wire N__53326;
    wire N__53323;
    wire N__53318;
    wire N__53313;
    wire N__53310;
    wire N__53307;
    wire N__53304;
    wire N__53301;
    wire N__53298;
    wire N__53295;
    wire N__53292;
    wire N__53289;
    wire N__53286;
    wire N__53285;
    wire N__53282;
    wire N__53279;
    wire N__53274;
    wire N__53271;
    wire N__53268;
    wire N__53265;
    wire N__53262;
    wire N__53259;
    wire N__53256;
    wire N__53255;
    wire N__53252;
    wire N__53251;
    wire N__53248;
    wire N__53245;
    wire N__53242;
    wire N__53235;
    wire N__53232;
    wire N__53231;
    wire N__53230;
    wire N__53227;
    wire N__53226;
    wire N__53223;
    wire N__53218;
    wire N__53215;
    wire N__53212;
    wire N__53209;
    wire N__53206;
    wire N__53203;
    wire N__53200;
    wire N__53193;
    wire N__53190;
    wire N__53187;
    wire N__53184;
    wire N__53181;
    wire N__53178;
    wire N__53175;
    wire N__53172;
    wire N__53169;
    wire N__53166;
    wire N__53163;
    wire N__53160;
    wire N__53157;
    wire N__53156;
    wire N__53153;
    wire N__53150;
    wire N__53145;
    wire N__53142;
    wire N__53139;
    wire N__53138;
    wire N__53137;
    wire N__53130;
    wire N__53127;
    wire N__53126;
    wire N__53125;
    wire N__53122;
    wire N__53119;
    wire N__53112;
    wire N__53109;
    wire N__53106;
    wire N__53105;
    wire N__53102;
    wire N__53099;
    wire N__53096;
    wire N__53093;
    wire N__53090;
    wire N__53087;
    wire N__53082;
    wire N__53079;
    wire N__53076;
    wire N__53073;
    wire N__53070;
    wire N__53067;
    wire N__53064;
    wire N__53063;
    wire N__53062;
    wire N__53059;
    wire N__53056;
    wire N__53055;
    wire N__53050;
    wire N__53047;
    wire N__53044;
    wire N__53041;
    wire N__53038;
    wire N__53035;
    wire N__53032;
    wire N__53025;
    wire N__53022;
    wire N__53019;
    wire N__53016;
    wire N__53015;
    wire N__53012;
    wire N__53009;
    wire N__53004;
    wire N__53001;
    wire N__52998;
    wire N__52995;
    wire N__52992;
    wire N__52989;
    wire N__52986;
    wire N__52983;
    wire N__52980;
    wire N__52977;
    wire N__52974;
    wire N__52971;
    wire N__52968;
    wire N__52965;
    wire N__52962;
    wire N__52959;
    wire N__52956;
    wire N__52953;
    wire N__52950;
    wire N__52947;
    wire N__52946;
    wire N__52945;
    wire N__52944;
    wire N__52943;
    wire N__52938;
    wire N__52935;
    wire N__52934;
    wire N__52931;
    wire N__52928;
    wire N__52923;
    wire N__52920;
    wire N__52917;
    wire N__52914;
    wire N__52913;
    wire N__52912;
    wire N__52911;
    wire N__52910;
    wire N__52909;
    wire N__52908;
    wire N__52905;
    wire N__52902;
    wire N__52899;
    wire N__52896;
    wire N__52893;
    wire N__52890;
    wire N__52881;
    wire N__52866;
    wire N__52865;
    wire N__52862;
    wire N__52859;
    wire N__52856;
    wire N__52853;
    wire N__52852;
    wire N__52849;
    wire N__52846;
    wire N__52843;
    wire N__52838;
    wire N__52833;
    wire N__52830;
    wire N__52829;
    wire N__52828;
    wire N__52827;
    wire N__52826;
    wire N__52821;
    wire N__52818;
    wire N__52817;
    wire N__52814;
    wire N__52811;
    wire N__52806;
    wire N__52803;
    wire N__52800;
    wire N__52797;
    wire N__52796;
    wire N__52795;
    wire N__52794;
    wire N__52793;
    wire N__52792;
    wire N__52791;
    wire N__52788;
    wire N__52783;
    wire N__52780;
    wire N__52777;
    wire N__52772;
    wire N__52765;
    wire N__52752;
    wire N__52751;
    wire N__52748;
    wire N__52747;
    wire N__52744;
    wire N__52741;
    wire N__52738;
    wire N__52735;
    wire N__52728;
    wire N__52725;
    wire N__52722;
    wire N__52719;
    wire N__52716;
    wire N__52713;
    wire N__52710;
    wire N__52707;
    wire N__52704;
    wire N__52701;
    wire N__52698;
    wire N__52695;
    wire N__52694;
    wire N__52689;
    wire N__52686;
    wire N__52683;
    wire N__52682;
    wire N__52677;
    wire N__52674;
    wire N__52671;
    wire N__52670;
    wire N__52669;
    wire N__52666;
    wire N__52661;
    wire N__52656;
    wire N__52653;
    wire N__52650;
    wire N__52647;
    wire N__52644;
    wire N__52643;
    wire N__52638;
    wire N__52635;
    wire N__52634;
    wire N__52631;
    wire N__52630;
    wire N__52627;
    wire N__52624;
    wire N__52621;
    wire N__52618;
    wire N__52615;
    wire N__52612;
    wire N__52609;
    wire N__52606;
    wire N__52599;
    wire N__52596;
    wire N__52593;
    wire N__52590;
    wire N__52589;
    wire N__52588;
    wire N__52587;
    wire N__52586;
    wire N__52585;
    wire N__52582;
    wire N__52571;
    wire N__52566;
    wire N__52565;
    wire N__52562;
    wire N__52559;
    wire N__52558;
    wire N__52557;
    wire N__52554;
    wire N__52547;
    wire N__52542;
    wire N__52541;
    wire N__52538;
    wire N__52535;
    wire N__52532;
    wire N__52529;
    wire N__52524;
    wire N__52523;
    wire N__52522;
    wire N__52519;
    wire N__52516;
    wire N__52513;
    wire N__52506;
    wire N__52503;
    wire N__52502;
    wire N__52497;
    wire N__52494;
    wire N__52491;
    wire N__52490;
    wire N__52487;
    wire N__52484;
    wire N__52479;
    wire N__52476;
    wire N__52473;
    wire N__52470;
    wire N__52469;
    wire N__52468;
    wire N__52465;
    wire N__52460;
    wire N__52455;
    wire N__52452;
    wire N__52451;
    wire N__52448;
    wire N__52447;
    wire N__52444;
    wire N__52441;
    wire N__52438;
    wire N__52433;
    wire N__52428;
    wire N__52425;
    wire N__52424;
    wire N__52421;
    wire N__52418;
    wire N__52417;
    wire N__52416;
    wire N__52415;
    wire N__52414;
    wire N__52401;
    wire N__52398;
    wire N__52397;
    wire N__52396;
    wire N__52395;
    wire N__52394;
    wire N__52393;
    wire N__52392;
    wire N__52391;
    wire N__52390;
    wire N__52389;
    wire N__52388;
    wire N__52387;
    wire N__52386;
    wire N__52369;
    wire N__52358;
    wire N__52353;
    wire N__52350;
    wire N__52347;
    wire N__52344;
    wire N__52341;
    wire N__52338;
    wire N__52335;
    wire N__52332;
    wire N__52331;
    wire N__52328;
    wire N__52325;
    wire N__52320;
    wire N__52317;
    wire N__52314;
    wire N__52311;
    wire N__52308;
    wire N__52305;
    wire N__52304;
    wire N__52301;
    wire N__52298;
    wire N__52295;
    wire N__52292;
    wire N__52287;
    wire N__52284;
    wire N__52281;
    wire N__52280;
    wire N__52279;
    wire N__52276;
    wire N__52273;
    wire N__52270;
    wire N__52265;
    wire N__52260;
    wire N__52257;
    wire N__52254;
    wire N__52253;
    wire N__52252;
    wire N__52251;
    wire N__52250;
    wire N__52245;
    wire N__52238;
    wire N__52233;
    wire N__52232;
    wire N__52231;
    wire N__52230;
    wire N__52225;
    wire N__52220;
    wire N__52215;
    wire N__52214;
    wire N__52211;
    wire N__52208;
    wire N__52203;
    wire N__52200;
    wire N__52199;
    wire N__52196;
    wire N__52193;
    wire N__52190;
    wire N__52187;
    wire N__52182;
    wire N__52181;
    wire N__52178;
    wire N__52175;
    wire N__52170;
    wire N__52167;
    wire N__52164;
    wire N__52161;
    wire N__52158;
    wire N__52155;
    wire N__52152;
    wire N__52149;
    wire N__52148;
    wire N__52145;
    wire N__52142;
    wire N__52139;
    wire N__52138;
    wire N__52135;
    wire N__52132;
    wire N__52129;
    wire N__52124;
    wire N__52119;
    wire N__52116;
    wire N__52113;
    wire N__52110;
    wire N__52109;
    wire N__52108;
    wire N__52105;
    wire N__52100;
    wire N__52095;
    wire N__52092;
    wire N__52091;
    wire N__52090;
    wire N__52087;
    wire N__52082;
    wire N__52079;
    wire N__52076;
    wire N__52071;
    wire N__52068;
    wire N__52065;
    wire N__52062;
    wire N__52059;
    wire N__52056;
    wire N__52053;
    wire N__52050;
    wire N__52047;
    wire N__52046;
    wire N__52045;
    wire N__52042;
    wire N__52037;
    wire N__52032;
    wire N__52031;
    wire N__52030;
    wire N__52029;
    wire N__52020;
    wire N__52017;
    wire N__52014;
    wire N__52013;
    wire N__52012;
    wire N__52009;
    wire N__52004;
    wire N__51999;
    wire N__51996;
    wire N__51993;
    wire N__51990;
    wire N__51987;
    wire N__51984;
    wire N__51981;
    wire N__51978;
    wire N__51975;
    wire N__51972;
    wire N__51969;
    wire N__51966;
    wire N__51963;
    wire N__51962;
    wire N__51959;
    wire N__51956;
    wire N__51951;
    wire N__51948;
    wire N__51945;
    wire N__51942;
    wire N__51939;
    wire N__51936;
    wire N__51933;
    wire N__51930;
    wire N__51927;
    wire N__51926;
    wire N__51923;
    wire N__51920;
    wire N__51919;
    wire N__51916;
    wire N__51915;
    wire N__51910;
    wire N__51907;
    wire N__51904;
    wire N__51901;
    wire N__51896;
    wire N__51891;
    wire N__51888;
    wire N__51885;
    wire N__51882;
    wire N__51879;
    wire N__51878;
    wire N__51875;
    wire N__51872;
    wire N__51867;
    wire N__51864;
    wire N__51861;
    wire N__51858;
    wire N__51855;
    wire N__51852;
    wire N__51849;
    wire N__51846;
    wire N__51843;
    wire N__51840;
    wire N__51837;
    wire N__51836;
    wire N__51833;
    wire N__51830;
    wire N__51827;
    wire N__51822;
    wire N__51819;
    wire N__51816;
    wire N__51813;
    wire N__51812;
    wire N__51809;
    wire N__51806;
    wire N__51801;
    wire N__51798;
    wire N__51795;
    wire N__51792;
    wire N__51791;
    wire N__51788;
    wire N__51785;
    wire N__51780;
    wire N__51777;
    wire N__51774;
    wire N__51771;
    wire N__51768;
    wire N__51767;
    wire N__51762;
    wire N__51759;
    wire N__51756;
    wire N__51753;
    wire N__51750;
    wire N__51747;
    wire N__51746;
    wire N__51741;
    wire N__51738;
    wire N__51737;
    wire N__51732;
    wire N__51729;
    wire N__51726;
    wire N__51723;
    wire N__51720;
    wire N__51719;
    wire N__51716;
    wire N__51713;
    wire N__51710;
    wire N__51707;
    wire N__51704;
    wire N__51701;
    wire N__51696;
    wire N__51693;
    wire N__51692;
    wire N__51689;
    wire N__51686;
    wire N__51681;
    wire N__51680;
    wire N__51675;
    wire N__51672;
    wire N__51669;
    wire N__51666;
    wire N__51663;
    wire N__51660;
    wire N__51659;
    wire N__51654;
    wire N__51651;
    wire N__51650;
    wire N__51645;
    wire N__51642;
    wire N__51639;
    wire N__51636;
    wire N__51633;
    wire N__51632;
    wire N__51627;
    wire N__51624;
    wire N__51623;
    wire N__51618;
    wire N__51615;
    wire N__51612;
    wire N__51609;
    wire N__51606;
    wire N__51605;
    wire N__51602;
    wire N__51599;
    wire N__51596;
    wire N__51593;
    wire N__51590;
    wire N__51587;
    wire N__51584;
    wire N__51581;
    wire N__51576;
    wire N__51575;
    wire N__51570;
    wire N__51567;
    wire N__51564;
    wire N__51561;
    wire N__51558;
    wire N__51555;
    wire N__51554;
    wire N__51553;
    wire N__51548;
    wire N__51545;
    wire N__51542;
    wire N__51539;
    wire N__51536;
    wire N__51533;
    wire N__51530;
    wire N__51525;
    wire N__51522;
    wire N__51519;
    wire N__51516;
    wire N__51513;
    wire N__51510;
    wire N__51509;
    wire N__51506;
    wire N__51503;
    wire N__51500;
    wire N__51495;
    wire N__51494;
    wire N__51493;
    wire N__51492;
    wire N__51491;
    wire N__51490;
    wire N__51489;
    wire N__51488;
    wire N__51487;
    wire N__51486;
    wire N__51485;
    wire N__51484;
    wire N__51483;
    wire N__51482;
    wire N__51481;
    wire N__51480;
    wire N__51479;
    wire N__51478;
    wire N__51477;
    wire N__51476;
    wire N__51475;
    wire N__51474;
    wire N__51473;
    wire N__51472;
    wire N__51423;
    wire N__51420;
    wire N__51417;
    wire N__51414;
    wire N__51411;
    wire N__51408;
    wire N__51405;
    wire N__51402;
    wire N__51399;
    wire N__51396;
    wire N__51393;
    wire N__51390;
    wire N__51387;
    wire N__51384;
    wire N__51381;
    wire N__51378;
    wire N__51375;
    wire N__51372;
    wire N__51371;
    wire N__51368;
    wire N__51365;
    wire N__51362;
    wire N__51359;
    wire N__51356;
    wire N__51353;
    wire N__51348;
    wire N__51347;
    wire N__51342;
    wire N__51339;
    wire N__51336;
    wire N__51333;
    wire N__51330;
    wire N__51327;
    wire N__51324;
    wire N__51321;
    wire N__51318;
    wire N__51315;
    wire N__51314;
    wire N__51311;
    wire N__51308;
    wire N__51305;
    wire N__51302;
    wire N__51299;
    wire N__51296;
    wire N__51291;
    wire N__51288;
    wire N__51285;
    wire N__51284;
    wire N__51281;
    wire N__51278;
    wire N__51275;
    wire N__51272;
    wire N__51269;
    wire N__51266;
    wire N__51263;
    wire N__51260;
    wire N__51257;
    wire N__51254;
    wire N__51249;
    wire N__51246;
    wire N__51243;
    wire N__51242;
    wire N__51239;
    wire N__51236;
    wire N__51233;
    wire N__51230;
    wire N__51227;
    wire N__51224;
    wire N__51221;
    wire N__51218;
    wire N__51213;
    wire N__51210;
    wire N__51209;
    wire N__51206;
    wire N__51203;
    wire N__51200;
    wire N__51197;
    wire N__51194;
    wire N__51191;
    wire N__51186;
    wire N__51183;
    wire N__51180;
    wire N__51179;
    wire N__51176;
    wire N__51173;
    wire N__51168;
    wire N__51167;
    wire N__51166;
    wire N__51161;
    wire N__51158;
    wire N__51157;
    wire N__51156;
    wire N__51155;
    wire N__51154;
    wire N__51151;
    wire N__51148;
    wire N__51143;
    wire N__51138;
    wire N__51135;
    wire N__51128;
    wire N__51123;
    wire N__51120;
    wire N__51117;
    wire N__51114;
    wire N__51113;
    wire N__51112;
    wire N__51109;
    wire N__51106;
    wire N__51103;
    wire N__51098;
    wire N__51093;
    wire N__51090;
    wire N__51087;
    wire N__51084;
    wire N__51081;
    wire N__51078;
    wire N__51077;
    wire N__51074;
    wire N__51073;
    wire N__51068;
    wire N__51065;
    wire N__51062;
    wire N__51057;
    wire N__51054;
    wire N__51051;
    wire N__51048;
    wire N__51045;
    wire N__51042;
    wire N__51041;
    wire N__51040;
    wire N__51037;
    wire N__51032;
    wire N__51027;
    wire N__51024;
    wire N__51021;
    wire N__51018;
    wire N__51017;
    wire N__51016;
    wire N__51015;
    wire N__51010;
    wire N__51005;
    wire N__51000;
    wire N__50997;
    wire N__50994;
    wire N__50993;
    wire N__50992;
    wire N__50991;
    wire N__50990;
    wire N__50987;
    wire N__50986;
    wire N__50983;
    wire N__50978;
    wire N__50971;
    wire N__50964;
    wire N__50961;
    wire N__50960;
    wire N__50959;
    wire N__50958;
    wire N__50955;
    wire N__50948;
    wire N__50947;
    wire N__50946;
    wire N__50945;
    wire N__50944;
    wire N__50943;
    wire N__50942;
    wire N__50937;
    wire N__50936;
    wire N__50935;
    wire N__50930;
    wire N__50929;
    wire N__50928;
    wire N__50923;
    wire N__50918;
    wire N__50915;
    wire N__50910;
    wire N__50907;
    wire N__50904;
    wire N__50901;
    wire N__50886;
    wire N__50883;
    wire N__50880;
    wire N__50877;
    wire N__50874;
    wire N__50873;
    wire N__50868;
    wire N__50865;
    wire N__50862;
    wire N__50859;
    wire N__50858;
    wire N__50857;
    wire N__50854;
    wire N__50851;
    wire N__50848;
    wire N__50843;
    wire N__50838;
    wire N__50835;
    wire N__50834;
    wire N__50833;
    wire N__50832;
    wire N__50829;
    wire N__50824;
    wire N__50823;
    wire N__50820;
    wire N__50815;
    wire N__50814;
    wire N__50813;
    wire N__50812;
    wire N__50809;
    wire N__50806;
    wire N__50803;
    wire N__50796;
    wire N__50787;
    wire N__50786;
    wire N__50785;
    wire N__50784;
    wire N__50783;
    wire N__50782;
    wire N__50779;
    wire N__50774;
    wire N__50771;
    wire N__50770;
    wire N__50769;
    wire N__50764;
    wire N__50759;
    wire N__50758;
    wire N__50755;
    wire N__50750;
    wire N__50747;
    wire N__50744;
    wire N__50741;
    wire N__50736;
    wire N__50731;
    wire N__50724;
    wire N__50721;
    wire N__50718;
    wire N__50717;
    wire N__50714;
    wire N__50711;
    wire N__50706;
    wire N__50703;
    wire N__50702;
    wire N__50699;
    wire N__50696;
    wire N__50693;
    wire N__50690;
    wire N__50687;
    wire N__50684;
    wire N__50679;
    wire N__50676;
    wire N__50675;
    wire N__50672;
    wire N__50669;
    wire N__50666;
    wire N__50663;
    wire N__50660;
    wire N__50657;
    wire N__50652;
    wire N__50649;
    wire N__50646;
    wire N__50643;
    wire N__50640;
    wire N__50637;
    wire N__50634;
    wire N__50631;
    wire N__50628;
    wire N__50625;
    wire N__50622;
    wire N__50619;
    wire N__50616;
    wire N__50613;
    wire N__50610;
    wire N__50607;
    wire N__50604;
    wire N__50601;
    wire N__50598;
    wire N__50595;
    wire N__50592;
    wire N__50589;
    wire N__50586;
    wire N__50583;
    wire N__50580;
    wire N__50577;
    wire N__50574;
    wire N__50573;
    wire N__50570;
    wire N__50567;
    wire N__50564;
    wire N__50561;
    wire N__50556;
    wire N__50555;
    wire N__50552;
    wire N__50549;
    wire N__50546;
    wire N__50543;
    wire N__50538;
    wire N__50535;
    wire N__50532;
    wire N__50529;
    wire N__50526;
    wire N__50523;
    wire N__50522;
    wire N__50521;
    wire N__50518;
    wire N__50515;
    wire N__50512;
    wire N__50505;
    wire N__50502;
    wire N__50499;
    wire N__50498;
    wire N__50495;
    wire N__50492;
    wire N__50489;
    wire N__50484;
    wire N__50483;
    wire N__50480;
    wire N__50477;
    wire N__50474;
    wire N__50473;
    wire N__50470;
    wire N__50467;
    wire N__50464;
    wire N__50457;
    wire N__50454;
    wire N__50451;
    wire N__50448;
    wire N__50445;
    wire N__50444;
    wire N__50443;
    wire N__50440;
    wire N__50437;
    wire N__50436;
    wire N__50433;
    wire N__50428;
    wire N__50425;
    wire N__50422;
    wire N__50419;
    wire N__50416;
    wire N__50413;
    wire N__50408;
    wire N__50403;
    wire N__50400;
    wire N__50397;
    wire N__50394;
    wire N__50391;
    wire N__50388;
    wire N__50385;
    wire N__50382;
    wire N__50379;
    wire N__50376;
    wire N__50373;
    wire N__50370;
    wire N__50367;
    wire N__50364;
    wire N__50361;
    wire N__50360;
    wire N__50357;
    wire N__50354;
    wire N__50349;
    wire N__50346;
    wire N__50343;
    wire N__50340;
    wire N__50337;
    wire N__50334;
    wire N__50331;
    wire N__50328;
    wire N__50325;
    wire N__50322;
    wire N__50319;
    wire N__50316;
    wire N__50315;
    wire N__50312;
    wire N__50309;
    wire N__50304;
    wire N__50301;
    wire N__50298;
    wire N__50295;
    wire N__50292;
    wire N__50289;
    wire N__50286;
    wire N__50283;
    wire N__50280;
    wire N__50277;
    wire N__50276;
    wire N__50273;
    wire N__50270;
    wire N__50265;
    wire N__50262;
    wire N__50261;
    wire N__50256;
    wire N__50253;
    wire N__50250;
    wire N__50247;
    wire N__50244;
    wire N__50241;
    wire N__50240;
    wire N__50237;
    wire N__50234;
    wire N__50231;
    wire N__50230;
    wire N__50229;
    wire N__50226;
    wire N__50223;
    wire N__50220;
    wire N__50217;
    wire N__50208;
    wire N__50205;
    wire N__50202;
    wire N__50199;
    wire N__50196;
    wire N__50193;
    wire N__50190;
    wire N__50187;
    wire N__50184;
    wire N__50181;
    wire N__50178;
    wire N__50177;
    wire N__50174;
    wire N__50171;
    wire N__50168;
    wire N__50165;
    wire N__50160;
    wire N__50159;
    wire N__50158;
    wire N__50155;
    wire N__50154;
    wire N__50153;
    wire N__50150;
    wire N__50147;
    wire N__50146;
    wire N__50143;
    wire N__50140;
    wire N__50137;
    wire N__50134;
    wire N__50131;
    wire N__50128;
    wire N__50125;
    wire N__50122;
    wire N__50119;
    wire N__50116;
    wire N__50113;
    wire N__50108;
    wire N__50103;
    wire N__50100;
    wire N__50095;
    wire N__50092;
    wire N__50085;
    wire N__50082;
    wire N__50079;
    wire N__50076;
    wire N__50073;
    wire N__50070;
    wire N__50067;
    wire N__50064;
    wire N__50061;
    wire N__50058;
    wire N__50055;
    wire N__50052;
    wire N__50049;
    wire N__50046;
    wire N__50043;
    wire N__50040;
    wire N__50037;
    wire N__50034;
    wire N__50031;
    wire N__50028;
    wire N__50025;
    wire N__50022;
    wire N__50019;
    wire N__50016;
    wire N__50013;
    wire N__50010;
    wire N__50007;
    wire N__50004;
    wire N__50001;
    wire N__49998;
    wire N__49995;
    wire N__49992;
    wire N__49991;
    wire N__49988;
    wire N__49985;
    wire N__49980;
    wire N__49979;
    wire N__49976;
    wire N__49973;
    wire N__49968;
    wire N__49967;
    wire N__49962;
    wire N__49959;
    wire N__49956;
    wire N__49955;
    wire N__49950;
    wire N__49947;
    wire N__49944;
    wire N__49941;
    wire N__49938;
    wire N__49935;
    wire N__49932;
    wire N__49929;
    wire N__49926;
    wire N__49923;
    wire N__49920;
    wire N__49917;
    wire N__49914;
    wire N__49911;
    wire N__49908;
    wire N__49905;
    wire N__49902;
    wire N__49899;
    wire N__49896;
    wire N__49893;
    wire N__49890;
    wire N__49887;
    wire N__49884;
    wire N__49881;
    wire N__49878;
    wire N__49875;
    wire N__49872;
    wire N__49869;
    wire N__49866;
    wire N__49863;
    wire N__49860;
    wire N__49857;
    wire N__49854;
    wire N__49851;
    wire N__49848;
    wire N__49845;
    wire N__49842;
    wire N__49839;
    wire N__49836;
    wire N__49833;
    wire N__49830;
    wire N__49827;
    wire N__49824;
    wire N__49821;
    wire N__49818;
    wire N__49815;
    wire N__49812;
    wire N__49809;
    wire N__49806;
    wire N__49803;
    wire N__49800;
    wire N__49797;
    wire N__49794;
    wire N__49791;
    wire N__49788;
    wire N__49785;
    wire N__49782;
    wire N__49779;
    wire N__49778;
    wire N__49777;
    wire N__49776;
    wire N__49771;
    wire N__49766;
    wire N__49763;
    wire N__49760;
    wire N__49757;
    wire N__49752;
    wire N__49749;
    wire N__49746;
    wire N__49743;
    wire N__49740;
    wire N__49737;
    wire N__49734;
    wire N__49731;
    wire N__49730;
    wire N__49729;
    wire N__49728;
    wire N__49725;
    wire N__49718;
    wire N__49713;
    wire N__49710;
    wire N__49707;
    wire N__49704;
    wire N__49701;
    wire N__49698;
    wire N__49695;
    wire N__49692;
    wire N__49689;
    wire N__49688;
    wire N__49687;
    wire N__49686;
    wire N__49683;
    wire N__49678;
    wire N__49675;
    wire N__49670;
    wire N__49667;
    wire N__49664;
    wire N__49661;
    wire N__49656;
    wire N__49653;
    wire N__49652;
    wire N__49649;
    wire N__49646;
    wire N__49643;
    wire N__49640;
    wire N__49635;
    wire N__49632;
    wire N__49629;
    wire N__49628;
    wire N__49627;
    wire N__49626;
    wire N__49625;
    wire N__49624;
    wire N__49623;
    wire N__49622;
    wire N__49621;
    wire N__49616;
    wire N__49611;
    wire N__49608;
    wire N__49607;
    wire N__49604;
    wire N__49597;
    wire N__49592;
    wire N__49589;
    wire N__49586;
    wire N__49581;
    wire N__49576;
    wire N__49569;
    wire N__49566;
    wire N__49563;
    wire N__49560;
    wire N__49557;
    wire N__49554;
    wire N__49551;
    wire N__49548;
    wire N__49547;
    wire N__49544;
    wire N__49541;
    wire N__49536;
    wire N__49533;
    wire N__49530;
    wire N__49527;
    wire N__49524;
    wire N__49521;
    wire N__49518;
    wire N__49515;
    wire N__49512;
    wire N__49511;
    wire N__49508;
    wire N__49507;
    wire N__49504;
    wire N__49501;
    wire N__49496;
    wire N__49491;
    wire N__49488;
    wire N__49485;
    wire N__49482;
    wire N__49479;
    wire N__49478;
    wire N__49475;
    wire N__49474;
    wire N__49471;
    wire N__49468;
    wire N__49465;
    wire N__49464;
    wire N__49461;
    wire N__49456;
    wire N__49453;
    wire N__49450;
    wire N__49443;
    wire N__49440;
    wire N__49439;
    wire N__49438;
    wire N__49435;
    wire N__49432;
    wire N__49429;
    wire N__49422;
    wire N__49419;
    wire N__49416;
    wire N__49415;
    wire N__49412;
    wire N__49409;
    wire N__49404;
    wire N__49401;
    wire N__49398;
    wire N__49395;
    wire N__49392;
    wire N__49389;
    wire N__49386;
    wire N__49383;
    wire N__49380;
    wire N__49377;
    wire N__49376;
    wire N__49373;
    wire N__49370;
    wire N__49367;
    wire N__49364;
    wire N__49359;
    wire N__49358;
    wire N__49355;
    wire N__49352;
    wire N__49351;
    wire N__49348;
    wire N__49345;
    wire N__49342;
    wire N__49341;
    wire N__49338;
    wire N__49335;
    wire N__49332;
    wire N__49329;
    wire N__49328;
    wire N__49325;
    wire N__49322;
    wire N__49319;
    wire N__49316;
    wire N__49313;
    wire N__49302;
    wire N__49299;
    wire N__49298;
    wire N__49293;
    wire N__49290;
    wire N__49287;
    wire N__49286;
    wire N__49281;
    wire N__49278;
    wire N__49275;
    wire N__49272;
    wire N__49269;
    wire N__49266;
    wire N__49263;
    wire N__49262;
    wire N__49257;
    wire N__49254;
    wire N__49251;
    wire N__49248;
    wire N__49247;
    wire N__49246;
    wire N__49245;
    wire N__49240;
    wire N__49237;
    wire N__49234;
    wire N__49231;
    wire N__49224;
    wire N__49223;
    wire N__49220;
    wire N__49217;
    wire N__49216;
    wire N__49215;
    wire N__49212;
    wire N__49209;
    wire N__49204;
    wire N__49203;
    wire N__49200;
    wire N__49197;
    wire N__49194;
    wire N__49191;
    wire N__49182;
    wire N__49181;
    wire N__49178;
    wire N__49177;
    wire N__49174;
    wire N__49171;
    wire N__49168;
    wire N__49167;
    wire N__49164;
    wire N__49161;
    wire N__49158;
    wire N__49155;
    wire N__49154;
    wire N__49147;
    wire N__49142;
    wire N__49137;
    wire N__49136;
    wire N__49133;
    wire N__49130;
    wire N__49129;
    wire N__49128;
    wire N__49125;
    wire N__49122;
    wire N__49119;
    wire N__49118;
    wire N__49115;
    wire N__49108;
    wire N__49105;
    wire N__49102;
    wire N__49099;
    wire N__49096;
    wire N__49091;
    wire N__49088;
    wire N__49085;
    wire N__49082;
    wire N__49079;
    wire N__49074;
    wire N__49071;
    wire N__49068;
    wire N__49065;
    wire N__49062;
    wire N__49059;
    wire N__49056;
    wire N__49053;
    wire N__49052;
    wire N__49051;
    wire N__49044;
    wire N__49041;
    wire N__49038;
    wire N__49035;
    wire N__49032;
    wire N__49029;
    wire N__49026;
    wire N__49023;
    wire N__49022;
    wire N__49021;
    wire N__49020;
    wire N__49019;
    wire N__49016;
    wire N__49009;
    wire N__49006;
    wire N__49001;
    wire N__48996;
    wire N__48993;
    wire N__48990;
    wire N__48987;
    wire N__48984;
    wire N__48981;
    wire N__48978;
    wire N__48975;
    wire N__48972;
    wire N__48971;
    wire N__48970;
    wire N__48969;
    wire N__48968;
    wire N__48967;
    wire N__48964;
    wire N__48963;
    wire N__48960;
    wire N__48955;
    wire N__48950;
    wire N__48945;
    wire N__48942;
    wire N__48939;
    wire N__48934;
    wire N__48931;
    wire N__48926;
    wire N__48923;
    wire N__48920;
    wire N__48915;
    wire N__48912;
    wire N__48909;
    wire N__48908;
    wire N__48907;
    wire N__48906;
    wire N__48903;
    wire N__48900;
    wire N__48897;
    wire N__48894;
    wire N__48885;
    wire N__48884;
    wire N__48883;
    wire N__48882;
    wire N__48881;
    wire N__48880;
    wire N__48879;
    wire N__48876;
    wire N__48869;
    wire N__48866;
    wire N__48861;
    wire N__48858;
    wire N__48853;
    wire N__48850;
    wire N__48845;
    wire N__48842;
    wire N__48839;
    wire N__48836;
    wire N__48833;
    wire N__48830;
    wire N__48827;
    wire N__48822;
    wire N__48821;
    wire N__48820;
    wire N__48817;
    wire N__48816;
    wire N__48815;
    wire N__48814;
    wire N__48809;
    wire N__48802;
    wire N__48799;
    wire N__48796;
    wire N__48795;
    wire N__48790;
    wire N__48787;
    wire N__48784;
    wire N__48781;
    wire N__48774;
    wire N__48773;
    wire N__48772;
    wire N__48771;
    wire N__48770;
    wire N__48769;
    wire N__48768;
    wire N__48767;
    wire N__48762;
    wire N__48755;
    wire N__48752;
    wire N__48747;
    wire N__48740;
    wire N__48735;
    wire N__48732;
    wire N__48729;
    wire N__48726;
    wire N__48723;
    wire N__48720;
    wire N__48717;
    wire N__48714;
    wire N__48711;
    wire N__48708;
    wire N__48705;
    wire N__48702;
    wire N__48699;
    wire N__48696;
    wire N__48695;
    wire N__48692;
    wire N__48689;
    wire N__48686;
    wire N__48683;
    wire N__48680;
    wire N__48677;
    wire N__48672;
    wire N__48671;
    wire N__48668;
    wire N__48667;
    wire N__48664;
    wire N__48659;
    wire N__48658;
    wire N__48657;
    wire N__48654;
    wire N__48653;
    wire N__48652;
    wire N__48649;
    wire N__48646;
    wire N__48645;
    wire N__48642;
    wire N__48639;
    wire N__48634;
    wire N__48631;
    wire N__48626;
    wire N__48615;
    wire N__48614;
    wire N__48611;
    wire N__48608;
    wire N__48605;
    wire N__48600;
    wire N__48597;
    wire N__48594;
    wire N__48593;
    wire N__48588;
    wire N__48585;
    wire N__48582;
    wire N__48581;
    wire N__48576;
    wire N__48573;
    wire N__48570;
    wire N__48569;
    wire N__48568;
    wire N__48567;
    wire N__48564;
    wire N__48557;
    wire N__48552;
    wire N__48549;
    wire N__48548;
    wire N__48547;
    wire N__48542;
    wire N__48539;
    wire N__48536;
    wire N__48533;
    wire N__48528;
    wire N__48525;
    wire N__48524;
    wire N__48523;
    wire N__48522;
    wire N__48519;
    wire N__48514;
    wire N__48511;
    wire N__48508;
    wire N__48505;
    wire N__48498;
    wire N__48495;
    wire N__48492;
    wire N__48489;
    wire N__48486;
    wire N__48483;
    wire N__48480;
    wire N__48477;
    wire N__48474;
    wire N__48471;
    wire N__48468;
    wire N__48465;
    wire N__48462;
    wire N__48459;
    wire N__48458;
    wire N__48457;
    wire N__48454;
    wire N__48449;
    wire N__48448;
    wire N__48443;
    wire N__48440;
    wire N__48435;
    wire N__48432;
    wire N__48429;
    wire N__48428;
    wire N__48427;
    wire N__48426;
    wire N__48425;
    wire N__48424;
    wire N__48421;
    wire N__48410;
    wire N__48405;
    wire N__48402;
    wire N__48399;
    wire N__48398;
    wire N__48395;
    wire N__48392;
    wire N__48389;
    wire N__48384;
    wire N__48381;
    wire N__48378;
    wire N__48375;
    wire N__48372;
    wire N__48369;
    wire N__48368;
    wire N__48367;
    wire N__48364;
    wire N__48359;
    wire N__48354;
    wire N__48351;
    wire N__48350;
    wire N__48347;
    wire N__48344;
    wire N__48339;
    wire N__48338;
    wire N__48337;
    wire N__48336;
    wire N__48335;
    wire N__48334;
    wire N__48327;
    wire N__48324;
    wire N__48321;
    wire N__48320;
    wire N__48319;
    wire N__48318;
    wire N__48315;
    wire N__48314;
    wire N__48313;
    wire N__48312;
    wire N__48311;
    wire N__48310;
    wire N__48309;
    wire N__48304;
    wire N__48295;
    wire N__48288;
    wire N__48283;
    wire N__48278;
    wire N__48275;
    wire N__48270;
    wire N__48265;
    wire N__48262;
    wire N__48257;
    wire N__48254;
    wire N__48251;
    wire N__48248;
    wire N__48245;
    wire N__48240;
    wire N__48237;
    wire N__48236;
    wire N__48231;
    wire N__48228;
    wire N__48227;
    wire N__48222;
    wire N__48219;
    wire N__48216;
    wire N__48213;
    wire N__48210;
    wire N__48207;
    wire N__48206;
    wire N__48201;
    wire N__48198;
    wire N__48195;
    wire N__48192;
    wire N__48189;
    wire N__48186;
    wire N__48183;
    wire N__48180;
    wire N__48177;
    wire N__48176;
    wire N__48171;
    wire N__48168;
    wire N__48167;
    wire N__48164;
    wire N__48161;
    wire N__48158;
    wire N__48155;
    wire N__48150;
    wire N__48147;
    wire N__48144;
    wire N__48141;
    wire N__48138;
    wire N__48135;
    wire N__48132;
    wire N__48129;
    wire N__48126;
    wire N__48123;
    wire N__48120;
    wire N__48119;
    wire N__48114;
    wire N__48111;
    wire N__48108;
    wire N__48105;
    wire N__48102;
    wire N__48101;
    wire N__48100;
    wire N__48095;
    wire N__48092;
    wire N__48087;
    wire N__48084;
    wire N__48083;
    wire N__48078;
    wire N__48075;
    wire N__48072;
    wire N__48069;
    wire N__48066;
    wire N__48063;
    wire N__48060;
    wire N__48059;
    wire N__48056;
    wire N__48053;
    wire N__48050;
    wire N__48047;
    wire N__48042;
    wire N__48041;
    wire N__48038;
    wire N__48037;
    wire N__48034;
    wire N__48029;
    wire N__48024;
    wire N__48021;
    wire N__48018;
    wire N__48017;
    wire N__48014;
    wire N__48011;
    wire N__48008;
    wire N__48005;
    wire N__48002;
    wire N__47997;
    wire N__47996;
    wire N__47993;
    wire N__47992;
    wire N__47991;
    wire N__47990;
    wire N__47989;
    wire N__47988;
    wire N__47987;
    wire N__47986;
    wire N__47983;
    wire N__47982;
    wire N__47979;
    wire N__47978;
    wire N__47961;
    wire N__47958;
    wire N__47955;
    wire N__47952;
    wire N__47951;
    wire N__47950;
    wire N__47947;
    wire N__47944;
    wire N__47943;
    wire N__47940;
    wire N__47935;
    wire N__47932;
    wire N__47929;
    wire N__47926;
    wire N__47923;
    wire N__47920;
    wire N__47909;
    wire N__47904;
    wire N__47901;
    wire N__47898;
    wire N__47895;
    wire N__47894;
    wire N__47893;
    wire N__47890;
    wire N__47885;
    wire N__47880;
    wire N__47877;
    wire N__47876;
    wire N__47875;
    wire N__47874;
    wire N__47865;
    wire N__47862;
    wire N__47861;
    wire N__47860;
    wire N__47857;
    wire N__47854;
    wire N__47851;
    wire N__47850;
    wire N__47849;
    wire N__47846;
    wire N__47839;
    wire N__47836;
    wire N__47829;
    wire N__47826;
    wire N__47823;
    wire N__47822;
    wire N__47817;
    wire N__47816;
    wire N__47813;
    wire N__47810;
    wire N__47805;
    wire N__47802;
    wire N__47799;
    wire N__47798;
    wire N__47795;
    wire N__47792;
    wire N__47789;
    wire N__47786;
    wire N__47781;
    wire N__47778;
    wire N__47775;
    wire N__47772;
    wire N__47769;
    wire N__47766;
    wire N__47763;
    wire N__47760;
    wire N__47757;
    wire N__47754;
    wire N__47751;
    wire N__47748;
    wire N__47745;
    wire N__47742;
    wire N__47739;
    wire N__47736;
    wire N__47733;
    wire N__47730;
    wire N__47727;
    wire N__47724;
    wire N__47721;
    wire N__47718;
    wire N__47717;
    wire N__47714;
    wire N__47711;
    wire N__47708;
    wire N__47703;
    wire N__47702;
    wire N__47699;
    wire N__47696;
    wire N__47693;
    wire N__47688;
    wire N__47687;
    wire N__47684;
    wire N__47681;
    wire N__47678;
    wire N__47673;
    wire N__47672;
    wire N__47669;
    wire N__47666;
    wire N__47663;
    wire N__47658;
    wire N__47657;
    wire N__47654;
    wire N__47651;
    wire N__47648;
    wire N__47643;
    wire N__47642;
    wire N__47639;
    wire N__47636;
    wire N__47633;
    wire N__47628;
    wire N__47625;
    wire N__47622;
    wire N__47619;
    wire N__47616;
    wire N__47613;
    wire N__47610;
    wire N__47607;
    wire N__47604;
    wire N__47601;
    wire N__47598;
    wire N__47595;
    wire N__47592;
    wire N__47589;
    wire N__47588;
    wire N__47587;
    wire N__47586;
    wire N__47585;
    wire N__47584;
    wire N__47583;
    wire N__47582;
    wire N__47565;
    wire N__47562;
    wire N__47559;
    wire N__47556;
    wire N__47553;
    wire N__47550;
    wire N__47547;
    wire N__47544;
    wire N__47541;
    wire N__47540;
    wire N__47537;
    wire N__47534;
    wire N__47529;
    wire N__47528;
    wire N__47525;
    wire N__47522;
    wire N__47519;
    wire N__47514;
    wire N__47511;
    wire N__47508;
    wire N__47505;
    wire N__47502;
    wire N__47499;
    wire N__47496;
    wire N__47493;
    wire N__47490;
    wire N__47487;
    wire N__47484;
    wire N__47481;
    wire N__47478;
    wire N__47475;
    wire N__47472;
    wire N__47469;
    wire N__47466;
    wire N__47463;
    wire N__47460;
    wire N__47457;
    wire N__47454;
    wire N__47451;
    wire N__47448;
    wire N__47445;
    wire N__47442;
    wire N__47441;
    wire N__47438;
    wire N__47437;
    wire N__47434;
    wire N__47431;
    wire N__47428;
    wire N__47425;
    wire N__47422;
    wire N__47415;
    wire N__47414;
    wire N__47411;
    wire N__47408;
    wire N__47407;
    wire N__47404;
    wire N__47401;
    wire N__47398;
    wire N__47395;
    wire N__47388;
    wire N__47387;
    wire N__47384;
    wire N__47383;
    wire N__47380;
    wire N__47377;
    wire N__47374;
    wire N__47371;
    wire N__47368;
    wire N__47361;
    wire N__47358;
    wire N__47355;
    wire N__47352;
    wire N__47349;
    wire N__47346;
    wire N__47343;
    wire N__47340;
    wire N__47337;
    wire N__47334;
    wire N__47331;
    wire N__47328;
    wire N__47325;
    wire N__47322;
    wire N__47319;
    wire N__47316;
    wire N__47313;
    wire N__47312;
    wire N__47309;
    wire N__47306;
    wire N__47301;
    wire N__47298;
    wire N__47295;
    wire N__47292;
    wire N__47289;
    wire N__47286;
    wire N__47285;
    wire N__47284;
    wire N__47281;
    wire N__47278;
    wire N__47275;
    wire N__47272;
    wire N__47265;
    wire N__47262;
    wire N__47259;
    wire N__47258;
    wire N__47255;
    wire N__47252;
    wire N__47249;
    wire N__47246;
    wire N__47241;
    wire N__47238;
    wire N__47235;
    wire N__47232;
    wire N__47229;
    wire N__47228;
    wire N__47225;
    wire N__47224;
    wire N__47221;
    wire N__47218;
    wire N__47213;
    wire N__47208;
    wire N__47205;
    wire N__47202;
    wire N__47199;
    wire N__47196;
    wire N__47193;
    wire N__47190;
    wire N__47189;
    wire N__47188;
    wire N__47185;
    wire N__47182;
    wire N__47179;
    wire N__47174;
    wire N__47171;
    wire N__47168;
    wire N__47163;
    wire N__47160;
    wire N__47159;
    wire N__47158;
    wire N__47155;
    wire N__47152;
    wire N__47149;
    wire N__47146;
    wire N__47139;
    wire N__47136;
    wire N__47135;
    wire N__47132;
    wire N__47129;
    wire N__47124;
    wire N__47121;
    wire N__47118;
    wire N__47117;
    wire N__47116;
    wire N__47113;
    wire N__47108;
    wire N__47105;
    wire N__47100;
    wire N__47097;
    wire N__47094;
    wire N__47093;
    wire N__47092;
    wire N__47089;
    wire N__47084;
    wire N__47081;
    wire N__47076;
    wire N__47073;
    wire N__47070;
    wire N__47067;
    wire N__47064;
    wire N__47061;
    wire N__47058;
    wire N__47055;
    wire N__47052;
    wire N__47049;
    wire N__47046;
    wire N__47043;
    wire N__47040;
    wire N__47037;
    wire N__47034;
    wire N__47031;
    wire N__47028;
    wire N__47025;
    wire N__47022;
    wire N__47019;
    wire N__47016;
    wire N__47013;
    wire N__47010;
    wire N__47007;
    wire N__47004;
    wire N__47001;
    wire N__46998;
    wire N__46995;
    wire N__46992;
    wire N__46989;
    wire N__46986;
    wire N__46983;
    wire N__46980;
    wire N__46977;
    wire N__46974;
    wire N__46971;
    wire N__46968;
    wire N__46965;
    wire N__46962;
    wire N__46959;
    wire N__46956;
    wire N__46953;
    wire N__46950;
    wire N__46947;
    wire N__46944;
    wire N__46941;
    wire N__46938;
    wire N__46935;
    wire N__46932;
    wire N__46929;
    wire N__46926;
    wire N__46923;
    wire N__46920;
    wire N__46917;
    wire N__46914;
    wire N__46911;
    wire N__46908;
    wire N__46905;
    wire N__46902;
    wire N__46899;
    wire N__46896;
    wire N__46893;
    wire N__46890;
    wire N__46887;
    wire N__46884;
    wire N__46881;
    wire N__46878;
    wire N__46875;
    wire N__46872;
    wire N__46869;
    wire N__46866;
    wire N__46863;
    wire N__46860;
    wire N__46857;
    wire N__46854;
    wire N__46851;
    wire N__46848;
    wire N__46845;
    wire N__46842;
    wire N__46839;
    wire N__46836;
    wire N__46833;
    wire N__46830;
    wire N__46827;
    wire N__46824;
    wire N__46821;
    wire N__46818;
    wire N__46815;
    wire N__46812;
    wire N__46809;
    wire N__46806;
    wire N__46803;
    wire N__46800;
    wire N__46797;
    wire N__46794;
    wire N__46791;
    wire N__46788;
    wire N__46785;
    wire N__46782;
    wire N__46779;
    wire N__46776;
    wire N__46773;
    wire N__46770;
    wire N__46767;
    wire N__46764;
    wire N__46761;
    wire N__46758;
    wire N__46755;
    wire N__46754;
    wire N__46751;
    wire N__46748;
    wire N__46743;
    wire N__46740;
    wire N__46737;
    wire N__46734;
    wire N__46731;
    wire N__46728;
    wire N__46727;
    wire N__46724;
    wire N__46721;
    wire N__46716;
    wire N__46713;
    wire N__46710;
    wire N__46707;
    wire N__46704;
    wire N__46701;
    wire N__46698;
    wire N__46697;
    wire N__46696;
    wire N__46695;
    wire N__46694;
    wire N__46691;
    wire N__46682;
    wire N__46677;
    wire N__46674;
    wire N__46673;
    wire N__46672;
    wire N__46669;
    wire N__46666;
    wire N__46663;
    wire N__46662;
    wire N__46659;
    wire N__46652;
    wire N__46647;
    wire N__46644;
    wire N__46643;
    wire N__46638;
    wire N__46635;
    wire N__46632;
    wire N__46629;
    wire N__46626;
    wire N__46623;
    wire N__46620;
    wire N__46617;
    wire N__46614;
    wire N__46611;
    wire N__46608;
    wire N__46605;
    wire N__46602;
    wire N__46599;
    wire N__46596;
    wire N__46593;
    wire N__46590;
    wire N__46587;
    wire N__46584;
    wire N__46583;
    wire N__46582;
    wire N__46581;
    wire N__46578;
    wire N__46575;
    wire N__46570;
    wire N__46563;
    wire N__46560;
    wire N__46557;
    wire N__46554;
    wire N__46551;
    wire N__46548;
    wire N__46545;
    wire N__46542;
    wire N__46539;
    wire N__46536;
    wire N__46533;
    wire N__46532;
    wire N__46531;
    wire N__46528;
    wire N__46523;
    wire N__46520;
    wire N__46519;
    wire N__46516;
    wire N__46513;
    wire N__46510;
    wire N__46507;
    wire N__46500;
    wire N__46497;
    wire N__46496;
    wire N__46495;
    wire N__46492;
    wire N__46487;
    wire N__46486;
    wire N__46485;
    wire N__46484;
    wire N__46481;
    wire N__46478;
    wire N__46471;
    wire N__46464;
    wire N__46461;
    wire N__46460;
    wire N__46457;
    wire N__46454;
    wire N__46451;
    wire N__46446;
    wire N__46443;
    wire N__46440;
    wire N__46437;
    wire N__46434;
    wire N__46431;
    wire N__46428;
    wire N__46425;
    wire N__46422;
    wire N__46419;
    wire N__46416;
    wire N__46415;
    wire N__46412;
    wire N__46409;
    wire N__46404;
    wire N__46401;
    wire N__46400;
    wire N__46397;
    wire N__46394;
    wire N__46389;
    wire N__46386;
    wire N__46383;
    wire N__46380;
    wire N__46379;
    wire N__46378;
    wire N__46375;
    wire N__46372;
    wire N__46369;
    wire N__46362;
    wire N__46359;
    wire N__46356;
    wire N__46353;
    wire N__46350;
    wire N__46347;
    wire N__46344;
    wire N__46341;
    wire N__46340;
    wire N__46339;
    wire N__46338;
    wire N__46337;
    wire N__46336;
    wire N__46335;
    wire N__46334;
    wire N__46333;
    wire N__46332;
    wire N__46331;
    wire N__46328;
    wire N__46323;
    wire N__46322;
    wire N__46319;
    wire N__46316;
    wire N__46313;
    wire N__46312;
    wire N__46309;
    wire N__46306;
    wire N__46303;
    wire N__46300;
    wire N__46297;
    wire N__46294;
    wire N__46291;
    wire N__46282;
    wire N__46275;
    wire N__46268;
    wire N__46265;
    wire N__46262;
    wire N__46251;
    wire N__46250;
    wire N__46249;
    wire N__46242;
    wire N__46239;
    wire N__46236;
    wire N__46233;
    wire N__46230;
    wire N__46227;
    wire N__46224;
    wire N__46221;
    wire N__46218;
    wire N__46215;
    wire N__46212;
    wire N__46209;
    wire N__46206;
    wire N__46203;
    wire N__46200;
    wire N__46197;
    wire N__46194;
    wire N__46191;
    wire N__46188;
    wire N__46185;
    wire N__46182;
    wire N__46179;
    wire N__46176;
    wire N__46175;
    wire N__46170;
    wire N__46167;
    wire N__46164;
    wire N__46161;
    wire N__46158;
    wire N__46155;
    wire N__46152;
    wire N__46149;
    wire N__46148;
    wire N__46145;
    wire N__46142;
    wire N__46137;
    wire N__46134;
    wire N__46131;
    wire N__46128;
    wire N__46125;
    wire N__46122;
    wire N__46121;
    wire N__46116;
    wire N__46113;
    wire N__46110;
    wire N__46107;
    wire N__46104;
    wire N__46101;
    wire N__46098;
    wire N__46095;
    wire N__46092;
    wire N__46089;
    wire N__46086;
    wire N__46083;
    wire N__46080;
    wire N__46077;
    wire N__46074;
    wire N__46071;
    wire N__46068;
    wire N__46065;
    wire N__46062;
    wire N__46059;
    wire N__46056;
    wire N__46055;
    wire N__46052;
    wire N__46047;
    wire N__46044;
    wire N__46041;
    wire N__46038;
    wire N__46035;
    wire N__46032;
    wire N__46029;
    wire N__46026;
    wire N__46023;
    wire N__46022;
    wire N__46019;
    wire N__46016;
    wire N__46013;
    wire N__46008;
    wire N__46005;
    wire N__46002;
    wire N__45999;
    wire N__45996;
    wire N__45993;
    wire N__45992;
    wire N__45989;
    wire N__45986;
    wire N__45981;
    wire N__45978;
    wire N__45975;
    wire N__45974;
    wire N__45973;
    wire N__45970;
    wire N__45965;
    wire N__45960;
    wire N__45957;
    wire N__45954;
    wire N__45951;
    wire N__45948;
    wire N__45947;
    wire N__45944;
    wire N__45941;
    wire N__45936;
    wire N__45933;
    wire N__45930;
    wire N__45927;
    wire N__45924;
    wire N__45921;
    wire N__45918;
    wire N__45915;
    wire N__45914;
    wire N__45911;
    wire N__45908;
    wire N__45905;
    wire N__45902;
    wire N__45899;
    wire N__45896;
    wire N__45893;
    wire N__45890;
    wire N__45887;
    wire N__45884;
    wire N__45879;
    wire N__45876;
    wire N__45873;
    wire N__45872;
    wire N__45867;
    wire N__45864;
    wire N__45861;
    wire N__45858;
    wire N__45855;
    wire N__45852;
    wire N__45851;
    wire N__45848;
    wire N__45845;
    wire N__45840;
    wire N__45837;
    wire N__45834;
    wire N__45831;
    wire N__45828;
    wire N__45825;
    wire N__45822;
    wire N__45819;
    wire N__45816;
    wire N__45813;
    wire N__45810;
    wire N__45807;
    wire N__45804;
    wire N__45801;
    wire N__45800;
    wire N__45797;
    wire N__45794;
    wire N__45789;
    wire N__45788;
    wire N__45783;
    wire N__45780;
    wire N__45777;
    wire N__45774;
    wire N__45771;
    wire N__45770;
    wire N__45765;
    wire N__45762;
    wire N__45759;
    wire N__45756;
    wire N__45753;
    wire N__45750;
    wire N__45747;
    wire N__45744;
    wire N__45743;
    wire N__45740;
    wire N__45737;
    wire N__45732;
    wire N__45729;
    wire N__45726;
    wire N__45723;
    wire N__45720;
    wire N__45717;
    wire N__45714;
    wire N__45713;
    wire N__45710;
    wire N__45707;
    wire N__45702;
    wire N__45699;
    wire N__45698;
    wire N__45697;
    wire N__45694;
    wire N__45691;
    wire N__45690;
    wire N__45687;
    wire N__45684;
    wire N__45681;
    wire N__45678;
    wire N__45675;
    wire N__45672;
    wire N__45667;
    wire N__45664;
    wire N__45657;
    wire N__45656;
    wire N__45655;
    wire N__45654;
    wire N__45653;
    wire N__45650;
    wire N__45647;
    wire N__45644;
    wire N__45639;
    wire N__45638;
    wire N__45633;
    wire N__45628;
    wire N__45625;
    wire N__45622;
    wire N__45619;
    wire N__45616;
    wire N__45609;
    wire N__45608;
    wire N__45605;
    wire N__45602;
    wire N__45599;
    wire N__45598;
    wire N__45595;
    wire N__45592;
    wire N__45589;
    wire N__45588;
    wire N__45587;
    wire N__45584;
    wire N__45579;
    wire N__45574;
    wire N__45567;
    wire N__45564;
    wire N__45563;
    wire N__45560;
    wire N__45557;
    wire N__45552;
    wire N__45549;
    wire N__45548;
    wire N__45545;
    wire N__45542;
    wire N__45539;
    wire N__45536;
    wire N__45535;
    wire N__45532;
    wire N__45529;
    wire N__45526;
    wire N__45519;
    wire N__45518;
    wire N__45515;
    wire N__45512;
    wire N__45509;
    wire N__45506;
    wire N__45501;
    wire N__45500;
    wire N__45499;
    wire N__45496;
    wire N__45493;
    wire N__45490;
    wire N__45487;
    wire N__45482;
    wire N__45477;
    wire N__45476;
    wire N__45473;
    wire N__45470;
    wire N__45465;
    wire N__45462;
    wire N__45461;
    wire N__45460;
    wire N__45459;
    wire N__45458;
    wire N__45457;
    wire N__45456;
    wire N__45455;
    wire N__45454;
    wire N__45453;
    wire N__45450;
    wire N__45447;
    wire N__45446;
    wire N__45445;
    wire N__45442;
    wire N__45439;
    wire N__45436;
    wire N__45429;
    wire N__45420;
    wire N__45415;
    wire N__45410;
    wire N__45405;
    wire N__45400;
    wire N__45397;
    wire N__45394;
    wire N__45391;
    wire N__45384;
    wire N__45383;
    wire N__45382;
    wire N__45381;
    wire N__45380;
    wire N__45379;
    wire N__45378;
    wire N__45377;
    wire N__45376;
    wire N__45375;
    wire N__45374;
    wire N__45373;
    wire N__45370;
    wire N__45367;
    wire N__45366;
    wire N__45365;
    wire N__45362;
    wire N__45359;
    wire N__45356;
    wire N__45353;
    wire N__45352;
    wire N__45351;
    wire N__45350;
    wire N__45349;
    wire N__45344;
    wire N__45339;
    wire N__45334;
    wire N__45331;
    wire N__45328;
    wire N__45323;
    wire N__45320;
    wire N__45313;
    wire N__45304;
    wire N__45299;
    wire N__45296;
    wire N__45293;
    wire N__45290;
    wire N__45281;
    wire N__45278;
    wire N__45275;
    wire N__45272;
    wire N__45267;
    wire N__45258;
    wire N__45255;
    wire N__45254;
    wire N__45253;
    wire N__45250;
    wire N__45245;
    wire N__45240;
    wire N__45237;
    wire N__45236;
    wire N__45233;
    wire N__45230;
    wire N__45225;
    wire N__45222;
    wire N__45219;
    wire N__45216;
    wire N__45215;
    wire N__45214;
    wire N__45213;
    wire N__45212;
    wire N__45211;
    wire N__45208;
    wire N__45205;
    wire N__45202;
    wire N__45199;
    wire N__45196;
    wire N__45193;
    wire N__45180;
    wire N__45177;
    wire N__45176;
    wire N__45173;
    wire N__45170;
    wire N__45169;
    wire N__45168;
    wire N__45167;
    wire N__45166;
    wire N__45161;
    wire N__45158;
    wire N__45155;
    wire N__45152;
    wire N__45149;
    wire N__45144;
    wire N__45141;
    wire N__45138;
    wire N__45133;
    wire N__45126;
    wire N__45123;
    wire N__45120;
    wire N__45117;
    wire N__45114;
    wire N__45111;
    wire N__45110;
    wire N__45107;
    wire N__45104;
    wire N__45101;
    wire N__45098;
    wire N__45095;
    wire N__45092;
    wire N__45087;
    wire N__45084;
    wire N__45081;
    wire N__45078;
    wire N__45075;
    wire N__45072;
    wire N__45069;
    wire N__45066;
    wire N__45063;
    wire N__45060;
    wire N__45057;
    wire N__45054;
    wire N__45051;
    wire N__45050;
    wire N__45047;
    wire N__45044;
    wire N__45039;
    wire N__45036;
    wire N__45033;
    wire N__45030;
    wire N__45027;
    wire N__45024;
    wire N__45021;
    wire N__45018;
    wire N__45015;
    wire N__45012;
    wire N__45009;
    wire N__45006;
    wire N__45003;
    wire N__45000;
    wire N__44997;
    wire N__44994;
    wire N__44991;
    wire N__44988;
    wire N__44985;
    wire N__44982;
    wire N__44979;
    wire N__44976;
    wire N__44973;
    wire N__44972;
    wire N__44967;
    wire N__44966;
    wire N__44965;
    wire N__44964;
    wire N__44963;
    wire N__44960;
    wire N__44955;
    wire N__44954;
    wire N__44953;
    wire N__44950;
    wire N__44947;
    wire N__44944;
    wire N__44941;
    wire N__44934;
    wire N__44925;
    wire N__44922;
    wire N__44919;
    wire N__44916;
    wire N__44915;
    wire N__44912;
    wire N__44909;
    wire N__44904;
    wire N__44901;
    wire N__44898;
    wire N__44895;
    wire N__44892;
    wire N__44889;
    wire N__44886;
    wire N__44883;
    wire N__44882;
    wire N__44879;
    wire N__44876;
    wire N__44871;
    wire N__44868;
    wire N__44865;
    wire N__44862;
    wire N__44859;
    wire N__44856;
    wire N__44853;
    wire N__44850;
    wire N__44849;
    wire N__44846;
    wire N__44843;
    wire N__44840;
    wire N__44837;
    wire N__44834;
    wire N__44831;
    wire N__44826;
    wire N__44823;
    wire N__44820;
    wire N__44817;
    wire N__44814;
    wire N__44813;
    wire N__44810;
    wire N__44807;
    wire N__44804;
    wire N__44801;
    wire N__44798;
    wire N__44795;
    wire N__44790;
    wire N__44787;
    wire N__44784;
    wire N__44781;
    wire N__44778;
    wire N__44775;
    wire N__44774;
    wire N__44773;
    wire N__44770;
    wire N__44765;
    wire N__44762;
    wire N__44759;
    wire N__44754;
    wire N__44751;
    wire N__44750;
    wire N__44747;
    wire N__44744;
    wire N__44741;
    wire N__44740;
    wire N__44739;
    wire N__44734;
    wire N__44731;
    wire N__44728;
    wire N__44725;
    wire N__44722;
    wire N__44715;
    wire N__44712;
    wire N__44711;
    wire N__44710;
    wire N__44709;
    wire N__44708;
    wire N__44703;
    wire N__44700;
    wire N__44699;
    wire N__44694;
    wire N__44691;
    wire N__44688;
    wire N__44685;
    wire N__44676;
    wire N__44673;
    wire N__44670;
    wire N__44667;
    wire N__44664;
    wire N__44661;
    wire N__44658;
    wire N__44657;
    wire N__44656;
    wire N__44653;
    wire N__44650;
    wire N__44647;
    wire N__44644;
    wire N__44641;
    wire N__44638;
    wire N__44635;
    wire N__44632;
    wire N__44625;
    wire N__44622;
    wire N__44621;
    wire N__44618;
    wire N__44615;
    wire N__44612;
    wire N__44609;
    wire N__44606;
    wire N__44603;
    wire N__44598;
    wire N__44595;
    wire N__44592;
    wire N__44589;
    wire N__44586;
    wire N__44583;
    wire N__44580;
    wire N__44577;
    wire N__44574;
    wire N__44571;
    wire N__44570;
    wire N__44567;
    wire N__44564;
    wire N__44559;
    wire N__44556;
    wire N__44553;
    wire N__44552;
    wire N__44551;
    wire N__44548;
    wire N__44545;
    wire N__44542;
    wire N__44539;
    wire N__44536;
    wire N__44533;
    wire N__44530;
    wire N__44527;
    wire N__44520;
    wire N__44517;
    wire N__44514;
    wire N__44511;
    wire N__44510;
    wire N__44507;
    wire N__44504;
    wire N__44499;
    wire N__44496;
    wire N__44493;
    wire N__44490;
    wire N__44489;
    wire N__44486;
    wire N__44483;
    wire N__44480;
    wire N__44477;
    wire N__44474;
    wire N__44471;
    wire N__44466;
    wire N__44463;
    wire N__44460;
    wire N__44459;
    wire N__44456;
    wire N__44453;
    wire N__44450;
    wire N__44447;
    wire N__44442;
    wire N__44439;
    wire N__44436;
    wire N__44433;
    wire N__44432;
    wire N__44429;
    wire N__44426;
    wire N__44423;
    wire N__44420;
    wire N__44415;
    wire N__44414;
    wire N__44411;
    wire N__44408;
    wire N__44405;
    wire N__44400;
    wire N__44397;
    wire N__44394;
    wire N__44391;
    wire N__44388;
    wire N__44385;
    wire N__44382;
    wire N__44381;
    wire N__44378;
    wire N__44375;
    wire N__44370;
    wire N__44367;
    wire N__44364;
    wire N__44361;
    wire N__44358;
    wire N__44355;
    wire N__44352;
    wire N__44349;
    wire N__44346;
    wire N__44343;
    wire N__44340;
    wire N__44337;
    wire N__44334;
    wire N__44331;
    wire N__44328;
    wire N__44325;
    wire N__44322;
    wire N__44319;
    wire N__44316;
    wire N__44313;
    wire N__44310;
    wire N__44309;
    wire N__44306;
    wire N__44303;
    wire N__44298;
    wire N__44295;
    wire N__44292;
    wire N__44289;
    wire N__44286;
    wire N__44283;
    wire N__44280;
    wire N__44277;
    wire N__44274;
    wire N__44271;
    wire N__44268;
    wire N__44265;
    wire N__44262;
    wire N__44259;
    wire N__44258;
    wire N__44255;
    wire N__44252;
    wire N__44247;
    wire N__44244;
    wire N__44241;
    wire N__44238;
    wire N__44235;
    wire N__44232;
    wire N__44229;
    wire N__44226;
    wire N__44223;
    wire N__44220;
    wire N__44217;
    wire N__44214;
    wire N__44211;
    wire N__44208;
    wire N__44205;
    wire N__44204;
    wire N__44201;
    wire N__44198;
    wire N__44195;
    wire N__44192;
    wire N__44187;
    wire N__44184;
    wire N__44181;
    wire N__44178;
    wire N__44175;
    wire N__44172;
    wire N__44169;
    wire N__44166;
    wire N__44163;
    wire N__44160;
    wire N__44157;
    wire N__44156;
    wire N__44153;
    wire N__44150;
    wire N__44145;
    wire N__44142;
    wire N__44139;
    wire N__44136;
    wire N__44133;
    wire N__44130;
    wire N__44127;
    wire N__44126;
    wire N__44123;
    wire N__44120;
    wire N__44115;
    wire N__44112;
    wire N__44109;
    wire N__44106;
    wire N__44105;
    wire N__44100;
    wire N__44097;
    wire N__44094;
    wire N__44091;
    wire N__44088;
    wire N__44085;
    wire N__44082;
    wire N__44081;
    wire N__44076;
    wire N__44073;
    wire N__44070;
    wire N__44069;
    wire N__44068;
    wire N__44065;
    wire N__44060;
    wire N__44055;
    wire N__44052;
    wire N__44049;
    wire N__44048;
    wire N__44045;
    wire N__44042;
    wire N__44037;
    wire N__44034;
    wire N__44031;
    wire N__44028;
    wire N__44025;
    wire N__44022;
    wire N__44019;
    wire N__44016;
    wire N__44013;
    wire N__44010;
    wire N__44007;
    wire N__44006;
    wire N__44001;
    wire N__43998;
    wire N__43997;
    wire N__43992;
    wire N__43989;
    wire N__43986;
    wire N__43983;
    wire N__43980;
    wire N__43977;
    wire N__43974;
    wire N__43971;
    wire N__43968;
    wire N__43965;
    wire N__43962;
    wire N__43959;
    wire N__43958;
    wire N__43955;
    wire N__43952;
    wire N__43947;
    wire N__43944;
    wire N__43943;
    wire N__43940;
    wire N__43937;
    wire N__43932;
    wire N__43931;
    wire N__43930;
    wire N__43927;
    wire N__43922;
    wire N__43917;
    wire N__43914;
    wire N__43911;
    wire N__43910;
    wire N__43905;
    wire N__43902;
    wire N__43899;
    wire N__43898;
    wire N__43893;
    wire N__43890;
    wire N__43889;
    wire N__43884;
    wire N__43881;
    wire N__43878;
    wire N__43875;
    wire N__43872;
    wire N__43869;
    wire N__43866;
    wire N__43865;
    wire N__43860;
    wire N__43857;
    wire N__43854;
    wire N__43851;
    wire N__43848;
    wire N__43845;
    wire N__43842;
    wire N__43839;
    wire N__43836;
    wire N__43833;
    wire N__43830;
    wire N__43829;
    wire N__43824;
    wire N__43821;
    wire N__43818;
    wire N__43815;
    wire N__43812;
    wire N__43809;
    wire N__43806;
    wire N__43803;
    wire N__43800;
    wire N__43797;
    wire N__43794;
    wire N__43791;
    wire N__43788;
    wire N__43785;
    wire N__43782;
    wire N__43779;
    wire N__43776;
    wire N__43773;
    wire N__43770;
    wire N__43767;
    wire N__43764;
    wire N__43763;
    wire N__43760;
    wire N__43757;
    wire N__43752;
    wire N__43749;
    wire N__43746;
    wire N__43745;
    wire N__43742;
    wire N__43739;
    wire N__43734;
    wire N__43731;
    wire N__43730;
    wire N__43727;
    wire N__43724;
    wire N__43719;
    wire N__43716;
    wire N__43713;
    wire N__43710;
    wire N__43707;
    wire N__43704;
    wire N__43701;
    wire N__43698;
    wire N__43695;
    wire N__43692;
    wire N__43689;
    wire N__43686;
    wire N__43683;
    wire N__43680;
    wire N__43677;
    wire N__43674;
    wire N__43671;
    wire N__43668;
    wire N__43665;
    wire N__43662;
    wire N__43659;
    wire N__43656;
    wire N__43653;
    wire N__43650;
    wire N__43647;
    wire N__43644;
    wire N__43641;
    wire N__43638;
    wire N__43635;
    wire N__43632;
    wire N__43629;
    wire N__43626;
    wire N__43623;
    wire N__43620;
    wire N__43617;
    wire N__43614;
    wire N__43611;
    wire N__43608;
    wire N__43605;
    wire N__43602;
    wire N__43599;
    wire N__43596;
    wire N__43593;
    wire N__43590;
    wire N__43587;
    wire N__43584;
    wire N__43581;
    wire N__43578;
    wire N__43575;
    wire N__43572;
    wire N__43569;
    wire N__43566;
    wire N__43563;
    wire N__43560;
    wire N__43557;
    wire N__43554;
    wire N__43551;
    wire N__43548;
    wire N__43545;
    wire N__43542;
    wire N__43539;
    wire N__43536;
    wire N__43533;
    wire N__43530;
    wire N__43527;
    wire N__43524;
    wire N__43521;
    wire N__43518;
    wire N__43515;
    wire N__43512;
    wire N__43509;
    wire N__43506;
    wire N__43503;
    wire N__43500;
    wire N__43497;
    wire N__43494;
    wire N__43491;
    wire N__43488;
    wire N__43485;
    wire N__43482;
    wire N__43479;
    wire N__43476;
    wire N__43473;
    wire N__43470;
    wire N__43467;
    wire N__43464;
    wire N__43461;
    wire N__43458;
    wire N__43455;
    wire N__43452;
    wire N__43449;
    wire N__43446;
    wire N__43443;
    wire N__43440;
    wire N__43437;
    wire N__43434;
    wire N__43431;
    wire N__43428;
    wire N__43425;
    wire N__43424;
    wire N__43421;
    wire N__43418;
    wire N__43415;
    wire N__43414;
    wire N__43411;
    wire N__43408;
    wire N__43405;
    wire N__43398;
    wire N__43395;
    wire N__43392;
    wire N__43389;
    wire N__43386;
    wire N__43383;
    wire N__43380;
    wire N__43377;
    wire N__43374;
    wire N__43371;
    wire N__43370;
    wire N__43367;
    wire N__43364;
    wire N__43359;
    wire N__43356;
    wire N__43353;
    wire N__43350;
    wire N__43347;
    wire N__43344;
    wire N__43341;
    wire N__43338;
    wire N__43337;
    wire N__43336;
    wire N__43333;
    wire N__43330;
    wire N__43327;
    wire N__43320;
    wire N__43317;
    wire N__43314;
    wire N__43313;
    wire N__43312;
    wire N__43309;
    wire N__43304;
    wire N__43299;
    wire N__43296;
    wire N__43295;
    wire N__43294;
    wire N__43287;
    wire N__43284;
    wire N__43281;
    wire N__43280;
    wire N__43277;
    wire N__43276;
    wire N__43273;
    wire N__43270;
    wire N__43265;
    wire N__43260;
    wire N__43257;
    wire N__43256;
    wire N__43253;
    wire N__43250;
    wire N__43247;
    wire N__43244;
    wire N__43243;
    wire N__43242;
    wire N__43237;
    wire N__43232;
    wire N__43227;
    wire N__43224;
    wire N__43223;
    wire N__43220;
    wire N__43217;
    wire N__43216;
    wire N__43213;
    wire N__43212;
    wire N__43209;
    wire N__43206;
    wire N__43203;
    wire N__43200;
    wire N__43191;
    wire N__43188;
    wire N__43187;
    wire N__43186;
    wire N__43183;
    wire N__43180;
    wire N__43177;
    wire N__43174;
    wire N__43171;
    wire N__43166;
    wire N__43161;
    wire N__43158;
    wire N__43157;
    wire N__43156;
    wire N__43153;
    wire N__43148;
    wire N__43145;
    wire N__43142;
    wire N__43137;
    wire N__43134;
    wire N__43131;
    wire N__43128;
    wire N__43127;
    wire N__43124;
    wire N__43121;
    wire N__43116;
    wire N__43113;
    wire N__43110;
    wire N__43107;
    wire N__43104;
    wire N__43101;
    wire N__43098;
    wire N__43097;
    wire N__43096;
    wire N__43095;
    wire N__43094;
    wire N__43093;
    wire N__43084;
    wire N__43079;
    wire N__43076;
    wire N__43073;
    wire N__43070;
    wire N__43065;
    wire N__43064;
    wire N__43063;
    wire N__43060;
    wire N__43057;
    wire N__43052;
    wire N__43047;
    wire N__43046;
    wire N__43045;
    wire N__43042;
    wire N__43039;
    wire N__43036;
    wire N__43029;
    wire N__43026;
    wire N__43023;
    wire N__43020;
    wire N__43017;
    wire N__43016;
    wire N__43013;
    wire N__43010;
    wire N__43005;
    wire N__43002;
    wire N__42999;
    wire N__42996;
    wire N__42993;
    wire N__42990;
    wire N__42987;
    wire N__42984;
    wire N__42981;
    wire N__42980;
    wire N__42975;
    wire N__42972;
    wire N__42969;
    wire N__42966;
    wire N__42965;
    wire N__42962;
    wire N__42959;
    wire N__42956;
    wire N__42953;
    wire N__42948;
    wire N__42945;
    wire N__42942;
    wire N__42939;
    wire N__42936;
    wire N__42933;
    wire N__42930;
    wire N__42929;
    wire N__42926;
    wire N__42923;
    wire N__42920;
    wire N__42915;
    wire N__42914;
    wire N__42911;
    wire N__42908;
    wire N__42903;
    wire N__42902;
    wire N__42899;
    wire N__42896;
    wire N__42893;
    wire N__42888;
    wire N__42887;
    wire N__42884;
    wire N__42881;
    wire N__42876;
    wire N__42873;
    wire N__42872;
    wire N__42869;
    wire N__42866;
    wire N__42863;
    wire N__42858;
    wire N__42857;
    wire N__42854;
    wire N__42851;
    wire N__42846;
    wire N__42845;
    wire N__42842;
    wire N__42839;
    wire N__42834;
    wire N__42833;
    wire N__42830;
    wire N__42827;
    wire N__42824;
    wire N__42819;
    wire N__42816;
    wire N__42813;
    wire N__42810;
    wire N__42807;
    wire N__42806;
    wire N__42805;
    wire N__42802;
    wire N__42797;
    wire N__42792;
    wire N__42791;
    wire N__42790;
    wire N__42789;
    wire N__42786;
    wire N__42783;
    wire N__42778;
    wire N__42771;
    wire N__42768;
    wire N__42767;
    wire N__42766;
    wire N__42763;
    wire N__42758;
    wire N__42753;
    wire N__42750;
    wire N__42749;
    wire N__42748;
    wire N__42747;
    wire N__42744;
    wire N__42741;
    wire N__42738;
    wire N__42735;
    wire N__42726;
    wire N__42723;
    wire N__42722;
    wire N__42721;
    wire N__42718;
    wire N__42715;
    wire N__42714;
    wire N__42711;
    wire N__42708;
    wire N__42705;
    wire N__42702;
    wire N__42699;
    wire N__42690;
    wire N__42687;
    wire N__42684;
    wire N__42681;
    wire N__42678;
    wire N__42675;
    wire N__42674;
    wire N__42673;
    wire N__42670;
    wire N__42667;
    wire N__42664;
    wire N__42663;
    wire N__42658;
    wire N__42653;
    wire N__42650;
    wire N__42647;
    wire N__42642;
    wire N__42639;
    wire N__42636;
    wire N__42633;
    wire N__42630;
    wire N__42627;
    wire N__42624;
    wire N__42621;
    wire N__42620;
    wire N__42615;
    wire N__42612;
    wire N__42609;
    wire N__42606;
    wire N__42603;
    wire N__42600;
    wire N__42597;
    wire N__42594;
    wire N__42591;
    wire N__42588;
    wire N__42587;
    wire N__42582;
    wire N__42579;
    wire N__42576;
    wire N__42573;
    wire N__42570;
    wire N__42567;
    wire N__42564;
    wire N__42561;
    wire N__42558;
    wire N__42555;
    wire N__42554;
    wire N__42549;
    wire N__42546;
    wire N__42543;
    wire N__42540;
    wire N__42537;
    wire N__42534;
    wire N__42531;
    wire N__42528;
    wire N__42525;
    wire N__42522;
    wire N__42521;
    wire N__42516;
    wire N__42513;
    wire N__42510;
    wire N__42507;
    wire N__42504;
    wire N__42501;
    wire N__42498;
    wire N__42495;
    wire N__42492;
    wire N__42489;
    wire N__42488;
    wire N__42483;
    wire N__42480;
    wire N__42477;
    wire N__42474;
    wire N__42471;
    wire N__42468;
    wire N__42465;
    wire N__42462;
    wire N__42459;
    wire N__42456;
    wire N__42453;
    wire N__42450;
    wire N__42447;
    wire N__42444;
    wire N__42441;
    wire N__42438;
    wire N__42435;
    wire N__42432;
    wire N__42429;
    wire N__42426;
    wire N__42425;
    wire N__42422;
    wire N__42421;
    wire N__42418;
    wire N__42415;
    wire N__42412;
    wire N__42409;
    wire N__42406;
    wire N__42403;
    wire N__42396;
    wire N__42393;
    wire N__42390;
    wire N__42387;
    wire N__42384;
    wire N__42381;
    wire N__42378;
    wire N__42375;
    wire N__42372;
    wire N__42369;
    wire N__42366;
    wire N__42363;
    wire N__42360;
    wire N__42357;
    wire N__42356;
    wire N__42353;
    wire N__42350;
    wire N__42347;
    wire N__42344;
    wire N__42339;
    wire N__42336;
    wire N__42333;
    wire N__42330;
    wire N__42327;
    wire N__42324;
    wire N__42321;
    wire N__42318;
    wire N__42315;
    wire N__42314;
    wire N__42311;
    wire N__42308;
    wire N__42305;
    wire N__42302;
    wire N__42299;
    wire N__42296;
    wire N__42293;
    wire N__42288;
    wire N__42287;
    wire N__42286;
    wire N__42283;
    wire N__42276;
    wire N__42273;
    wire N__42270;
    wire N__42267;
    wire N__42264;
    wire N__42261;
    wire N__42258;
    wire N__42255;
    wire N__42252;
    wire N__42249;
    wire N__42246;
    wire N__42243;
    wire N__42240;
    wire N__42237;
    wire N__42234;
    wire N__42233;
    wire N__42228;
    wire N__42225;
    wire N__42222;
    wire N__42219;
    wire N__42218;
    wire N__42217;
    wire N__42210;
    wire N__42207;
    wire N__42206;
    wire N__42203;
    wire N__42202;
    wire N__42199;
    wire N__42192;
    wire N__42189;
    wire N__42188;
    wire N__42187;
    wire N__42186;
    wire N__42185;
    wire N__42174;
    wire N__42171;
    wire N__42168;
    wire N__42167;
    wire N__42166;
    wire N__42163;
    wire N__42158;
    wire N__42153;
    wire N__42150;
    wire N__42147;
    wire N__42146;
    wire N__42145;
    wire N__42142;
    wire N__42137;
    wire N__42134;
    wire N__42129;
    wire N__42126;
    wire N__42125;
    wire N__42122;
    wire N__42119;
    wire N__42114;
    wire N__42113;
    wire N__42112;
    wire N__42105;
    wire N__42102;
    wire N__42099;
    wire N__42096;
    wire N__42095;
    wire N__42092;
    wire N__42089;
    wire N__42084;
    wire N__42081;
    wire N__42078;
    wire N__42075;
    wire N__42072;
    wire N__42069;
    wire N__42068;
    wire N__42063;
    wire N__42060;
    wire N__42057;
    wire N__42056;
    wire N__42053;
    wire N__42050;
    wire N__42045;
    wire N__42042;
    wire N__42039;
    wire N__42036;
    wire N__42033;
    wire N__42030;
    wire N__42027;
    wire N__42024;
    wire N__42021;
    wire N__42018;
    wire N__42017;
    wire N__42016;
    wire N__42013;
    wire N__42008;
    wire N__42003;
    wire N__42000;
    wire N__41997;
    wire N__41994;
    wire N__41993;
    wire N__41990;
    wire N__41987;
    wire N__41984;
    wire N__41979;
    wire N__41976;
    wire N__41973;
    wire N__41970;
    wire N__41967;
    wire N__41964;
    wire N__41961;
    wire N__41960;
    wire N__41957;
    wire N__41956;
    wire N__41955;
    wire N__41952;
    wire N__41951;
    wire N__41944;
    wire N__41941;
    wire N__41938;
    wire N__41935;
    wire N__41930;
    wire N__41927;
    wire N__41924;
    wire N__41919;
    wire N__41916;
    wire N__41915;
    wire N__41914;
    wire N__41913;
    wire N__41910;
    wire N__41907;
    wire N__41906;
    wire N__41903;
    wire N__41900;
    wire N__41897;
    wire N__41894;
    wire N__41887;
    wire N__41880;
    wire N__41877;
    wire N__41874;
    wire N__41873;
    wire N__41872;
    wire N__41869;
    wire N__41868;
    wire N__41865;
    wire N__41862;
    wire N__41859;
    wire N__41854;
    wire N__41847;
    wire N__41846;
    wire N__41843;
    wire N__41840;
    wire N__41835;
    wire N__41832;
    wire N__41829;
    wire N__41826;
    wire N__41823;
    wire N__41820;
    wire N__41817;
    wire N__41814;
    wire N__41811;
    wire N__41810;
    wire N__41807;
    wire N__41804;
    wire N__41801;
    wire N__41798;
    wire N__41795;
    wire N__41790;
    wire N__41787;
    wire N__41784;
    wire N__41781;
    wire N__41778;
    wire N__41775;
    wire N__41772;
    wire N__41769;
    wire N__41766;
    wire N__41763;
    wire N__41760;
    wire N__41757;
    wire N__41754;
    wire N__41751;
    wire N__41748;
    wire N__41745;
    wire N__41742;
    wire N__41739;
    wire N__41736;
    wire N__41733;
    wire N__41730;
    wire N__41727;
    wire N__41724;
    wire N__41721;
    wire N__41718;
    wire N__41715;
    wire N__41714;
    wire N__41711;
    wire N__41708;
    wire N__41707;
    wire N__41704;
    wire N__41701;
    wire N__41700;
    wire N__41697;
    wire N__41694;
    wire N__41691;
    wire N__41688;
    wire N__41679;
    wire N__41678;
    wire N__41677;
    wire N__41674;
    wire N__41671;
    wire N__41668;
    wire N__41665;
    wire N__41662;
    wire N__41659;
    wire N__41652;
    wire N__41651;
    wire N__41650;
    wire N__41649;
    wire N__41646;
    wire N__41645;
    wire N__41642;
    wire N__41639;
    wire N__41636;
    wire N__41633;
    wire N__41630;
    wire N__41629;
    wire N__41628;
    wire N__41627;
    wire N__41624;
    wire N__41619;
    wire N__41616;
    wire N__41611;
    wire N__41606;
    wire N__41601;
    wire N__41596;
    wire N__41589;
    wire N__41588;
    wire N__41587;
    wire N__41586;
    wire N__41585;
    wire N__41584;
    wire N__41583;
    wire N__41568;
    wire N__41567;
    wire N__41566;
    wire N__41565;
    wire N__41562;
    wire N__41559;
    wire N__41556;
    wire N__41555;
    wire N__41552;
    wire N__41549;
    wire N__41544;
    wire N__41541;
    wire N__41532;
    wire N__41531;
    wire N__41528;
    wire N__41525;
    wire N__41522;
    wire N__41519;
    wire N__41516;
    wire N__41513;
    wire N__41510;
    wire N__41507;
    wire N__41502;
    wire N__41501;
    wire N__41500;
    wire N__41497;
    wire N__41494;
    wire N__41491;
    wire N__41488;
    wire N__41485;
    wire N__41482;
    wire N__41479;
    wire N__41476;
    wire N__41469;
    wire N__41466;
    wire N__41463;
    wire N__41460;
    wire N__41457;
    wire N__41454;
    wire N__41451;
    wire N__41448;
    wire N__41445;
    wire N__41442;
    wire N__41439;
    wire N__41436;
    wire N__41435;
    wire N__41432;
    wire N__41431;
    wire N__41428;
    wire N__41425;
    wire N__41422;
    wire N__41419;
    wire N__41416;
    wire N__41409;
    wire N__41408;
    wire N__41407;
    wire N__41404;
    wire N__41401;
    wire N__41398;
    wire N__41395;
    wire N__41392;
    wire N__41389;
    wire N__41386;
    wire N__41379;
    wire N__41376;
    wire N__41373;
    wire N__41370;
    wire N__41367;
    wire N__41364;
    wire N__41363;
    wire N__41362;
    wire N__41359;
    wire N__41354;
    wire N__41351;
    wire N__41348;
    wire N__41345;
    wire N__41344;
    wire N__41341;
    wire N__41338;
    wire N__41335;
    wire N__41332;
    wire N__41325;
    wire N__41322;
    wire N__41321;
    wire N__41318;
    wire N__41315;
    wire N__41310;
    wire N__41307;
    wire N__41304;
    wire N__41301;
    wire N__41298;
    wire N__41295;
    wire N__41292;
    wire N__41291;
    wire N__41288;
    wire N__41285;
    wire N__41282;
    wire N__41279;
    wire N__41276;
    wire N__41273;
    wire N__41270;
    wire N__41267;
    wire N__41264;
    wire N__41261;
    wire N__41256;
    wire N__41253;
    wire N__41250;
    wire N__41247;
    wire N__41244;
    wire N__41241;
    wire N__41238;
    wire N__41235;
    wire N__41232;
    wire N__41231;
    wire N__41228;
    wire N__41225;
    wire N__41224;
    wire N__41219;
    wire N__41216;
    wire N__41213;
    wire N__41208;
    wire N__41205;
    wire N__41202;
    wire N__41199;
    wire N__41196;
    wire N__41193;
    wire N__41190;
    wire N__41187;
    wire N__41184;
    wire N__41183;
    wire N__41180;
    wire N__41177;
    wire N__41174;
    wire N__41169;
    wire N__41166;
    wire N__41163;
    wire N__41162;
    wire N__41159;
    wire N__41156;
    wire N__41151;
    wire N__41150;
    wire N__41147;
    wire N__41144;
    wire N__41139;
    wire N__41136;
    wire N__41133;
    wire N__41132;
    wire N__41129;
    wire N__41126;
    wire N__41121;
    wire N__41118;
    wire N__41117;
    wire N__41114;
    wire N__41111;
    wire N__41106;
    wire N__41105;
    wire N__41102;
    wire N__41099;
    wire N__41096;
    wire N__41091;
    wire N__41088;
    wire N__41087;
    wire N__41084;
    wire N__41081;
    wire N__41076;
    wire N__41073;
    wire N__41070;
    wire N__41067;
    wire N__41064;
    wire N__41061;
    wire N__41058;
    wire N__41055;
    wire N__41052;
    wire N__41051;
    wire N__41050;
    wire N__41049;
    wire N__41046;
    wire N__41041;
    wire N__41038;
    wire N__41031;
    wire N__41030;
    wire N__41027;
    wire N__41026;
    wire N__41023;
    wire N__41018;
    wire N__41017;
    wire N__41012;
    wire N__41009;
    wire N__41006;
    wire N__41001;
    wire N__40998;
    wire N__40997;
    wire N__40996;
    wire N__40993;
    wire N__40988;
    wire N__40983;
    wire N__40980;
    wire N__40977;
    wire N__40974;
    wire N__40973;
    wire N__40972;
    wire N__40971;
    wire N__40968;
    wire N__40965;
    wire N__40962;
    wire N__40959;
    wire N__40950;
    wire N__40949;
    wire N__40946;
    wire N__40945;
    wire N__40942;
    wire N__40939;
    wire N__40936;
    wire N__40933;
    wire N__40930;
    wire N__40923;
    wire N__40920;
    wire N__40917;
    wire N__40914;
    wire N__40913;
    wire N__40910;
    wire N__40907;
    wire N__40902;
    wire N__40899;
    wire N__40896;
    wire N__40895;
    wire N__40892;
    wire N__40889;
    wire N__40884;
    wire N__40881;
    wire N__40878;
    wire N__40875;
    wire N__40874;
    wire N__40871;
    wire N__40868;
    wire N__40863;
    wire N__40860;
    wire N__40859;
    wire N__40856;
    wire N__40853;
    wire N__40850;
    wire N__40845;
    wire N__40842;
    wire N__40841;
    wire N__40838;
    wire N__40835;
    wire N__40832;
    wire N__40827;
    wire N__40824;
    wire N__40821;
    wire N__40820;
    wire N__40817;
    wire N__40814;
    wire N__40809;
    wire N__40806;
    wire N__40803;
    wire N__40800;
    wire N__40799;
    wire N__40796;
    wire N__40793;
    wire N__40788;
    wire N__40785;
    wire N__40784;
    wire N__40781;
    wire N__40778;
    wire N__40773;
    wire N__40770;
    wire N__40769;
    wire N__40766;
    wire N__40763;
    wire N__40758;
    wire N__40755;
    wire N__40754;
    wire N__40751;
    wire N__40748;
    wire N__40743;
    wire N__40740;
    wire N__40739;
    wire N__40736;
    wire N__40733;
    wire N__40728;
    wire N__40725;
    wire N__40724;
    wire N__40721;
    wire N__40718;
    wire N__40713;
    wire N__40710;
    wire N__40709;
    wire N__40706;
    wire N__40703;
    wire N__40700;
    wire N__40695;
    wire N__40692;
    wire N__40689;
    wire N__40686;
    wire N__40683;
    wire N__40680;
    wire N__40677;
    wire N__40674;
    wire N__40671;
    wire N__40668;
    wire N__40665;
    wire N__40662;
    wire N__40659;
    wire N__40656;
    wire N__40653;
    wire N__40650;
    wire N__40647;
    wire N__40644;
    wire N__40641;
    wire N__40638;
    wire N__40635;
    wire N__40632;
    wire N__40629;
    wire N__40626;
    wire N__40623;
    wire N__40620;
    wire N__40617;
    wire N__40614;
    wire N__40611;
    wire N__40608;
    wire N__40605;
    wire N__40602;
    wire N__40599;
    wire N__40596;
    wire N__40593;
    wire N__40590;
    wire N__40587;
    wire N__40584;
    wire N__40581;
    wire N__40578;
    wire N__40577;
    wire N__40574;
    wire N__40571;
    wire N__40566;
    wire N__40563;
    wire N__40560;
    wire N__40559;
    wire N__40556;
    wire N__40553;
    wire N__40552;
    wire N__40551;
    wire N__40546;
    wire N__40543;
    wire N__40540;
    wire N__40535;
    wire N__40532;
    wire N__40531;
    wire N__40528;
    wire N__40525;
    wire N__40522;
    wire N__40521;
    wire N__40514;
    wire N__40511;
    wire N__40506;
    wire N__40503;
    wire N__40500;
    wire N__40497;
    wire N__40494;
    wire N__40493;
    wire N__40492;
    wire N__40491;
    wire N__40490;
    wire N__40489;
    wire N__40488;
    wire N__40487;
    wire N__40482;
    wire N__40469;
    wire N__40466;
    wire N__40463;
    wire N__40460;
    wire N__40455;
    wire N__40452;
    wire N__40449;
    wire N__40446;
    wire N__40443;
    wire N__40442;
    wire N__40441;
    wire N__40440;
    wire N__40439;
    wire N__40436;
    wire N__40429;
    wire N__40428;
    wire N__40427;
    wire N__40424;
    wire N__40423;
    wire N__40420;
    wire N__40417;
    wire N__40410;
    wire N__40407;
    wire N__40402;
    wire N__40399;
    wire N__40392;
    wire N__40389;
    wire N__40386;
    wire N__40385;
    wire N__40384;
    wire N__40383;
    wire N__40382;
    wire N__40379;
    wire N__40372;
    wire N__40371;
    wire N__40370;
    wire N__40369;
    wire N__40366;
    wire N__40365;
    wire N__40362;
    wire N__40359;
    wire N__40352;
    wire N__40349;
    wire N__40346;
    wire N__40341;
    wire N__40338;
    wire N__40329;
    wire N__40326;
    wire N__40323;
    wire N__40322;
    wire N__40319;
    wire N__40316;
    wire N__40313;
    wire N__40312;
    wire N__40309;
    wire N__40306;
    wire N__40303;
    wire N__40298;
    wire N__40293;
    wire N__40290;
    wire N__40287;
    wire N__40284;
    wire N__40283;
    wire N__40280;
    wire N__40277;
    wire N__40274;
    wire N__40271;
    wire N__40266;
    wire N__40263;
    wire N__40260;
    wire N__40257;
    wire N__40254;
    wire N__40251;
    wire N__40250;
    wire N__40247;
    wire N__40244;
    wire N__40243;
    wire N__40242;
    wire N__40241;
    wire N__40240;
    wire N__40239;
    wire N__40238;
    wire N__40237;
    wire N__40234;
    wire N__40231;
    wire N__40228;
    wire N__40225;
    wire N__40222;
    wire N__40219;
    wire N__40216;
    wire N__40215;
    wire N__40214;
    wire N__40213;
    wire N__40212;
    wire N__40209;
    wire N__40206;
    wire N__40205;
    wire N__40202;
    wire N__40197;
    wire N__40180;
    wire N__40177;
    wire N__40174;
    wire N__40171;
    wire N__40168;
    wire N__40165;
    wire N__40156;
    wire N__40151;
    wire N__40148;
    wire N__40143;
    wire N__40142;
    wire N__40139;
    wire N__40138;
    wire N__40133;
    wire N__40130;
    wire N__40127;
    wire N__40122;
    wire N__40119;
    wire N__40118;
    wire N__40115;
    wire N__40114;
    wire N__40111;
    wire N__40108;
    wire N__40107;
    wire N__40104;
    wire N__40099;
    wire N__40096;
    wire N__40089;
    wire N__40086;
    wire N__40085;
    wire N__40082;
    wire N__40079;
    wire N__40076;
    wire N__40071;
    wire N__40070;
    wire N__40069;
    wire N__40066;
    wire N__40063;
    wire N__40058;
    wire N__40053;
    wire N__40050;
    wire N__40047;
    wire N__40044;
    wire N__40041;
    wire N__40038;
    wire N__40035;
    wire N__40032;
    wire N__40031;
    wire N__40028;
    wire N__40025;
    wire N__40020;
    wire N__40019;
    wire N__40014;
    wire N__40011;
    wire N__40008;
    wire N__40007;
    wire N__40006;
    wire N__40005;
    wire N__40002;
    wire N__40001;
    wire N__39998;
    wire N__39997;
    wire N__39994;
    wire N__39993;
    wire N__39992;
    wire N__39991;
    wire N__39976;
    wire N__39971;
    wire N__39968;
    wire N__39967;
    wire N__39962;
    wire N__39959;
    wire N__39954;
    wire N__39953;
    wire N__39952;
    wire N__39951;
    wire N__39950;
    wire N__39949;
    wire N__39948;
    wire N__39933;
    wire N__39932;
    wire N__39929;
    wire N__39928;
    wire N__39925;
    wire N__39922;
    wire N__39919;
    wire N__39912;
    wire N__39909;
    wire N__39906;
    wire N__39903;
    wire N__39900;
    wire N__39897;
    wire N__39896;
    wire N__39893;
    wire N__39890;
    wire N__39887;
    wire N__39884;
    wire N__39881;
    wire N__39876;
    wire N__39873;
    wire N__39872;
    wire N__39869;
    wire N__39868;
    wire N__39867;
    wire N__39860;
    wire N__39857;
    wire N__39854;
    wire N__39849;
    wire N__39846;
    wire N__39843;
    wire N__39840;
    wire N__39839;
    wire N__39836;
    wire N__39835;
    wire N__39830;
    wire N__39827;
    wire N__39824;
    wire N__39819;
    wire N__39816;
    wire N__39813;
    wire N__39812;
    wire N__39811;
    wire N__39810;
    wire N__39807;
    wire N__39802;
    wire N__39799;
    wire N__39798;
    wire N__39797;
    wire N__39792;
    wire N__39789;
    wire N__39784;
    wire N__39777;
    wire N__39776;
    wire N__39775;
    wire N__39774;
    wire N__39771;
    wire N__39768;
    wire N__39767;
    wire N__39764;
    wire N__39761;
    wire N__39756;
    wire N__39753;
    wire N__39748;
    wire N__39745;
    wire N__39742;
    wire N__39737;
    wire N__39734;
    wire N__39729;
    wire N__39726;
    wire N__39723;
    wire N__39720;
    wire N__39717;
    wire N__39714;
    wire N__39711;
    wire N__39708;
    wire N__39705;
    wire N__39702;
    wire N__39701;
    wire N__39696;
    wire N__39693;
    wire N__39692;
    wire N__39691;
    wire N__39688;
    wire N__39683;
    wire N__39678;
    wire N__39675;
    wire N__39672;
    wire N__39669;
    wire N__39666;
    wire N__39663;
    wire N__39660;
    wire N__39657;
    wire N__39654;
    wire N__39651;
    wire N__39648;
    wire N__39645;
    wire N__39642;
    wire N__39639;
    wire N__39636;
    wire N__39633;
    wire N__39630;
    wire N__39627;
    wire N__39624;
    wire N__39621;
    wire N__39620;
    wire N__39617;
    wire N__39614;
    wire N__39611;
    wire N__39606;
    wire N__39605;
    wire N__39604;
    wire N__39601;
    wire N__39598;
    wire N__39595;
    wire N__39592;
    wire N__39589;
    wire N__39586;
    wire N__39581;
    wire N__39576;
    wire N__39573;
    wire N__39572;
    wire N__39569;
    wire N__39566;
    wire N__39563;
    wire N__39558;
    wire N__39557;
    wire N__39556;
    wire N__39553;
    wire N__39550;
    wire N__39547;
    wire N__39544;
    wire N__39541;
    wire N__39538;
    wire N__39535;
    wire N__39532;
    wire N__39529;
    wire N__39522;
    wire N__39519;
    wire N__39518;
    wire N__39515;
    wire N__39512;
    wire N__39509;
    wire N__39504;
    wire N__39501;
    wire N__39500;
    wire N__39499;
    wire N__39496;
    wire N__39493;
    wire N__39490;
    wire N__39487;
    wire N__39480;
    wire N__39479;
    wire N__39476;
    wire N__39473;
    wire N__39470;
    wire N__39467;
    wire N__39464;
    wire N__39459;
    wire N__39458;
    wire N__39455;
    wire N__39452;
    wire N__39451;
    wire N__39450;
    wire N__39449;
    wire N__39448;
    wire N__39443;
    wire N__39434;
    wire N__39433;
    wire N__39432;
    wire N__39431;
    wire N__39426;
    wire N__39419;
    wire N__39414;
    wire N__39411;
    wire N__39410;
    wire N__39407;
    wire N__39404;
    wire N__39399;
    wire N__39398;
    wire N__39395;
    wire N__39392;
    wire N__39387;
    wire N__39386;
    wire N__39383;
    wire N__39380;
    wire N__39377;
    wire N__39372;
    wire N__39369;
    wire N__39368;
    wire N__39365;
    wire N__39362;
    wire N__39361;
    wire N__39358;
    wire N__39355;
    wire N__39352;
    wire N__39349;
    wire N__39342;
    wire N__39341;
    wire N__39338;
    wire N__39335;
    wire N__39330;
    wire N__39329;
    wire N__39326;
    wire N__39323;
    wire N__39320;
    wire N__39317;
    wire N__39314;
    wire N__39309;
    wire N__39308;
    wire N__39307;
    wire N__39304;
    wire N__39299;
    wire N__39298;
    wire N__39295;
    wire N__39292;
    wire N__39291;
    wire N__39290;
    wire N__39289;
    wire N__39288;
    wire N__39287;
    wire N__39286;
    wire N__39285;
    wire N__39284;
    wire N__39283;
    wire N__39280;
    wire N__39277;
    wire N__39274;
    wire N__39271;
    wire N__39264;
    wire N__39253;
    wire N__39240;
    wire N__39239;
    wire N__39236;
    wire N__39233;
    wire N__39230;
    wire N__39227;
    wire N__39224;
    wire N__39221;
    wire N__39220;
    wire N__39217;
    wire N__39214;
    wire N__39211;
    wire N__39208;
    wire N__39205;
    wire N__39198;
    wire N__39195;
    wire N__39192;
    wire N__39189;
    wire N__39186;
    wire N__39183;
    wire N__39180;
    wire N__39177;
    wire N__39174;
    wire N__39171;
    wire N__39168;
    wire N__39165;
    wire N__39162;
    wire N__39159;
    wire N__39156;
    wire N__39153;
    wire N__39150;
    wire N__39147;
    wire N__39144;
    wire N__39141;
    wire N__39138;
    wire N__39135;
    wire N__39132;
    wire N__39129;
    wire N__39126;
    wire N__39123;
    wire N__39120;
    wire N__39117;
    wire N__39114;
    wire N__39111;
    wire N__39108;
    wire N__39105;
    wire N__39102;
    wire N__39099;
    wire N__39096;
    wire N__39095;
    wire N__39094;
    wire N__39091;
    wire N__39088;
    wire N__39085;
    wire N__39078;
    wire N__39075;
    wire N__39074;
    wire N__39071;
    wire N__39068;
    wire N__39065;
    wire N__39060;
    wire N__39059;
    wire N__39056;
    wire N__39053;
    wire N__39052;
    wire N__39049;
    wire N__39046;
    wire N__39043;
    wire N__39038;
    wire N__39035;
    wire N__39030;
    wire N__39027;
    wire N__39024;
    wire N__39021;
    wire N__39018;
    wire N__39015;
    wire N__39012;
    wire N__39009;
    wire N__39006;
    wire N__39003;
    wire N__39000;
    wire N__38997;
    wire N__38994;
    wire N__38991;
    wire N__38988;
    wire N__38985;
    wire N__38982;
    wire N__38979;
    wire N__38976;
    wire N__38973;
    wire N__38970;
    wire N__38967;
    wire N__38964;
    wire N__38961;
    wire N__38958;
    wire N__38955;
    wire N__38952;
    wire N__38949;
    wire N__38946;
    wire N__38943;
    wire N__38940;
    wire N__38937;
    wire N__38934;
    wire N__38931;
    wire N__38928;
    wire N__38925;
    wire N__38922;
    wire N__38919;
    wire N__38916;
    wire N__38915;
    wire N__38912;
    wire N__38911;
    wire N__38908;
    wire N__38905;
    wire N__38902;
    wire N__38897;
    wire N__38894;
    wire N__38891;
    wire N__38890;
    wire N__38887;
    wire N__38884;
    wire N__38881;
    wire N__38874;
    wire N__38871;
    wire N__38868;
    wire N__38865;
    wire N__38862;
    wire N__38859;
    wire N__38856;
    wire N__38853;
    wire N__38850;
    wire N__38847;
    wire N__38844;
    wire N__38841;
    wire N__38838;
    wire N__38835;
    wire N__38832;
    wire N__38829;
    wire N__38828;
    wire N__38827;
    wire N__38822;
    wire N__38819;
    wire N__38816;
    wire N__38813;
    wire N__38810;
    wire N__38805;
    wire N__38802;
    wire N__38799;
    wire N__38798;
    wire N__38795;
    wire N__38792;
    wire N__38789;
    wire N__38784;
    wire N__38783;
    wire N__38780;
    wire N__38777;
    wire N__38774;
    wire N__38771;
    wire N__38766;
    wire N__38763;
    wire N__38760;
    wire N__38759;
    wire N__38756;
    wire N__38753;
    wire N__38750;
    wire N__38747;
    wire N__38742;
    wire N__38739;
    wire N__38736;
    wire N__38733;
    wire N__38730;
    wire N__38729;
    wire N__38726;
    wire N__38723;
    wire N__38720;
    wire N__38719;
    wire N__38716;
    wire N__38713;
    wire N__38710;
    wire N__38707;
    wire N__38702;
    wire N__38699;
    wire N__38696;
    wire N__38691;
    wire N__38690;
    wire N__38685;
    wire N__38682;
    wire N__38681;
    wire N__38678;
    wire N__38675;
    wire N__38672;
    wire N__38669;
    wire N__38666;
    wire N__38661;
    wire N__38660;
    wire N__38655;
    wire N__38652;
    wire N__38651;
    wire N__38646;
    wire N__38643;
    wire N__38640;
    wire N__38637;
    wire N__38634;
    wire N__38633;
    wire N__38632;
    wire N__38627;
    wire N__38624;
    wire N__38619;
    wire N__38616;
    wire N__38613;
    wire N__38610;
    wire N__38607;
    wire N__38606;
    wire N__38603;
    wire N__38600;
    wire N__38597;
    wire N__38594;
    wire N__38589;
    wire N__38586;
    wire N__38585;
    wire N__38580;
    wire N__38577;
    wire N__38574;
    wire N__38571;
    wire N__38570;
    wire N__38569;
    wire N__38566;
    wire N__38561;
    wire N__38558;
    wire N__38555;
    wire N__38552;
    wire N__38549;
    wire N__38544;
    wire N__38541;
    wire N__38538;
    wire N__38535;
    wire N__38534;
    wire N__38531;
    wire N__38528;
    wire N__38525;
    wire N__38522;
    wire N__38519;
    wire N__38514;
    wire N__38511;
    wire N__38510;
    wire N__38507;
    wire N__38506;
    wire N__38503;
    wire N__38502;
    wire N__38497;
    wire N__38492;
    wire N__38491;
    wire N__38486;
    wire N__38483;
    wire N__38478;
    wire N__38477;
    wire N__38472;
    wire N__38469;
    wire N__38466;
    wire N__38465;
    wire N__38464;
    wire N__38463;
    wire N__38462;
    wire N__38461;
    wire N__38460;
    wire N__38459;
    wire N__38454;
    wire N__38451;
    wire N__38450;
    wire N__38449;
    wire N__38448;
    wire N__38447;
    wire N__38444;
    wire N__38443;
    wire N__38442;
    wire N__38441;
    wire N__38440;
    wire N__38439;
    wire N__38430;
    wire N__38427;
    wire N__38414;
    wire N__38403;
    wire N__38402;
    wire N__38401;
    wire N__38400;
    wire N__38399;
    wire N__38398;
    wire N__38395;
    wire N__38388;
    wire N__38383;
    wire N__38378;
    wire N__38375;
    wire N__38374;
    wire N__38369;
    wire N__38368;
    wire N__38367;
    wire N__38366;
    wire N__38365;
    wire N__38362;
    wire N__38357;
    wire N__38354;
    wire N__38351;
    wire N__38348;
    wire N__38341;
    wire N__38338;
    wire N__38335;
    wire N__38322;
    wire N__38319;
    wire N__38316;
    wire N__38313;
    wire N__38310;
    wire N__38309;
    wire N__38306;
    wire N__38303;
    wire N__38300;
    wire N__38295;
    wire N__38292;
    wire N__38289;
    wire N__38286;
    wire N__38283;
    wire N__38280;
    wire N__38277;
    wire N__38274;
    wire N__38271;
    wire N__38268;
    wire N__38265;
    wire N__38262;
    wire N__38259;
    wire N__38256;
    wire N__38255;
    wire N__38252;
    wire N__38249;
    wire N__38244;
    wire N__38241;
    wire N__38238;
    wire N__38235;
    wire N__38232;
    wire N__38231;
    wire N__38228;
    wire N__38225;
    wire N__38222;
    wire N__38217;
    wire N__38214;
    wire N__38213;
    wire N__38210;
    wire N__38209;
    wire N__38206;
    wire N__38203;
    wire N__38202;
    wire N__38197;
    wire N__38194;
    wire N__38191;
    wire N__38184;
    wire N__38181;
    wire N__38178;
    wire N__38175;
    wire N__38174;
    wire N__38171;
    wire N__38168;
    wire N__38165;
    wire N__38160;
    wire N__38157;
    wire N__38154;
    wire N__38153;
    wire N__38152;
    wire N__38151;
    wire N__38148;
    wire N__38145;
    wire N__38140;
    wire N__38133;
    wire N__38130;
    wire N__38127;
    wire N__38126;
    wire N__38123;
    wire N__38120;
    wire N__38117;
    wire N__38114;
    wire N__38109;
    wire N__38106;
    wire N__38103;
    wire N__38102;
    wire N__38099;
    wire N__38096;
    wire N__38093;
    wire N__38090;
    wire N__38085;
    wire N__38082;
    wire N__38079;
    wire N__38078;
    wire N__38075;
    wire N__38072;
    wire N__38069;
    wire N__38064;
    wire N__38061;
    wire N__38058;
    wire N__38055;
    wire N__38054;
    wire N__38051;
    wire N__38048;
    wire N__38043;
    wire N__38040;
    wire N__38037;
    wire N__38034;
    wire N__38031;
    wire N__38030;
    wire N__38027;
    wire N__38024;
    wire N__38021;
    wire N__38016;
    wire N__38013;
    wire N__38010;
    wire N__38007;
    wire N__38006;
    wire N__38003;
    wire N__38000;
    wire N__37995;
    wire N__37992;
    wire N__37989;
    wire N__37986;
    wire N__37983;
    wire N__37980;
    wire N__37979;
    wire N__37976;
    wire N__37973;
    wire N__37968;
    wire N__37967;
    wire N__37962;
    wire N__37961;
    wire N__37958;
    wire N__37955;
    wire N__37952;
    wire N__37949;
    wire N__37946;
    wire N__37943;
    wire N__37938;
    wire N__37937;
    wire N__37932;
    wire N__37931;
    wire N__37928;
    wire N__37925;
    wire N__37922;
    wire N__37919;
    wire N__37916;
    wire N__37913;
    wire N__37908;
    wire N__37907;
    wire N__37902;
    wire N__37901;
    wire N__37898;
    wire N__37895;
    wire N__37892;
    wire N__37889;
    wire N__37886;
    wire N__37883;
    wire N__37878;
    wire N__37877;
    wire N__37874;
    wire N__37873;
    wire N__37868;
    wire N__37865;
    wire N__37862;
    wire N__37859;
    wire N__37856;
    wire N__37853;
    wire N__37850;
    wire N__37847;
    wire N__37842;
    wire N__37841;
    wire N__37840;
    wire N__37839;
    wire N__37836;
    wire N__37835;
    wire N__37834;
    wire N__37821;
    wire N__37818;
    wire N__37815;
    wire N__37814;
    wire N__37813;
    wire N__37812;
    wire N__37809;
    wire N__37806;
    wire N__37803;
    wire N__37800;
    wire N__37795;
    wire N__37790;
    wire N__37785;
    wire N__37782;
    wire N__37779;
    wire N__37776;
    wire N__37775;
    wire N__37774;
    wire N__37771;
    wire N__37770;
    wire N__37767;
    wire N__37764;
    wire N__37761;
    wire N__37760;
    wire N__37759;
    wire N__37756;
    wire N__37753;
    wire N__37750;
    wire N__37747;
    wire N__37744;
    wire N__37741;
    wire N__37738;
    wire N__37725;
    wire N__37722;
    wire N__37719;
    wire N__37718;
    wire N__37717;
    wire N__37714;
    wire N__37713;
    wire N__37712;
    wire N__37711;
    wire N__37710;
    wire N__37709;
    wire N__37708;
    wire N__37703;
    wire N__37700;
    wire N__37695;
    wire N__37694;
    wire N__37693;
    wire N__37684;
    wire N__37681;
    wire N__37678;
    wire N__37675;
    wire N__37670;
    wire N__37667;
    wire N__37664;
    wire N__37661;
    wire N__37658;
    wire N__37647;
    wire N__37646;
    wire N__37643;
    wire N__37642;
    wire N__37639;
    wire N__37638;
    wire N__37635;
    wire N__37632;
    wire N__37631;
    wire N__37630;
    wire N__37625;
    wire N__37624;
    wire N__37623;
    wire N__37620;
    wire N__37619;
    wire N__37618;
    wire N__37613;
    wire N__37610;
    wire N__37607;
    wire N__37604;
    wire N__37601;
    wire N__37598;
    wire N__37593;
    wire N__37590;
    wire N__37587;
    wire N__37584;
    wire N__37579;
    wire N__37576;
    wire N__37569;
    wire N__37566;
    wire N__37563;
    wire N__37560;
    wire N__37557;
    wire N__37548;
    wire N__37547;
    wire N__37546;
    wire N__37543;
    wire N__37540;
    wire N__37537;
    wire N__37536;
    wire N__37531;
    wire N__37528;
    wire N__37525;
    wire N__37522;
    wire N__37517;
    wire N__37512;
    wire N__37509;
    wire N__37508;
    wire N__37503;
    wire N__37500;
    wire N__37499;
    wire N__37494;
    wire N__37493;
    wire N__37490;
    wire N__37487;
    wire N__37484;
    wire N__37481;
    wire N__37478;
    wire N__37475;
    wire N__37470;
    wire N__37467;
    wire N__37464;
    wire N__37461;
    wire N__37458;
    wire N__37457;
    wire N__37456;
    wire N__37453;
    wire N__37448;
    wire N__37443;
    wire N__37440;
    wire N__37437;
    wire N__37434;
    wire N__37431;
    wire N__37428;
    wire N__37425;
    wire N__37422;
    wire N__37419;
    wire N__37416;
    wire N__37413;
    wire N__37410;
    wire N__37407;
    wire N__37404;
    wire N__37401;
    wire N__37398;
    wire N__37395;
    wire N__37392;
    wire N__37389;
    wire N__37386;
    wire N__37383;
    wire N__37382;
    wire N__37379;
    wire N__37376;
    wire N__37371;
    wire N__37368;
    wire N__37365;
    wire N__37362;
    wire N__37359;
    wire N__37356;
    wire N__37353;
    wire N__37352;
    wire N__37349;
    wire N__37346;
    wire N__37341;
    wire N__37338;
    wire N__37335;
    wire N__37332;
    wire N__37329;
    wire N__37326;
    wire N__37323;
    wire N__37322;
    wire N__37319;
    wire N__37316;
    wire N__37311;
    wire N__37310;
    wire N__37307;
    wire N__37304;
    wire N__37301;
    wire N__37296;
    wire N__37293;
    wire N__37290;
    wire N__37287;
    wire N__37284;
    wire N__37281;
    wire N__37280;
    wire N__37277;
    wire N__37274;
    wire N__37269;
    wire N__37266;
    wire N__37265;
    wire N__37262;
    wire N__37259;
    wire N__37258;
    wire N__37251;
    wire N__37248;
    wire N__37247;
    wire N__37244;
    wire N__37243;
    wire N__37242;
    wire N__37241;
    wire N__37240;
    wire N__37237;
    wire N__37226;
    wire N__37223;
    wire N__37218;
    wire N__37215;
    wire N__37212;
    wire N__37209;
    wire N__37206;
    wire N__37203;
    wire N__37202;
    wire N__37201;
    wire N__37198;
    wire N__37193;
    wire N__37190;
    wire N__37187;
    wire N__37184;
    wire N__37181;
    wire N__37176;
    wire N__37173;
    wire N__37172;
    wire N__37171;
    wire N__37168;
    wire N__37163;
    wire N__37160;
    wire N__37157;
    wire N__37152;
    wire N__37149;
    wire N__37146;
    wire N__37145;
    wire N__37144;
    wire N__37141;
    wire N__37136;
    wire N__37131;
    wire N__37128;
    wire N__37125;
    wire N__37122;
    wire N__37119;
    wire N__37116;
    wire N__37113;
    wire N__37110;
    wire N__37107;
    wire N__37104;
    wire N__37101;
    wire N__37098;
    wire N__37097;
    wire N__37096;
    wire N__37093;
    wire N__37090;
    wire N__37087;
    wire N__37082;
    wire N__37079;
    wire N__37076;
    wire N__37073;
    wire N__37068;
    wire N__37065;
    wire N__37062;
    wire N__37059;
    wire N__37058;
    wire N__37057;
    wire N__37054;
    wire N__37051;
    wire N__37048;
    wire N__37045;
    wire N__37042;
    wire N__37039;
    wire N__37036;
    wire N__37033;
    wire N__37030;
    wire N__37025;
    wire N__37022;
    wire N__37017;
    wire N__37014;
    wire N__37011;
    wire N__37010;
    wire N__37009;
    wire N__37006;
    wire N__37003;
    wire N__37000;
    wire N__36997;
    wire N__36994;
    wire N__36991;
    wire N__36988;
    wire N__36985;
    wire N__36982;
    wire N__36977;
    wire N__36974;
    wire N__36969;
    wire N__36966;
    wire N__36963;
    wire N__36960;
    wire N__36959;
    wire N__36956;
    wire N__36953;
    wire N__36952;
    wire N__36947;
    wire N__36944;
    wire N__36941;
    wire N__36938;
    wire N__36935;
    wire N__36932;
    wire N__36927;
    wire N__36924;
    wire N__36921;
    wire N__36918;
    wire N__36915;
    wire N__36914;
    wire N__36913;
    wire N__36910;
    wire N__36907;
    wire N__36904;
    wire N__36899;
    wire N__36896;
    wire N__36893;
    wire N__36890;
    wire N__36887;
    wire N__36884;
    wire N__36879;
    wire N__36876;
    wire N__36873;
    wire N__36872;
    wire N__36871;
    wire N__36868;
    wire N__36865;
    wire N__36862;
    wire N__36859;
    wire N__36856;
    wire N__36853;
    wire N__36850;
    wire N__36847;
    wire N__36840;
    wire N__36839;
    wire N__36836;
    wire N__36833;
    wire N__36830;
    wire N__36827;
    wire N__36824;
    wire N__36821;
    wire N__36818;
    wire N__36815;
    wire N__36810;
    wire N__36807;
    wire N__36804;
    wire N__36803;
    wire N__36802;
    wire N__36799;
    wire N__36796;
    wire N__36793;
    wire N__36790;
    wire N__36787;
    wire N__36784;
    wire N__36781;
    wire N__36778;
    wire N__36775;
    wire N__36770;
    wire N__36767;
    wire N__36762;
    wire N__36759;
    wire N__36756;
    wire N__36755;
    wire N__36752;
    wire N__36749;
    wire N__36746;
    wire N__36741;
    wire N__36738;
    wire N__36737;
    wire N__36736;
    wire N__36733;
    wire N__36730;
    wire N__36727;
    wire N__36722;
    wire N__36719;
    wire N__36716;
    wire N__36713;
    wire N__36710;
    wire N__36707;
    wire N__36702;
    wire N__36699;
    wire N__36696;
    wire N__36693;
    wire N__36692;
    wire N__36689;
    wire N__36686;
    wire N__36683;
    wire N__36678;
    wire N__36675;
    wire N__36674;
    wire N__36671;
    wire N__36670;
    wire N__36667;
    wire N__36664;
    wire N__36661;
    wire N__36658;
    wire N__36653;
    wire N__36650;
    wire N__36647;
    wire N__36644;
    wire N__36641;
    wire N__36638;
    wire N__36633;
    wire N__36630;
    wire N__36627;
    wire N__36626;
    wire N__36623;
    wire N__36620;
    wire N__36617;
    wire N__36612;
    wire N__36609;
    wire N__36608;
    wire N__36605;
    wire N__36604;
    wire N__36601;
    wire N__36598;
    wire N__36595;
    wire N__36592;
    wire N__36589;
    wire N__36586;
    wire N__36583;
    wire N__36580;
    wire N__36577;
    wire N__36574;
    wire N__36567;
    wire N__36564;
    wire N__36561;
    wire N__36558;
    wire N__36557;
    wire N__36554;
    wire N__36551;
    wire N__36548;
    wire N__36543;
    wire N__36540;
    wire N__36537;
    wire N__36536;
    wire N__36535;
    wire N__36532;
    wire N__36529;
    wire N__36526;
    wire N__36521;
    wire N__36518;
    wire N__36515;
    wire N__36512;
    wire N__36509;
    wire N__36506;
    wire N__36501;
    wire N__36498;
    wire N__36497;
    wire N__36496;
    wire N__36493;
    wire N__36490;
    wire N__36487;
    wire N__36484;
    wire N__36481;
    wire N__36478;
    wire N__36475;
    wire N__36470;
    wire N__36465;
    wire N__36462;
    wire N__36459;
    wire N__36456;
    wire N__36455;
    wire N__36454;
    wire N__36451;
    wire N__36448;
    wire N__36445;
    wire N__36440;
    wire N__36437;
    wire N__36434;
    wire N__36431;
    wire N__36428;
    wire N__36425;
    wire N__36420;
    wire N__36417;
    wire N__36414;
    wire N__36411;
    wire N__36410;
    wire N__36409;
    wire N__36406;
    wire N__36403;
    wire N__36400;
    wire N__36395;
    wire N__36392;
    wire N__36389;
    wire N__36386;
    wire N__36383;
    wire N__36380;
    wire N__36375;
    wire N__36372;
    wire N__36371;
    wire N__36370;
    wire N__36365;
    wire N__36362;
    wire N__36359;
    wire N__36356;
    wire N__36353;
    wire N__36348;
    wire N__36347;
    wire N__36344;
    wire N__36341;
    wire N__36338;
    wire N__36335;
    wire N__36330;
    wire N__36327;
    wire N__36324;
    wire N__36321;
    wire N__36318;
    wire N__36317;
    wire N__36314;
    wire N__36311;
    wire N__36306;
    wire N__36303;
    wire N__36300;
    wire N__36299;
    wire N__36296;
    wire N__36295;
    wire N__36292;
    wire N__36289;
    wire N__36286;
    wire N__36283;
    wire N__36280;
    wire N__36277;
    wire N__36274;
    wire N__36271;
    wire N__36266;
    wire N__36261;
    wire N__36258;
    wire N__36255;
    wire N__36252;
    wire N__36251;
    wire N__36250;
    wire N__36247;
    wire N__36244;
    wire N__36241;
    wire N__36236;
    wire N__36233;
    wire N__36230;
    wire N__36227;
    wire N__36224;
    wire N__36221;
    wire N__36216;
    wire N__36213;
    wire N__36210;
    wire N__36209;
    wire N__36206;
    wire N__36203;
    wire N__36198;
    wire N__36197;
    wire N__36192;
    wire N__36189;
    wire N__36186;
    wire N__36183;
    wire N__36180;
    wire N__36177;
    wire N__36174;
    wire N__36171;
    wire N__36168;
    wire N__36165;
    wire N__36162;
    wire N__36159;
    wire N__36156;
    wire N__36153;
    wire N__36152;
    wire N__36151;
    wire N__36146;
    wire N__36143;
    wire N__36140;
    wire N__36137;
    wire N__36134;
    wire N__36129;
    wire N__36126;
    wire N__36123;
    wire N__36120;
    wire N__36119;
    wire N__36116;
    wire N__36113;
    wire N__36110;
    wire N__36107;
    wire N__36102;
    wire N__36101;
    wire N__36096;
    wire N__36093;
    wire N__36092;
    wire N__36087;
    wire N__36084;
    wire N__36081;
    wire N__36078;
    wire N__36075;
    wire N__36072;
    wire N__36069;
    wire N__36066;
    wire N__36065;
    wire N__36064;
    wire N__36057;
    wire N__36054;
    wire N__36051;
    wire N__36048;
    wire N__36045;
    wire N__36042;
    wire N__36041;
    wire N__36036;
    wire N__36033;
    wire N__36030;
    wire N__36027;
    wire N__36026;
    wire N__36021;
    wire N__36018;
    wire N__36015;
    wire N__36012;
    wire N__36009;
    wire N__36006;
    wire N__36003;
    wire N__36000;
    wire N__35997;
    wire N__35994;
    wire N__35991;
    wire N__35990;
    wire N__35987;
    wire N__35984;
    wire N__35979;
    wire N__35978;
    wire N__35975;
    wire N__35972;
    wire N__35969;
    wire N__35966;
    wire N__35961;
    wire N__35958;
    wire N__35955;
    wire N__35952;
    wire N__35951;
    wire N__35948;
    wire N__35945;
    wire N__35942;
    wire N__35937;
    wire N__35936;
    wire N__35935;
    wire N__35932;
    wire N__35927;
    wire N__35924;
    wire N__35921;
    wire N__35918;
    wire N__35915;
    wire N__35912;
    wire N__35909;
    wire N__35906;
    wire N__35901;
    wire N__35898;
    wire N__35895;
    wire N__35892;
    wire N__35889;
    wire N__35886;
    wire N__35885;
    wire N__35884;
    wire N__35881;
    wire N__35876;
    wire N__35873;
    wire N__35870;
    wire N__35867;
    wire N__35864;
    wire N__35859;
    wire N__35856;
    wire N__35853;
    wire N__35852;
    wire N__35849;
    wire N__35846;
    wire N__35843;
    wire N__35838;
    wire N__35837;
    wire N__35836;
    wire N__35829;
    wire N__35826;
    wire N__35823;
    wire N__35820;
    wire N__35817;
    wire N__35814;
    wire N__35813;
    wire N__35808;
    wire N__35805;
    wire N__35804;
    wire N__35799;
    wire N__35796;
    wire N__35793;
    wire N__35790;
    wire N__35787;
    wire N__35784;
    wire N__35781;
    wire N__35780;
    wire N__35779;
    wire N__35778;
    wire N__35777;
    wire N__35774;
    wire N__35773;
    wire N__35760;
    wire N__35757;
    wire N__35756;
    wire N__35755;
    wire N__35754;
    wire N__35753;
    wire N__35752;
    wire N__35751;
    wire N__35750;
    wire N__35747;
    wire N__35734;
    wire N__35731;
    wire N__35728;
    wire N__35721;
    wire N__35718;
    wire N__35715;
    wire N__35712;
    wire N__35711;
    wire N__35708;
    wire N__35707;
    wire N__35700;
    wire N__35697;
    wire N__35694;
    wire N__35693;
    wire N__35688;
    wire N__35685;
    wire N__35682;
    wire N__35679;
    wire N__35678;
    wire N__35675;
    wire N__35672;
    wire N__35669;
    wire N__35666;
    wire N__35661;
    wire N__35660;
    wire N__35657;
    wire N__35654;
    wire N__35651;
    wire N__35648;
    wire N__35643;
    wire N__35642;
    wire N__35641;
    wire N__35640;
    wire N__35637;
    wire N__35632;
    wire N__35629;
    wire N__35624;
    wire N__35619;
    wire N__35616;
    wire N__35613;
    wire N__35610;
    wire N__35607;
    wire N__35604;
    wire N__35601;
    wire N__35598;
    wire N__35595;
    wire N__35594;
    wire N__35589;
    wire N__35586;
    wire N__35583;
    wire N__35580;
    wire N__35579;
    wire N__35578;
    wire N__35575;
    wire N__35570;
    wire N__35569;
    wire N__35568;
    wire N__35563;
    wire N__35558;
    wire N__35555;
    wire N__35550;
    wire N__35547;
    wire N__35544;
    wire N__35543;
    wire N__35540;
    wire N__35539;
    wire N__35532;
    wire N__35529;
    wire N__35526;
    wire N__35525;
    wire N__35524;
    wire N__35521;
    wire N__35518;
    wire N__35515;
    wire N__35510;
    wire N__35507;
    wire N__35504;
    wire N__35501;
    wire N__35496;
    wire N__35495;
    wire N__35490;
    wire N__35487;
    wire N__35484;
    wire N__35481;
    wire N__35478;
    wire N__35477;
    wire N__35472;
    wire N__35469;
    wire N__35466;
    wire N__35463;
    wire N__35462;
    wire N__35459;
    wire N__35454;
    wire N__35451;
    wire N__35448;
    wire N__35445;
    wire N__35444;
    wire N__35439;
    wire N__35436;
    wire N__35433;
    wire N__35430;
    wire N__35427;
    wire N__35424;
    wire N__35421;
    wire N__35420;
    wire N__35417;
    wire N__35414;
    wire N__35413;
    wire N__35410;
    wire N__35407;
    wire N__35404;
    wire N__35401;
    wire N__35398;
    wire N__35393;
    wire N__35388;
    wire N__35385;
    wire N__35382;
    wire N__35379;
    wire N__35376;
    wire N__35373;
    wire N__35370;
    wire N__35369;
    wire N__35368;
    wire N__35365;
    wire N__35360;
    wire N__35355;
    wire N__35352;
    wire N__35349;
    wire N__35346;
    wire N__35343;
    wire N__35342;
    wire N__35339;
    wire N__35336;
    wire N__35333;
    wire N__35328;
    wire N__35327;
    wire N__35322;
    wire N__35319;
    wire N__35316;
    wire N__35313;
    wire N__35310;
    wire N__35309;
    wire N__35304;
    wire N__35301;
    wire N__35300;
    wire N__35299;
    wire N__35292;
    wire N__35289;
    wire N__35286;
    wire N__35283;
    wire N__35280;
    wire N__35277;
    wire N__35274;
    wire N__35271;
    wire N__35268;
    wire N__35265;
    wire N__35262;
    wire N__35261;
    wire N__35260;
    wire N__35257;
    wire N__35252;
    wire N__35247;
    wire N__35244;
    wire N__35241;
    wire N__35238;
    wire N__35235;
    wire N__35234;
    wire N__35233;
    wire N__35230;
    wire N__35225;
    wire N__35222;
    wire N__35219;
    wire N__35214;
    wire N__35213;
    wire N__35212;
    wire N__35209;
    wire N__35206;
    wire N__35203;
    wire N__35200;
    wire N__35197;
    wire N__35192;
    wire N__35189;
    wire N__35186;
    wire N__35181;
    wire N__35180;
    wire N__35179;
    wire N__35178;
    wire N__35177;
    wire N__35174;
    wire N__35173;
    wire N__35170;
    wire N__35165;
    wire N__35158;
    wire N__35151;
    wire N__35150;
    wire N__35147;
    wire N__35144;
    wire N__35143;
    wire N__35142;
    wire N__35141;
    wire N__35140;
    wire N__35139;
    wire N__35134;
    wire N__35129;
    wire N__35122;
    wire N__35115;
    wire N__35112;
    wire N__35109;
    wire N__35106;
    wire N__35105;
    wire N__35104;
    wire N__35103;
    wire N__35100;
    wire N__35097;
    wire N__35094;
    wire N__35093;
    wire N__35092;
    wire N__35089;
    wire N__35084;
    wire N__35077;
    wire N__35072;
    wire N__35069;
    wire N__35066;
    wire N__35063;
    wire N__35058;
    wire N__35057;
    wire N__35056;
    wire N__35055;
    wire N__35054;
    wire N__35051;
    wire N__35046;
    wire N__35041;
    wire N__35034;
    wire N__35031;
    wire N__35028;
    wire N__35025;
    wire N__35022;
    wire N__35019;
    wire N__35018;
    wire N__35015;
    wire N__35012;
    wire N__35009;
    wire N__35006;
    wire N__35001;
    wire N__34998;
    wire N__34997;
    wire N__34994;
    wire N__34991;
    wire N__34986;
    wire N__34983;
    wire N__34982;
    wire N__34981;
    wire N__34978;
    wire N__34973;
    wire N__34968;
    wire N__34965;
    wire N__34962;
    wire N__34959;
    wire N__34958;
    wire N__34955;
    wire N__34952;
    wire N__34949;
    wire N__34946;
    wire N__34943;
    wire N__34938;
    wire N__34935;
    wire N__34932;
    wire N__34929;
    wire N__34926;
    wire N__34923;
    wire N__34920;
    wire N__34919;
    wire N__34914;
    wire N__34911;
    wire N__34908;
    wire N__34905;
    wire N__34902;
    wire N__34901;
    wire N__34898;
    wire N__34895;
    wire N__34892;
    wire N__34889;
    wire N__34886;
    wire N__34883;
    wire N__34878;
    wire N__34877;
    wire N__34874;
    wire N__34871;
    wire N__34868;
    wire N__34865;
    wire N__34862;
    wire N__34859;
    wire N__34856;
    wire N__34851;
    wire N__34848;
    wire N__34845;
    wire N__34844;
    wire N__34839;
    wire N__34836;
    wire N__34833;
    wire N__34830;
    wire N__34827;
    wire N__34824;
    wire N__34821;
    wire N__34820;
    wire N__34817;
    wire N__34814;
    wire N__34811;
    wire N__34808;
    wire N__34803;
    wire N__34802;
    wire N__34799;
    wire N__34796;
    wire N__34793;
    wire N__34788;
    wire N__34785;
    wire N__34782;
    wire N__34779;
    wire N__34776;
    wire N__34773;
    wire N__34770;
    wire N__34767;
    wire N__34764;
    wire N__34761;
    wire N__34758;
    wire N__34755;
    wire N__34754;
    wire N__34753;
    wire N__34750;
    wire N__34745;
    wire N__34740;
    wire N__34737;
    wire N__34734;
    wire N__34731;
    wire N__34728;
    wire N__34727;
    wire N__34722;
    wire N__34721;
    wire N__34718;
    wire N__34715;
    wire N__34712;
    wire N__34709;
    wire N__34706;
    wire N__34703;
    wire N__34698;
    wire N__34695;
    wire N__34694;
    wire N__34691;
    wire N__34688;
    wire N__34685;
    wire N__34680;
    wire N__34677;
    wire N__34674;
    wire N__34671;
    wire N__34668;
    wire N__34667;
    wire N__34664;
    wire N__34661;
    wire N__34656;
    wire N__34653;
    wire N__34650;
    wire N__34647;
    wire N__34644;
    wire N__34641;
    wire N__34638;
    wire N__34635;
    wire N__34632;
    wire N__34629;
    wire N__34626;
    wire N__34623;
    wire N__34620;
    wire N__34617;
    wire N__34614;
    wire N__34611;
    wire N__34610;
    wire N__34607;
    wire N__34604;
    wire N__34601;
    wire N__34596;
    wire N__34593;
    wire N__34590;
    wire N__34587;
    wire N__34584;
    wire N__34581;
    wire N__34578;
    wire N__34575;
    wire N__34572;
    wire N__34569;
    wire N__34566;
    wire N__34563;
    wire N__34560;
    wire N__34557;
    wire N__34554;
    wire N__34551;
    wire N__34548;
    wire N__34545;
    wire N__34542;
    wire N__34539;
    wire N__34536;
    wire N__34533;
    wire N__34530;
    wire N__34527;
    wire N__34524;
    wire N__34521;
    wire N__34518;
    wire N__34515;
    wire N__34512;
    wire N__34511;
    wire N__34510;
    wire N__34507;
    wire N__34502;
    wire N__34497;
    wire N__34496;
    wire N__34493;
    wire N__34490;
    wire N__34487;
    wire N__34484;
    wire N__34481;
    wire N__34478;
    wire N__34473;
    wire N__34470;
    wire N__34467;
    wire N__34464;
    wire N__34461;
    wire N__34458;
    wire N__34455;
    wire N__34452;
    wire N__34449;
    wire N__34446;
    wire N__34443;
    wire N__34440;
    wire N__34437;
    wire N__34434;
    wire N__34431;
    wire N__34428;
    wire N__34425;
    wire N__34422;
    wire N__34419;
    wire N__34416;
    wire N__34413;
    wire N__34410;
    wire N__34407;
    wire N__34404;
    wire N__34401;
    wire N__34398;
    wire N__34395;
    wire N__34392;
    wire N__34389;
    wire N__34386;
    wire N__34383;
    wire N__34380;
    wire N__34377;
    wire N__34374;
    wire N__34371;
    wire N__34368;
    wire N__34367;
    wire N__34364;
    wire N__34361;
    wire N__34356;
    wire N__34353;
    wire N__34350;
    wire N__34347;
    wire N__34344;
    wire N__34341;
    wire N__34338;
    wire N__34335;
    wire N__34332;
    wire N__34329;
    wire N__34326;
    wire N__34323;
    wire N__34320;
    wire N__34319;
    wire N__34316;
    wire N__34313;
    wire N__34310;
    wire N__34305;
    wire N__34302;
    wire N__34299;
    wire N__34296;
    wire N__34293;
    wire N__34290;
    wire N__34287;
    wire N__34284;
    wire N__34281;
    wire N__34278;
    wire N__34275;
    wire N__34272;
    wire N__34269;
    wire N__34266;
    wire N__34265;
    wire N__34262;
    wire N__34259;
    wire N__34254;
    wire N__34251;
    wire N__34248;
    wire N__34245;
    wire N__34242;
    wire N__34239;
    wire N__34238;
    wire N__34235;
    wire N__34232;
    wire N__34229;
    wire N__34226;
    wire N__34223;
    wire N__34218;
    wire N__34215;
    wire N__34214;
    wire N__34211;
    wire N__34210;
    wire N__34207;
    wire N__34202;
    wire N__34197;
    wire N__34196;
    wire N__34191;
    wire N__34188;
    wire N__34185;
    wire N__34184;
    wire N__34181;
    wire N__34178;
    wire N__34173;
    wire N__34170;
    wire N__34167;
    wire N__34164;
    wire N__34163;
    wire N__34160;
    wire N__34159;
    wire N__34158;
    wire N__34157;
    wire N__34154;
    wire N__34151;
    wire N__34148;
    wire N__34143;
    wire N__34134;
    wire N__34133;
    wire N__34130;
    wire N__34129;
    wire N__34128;
    wire N__34127;
    wire N__34124;
    wire N__34121;
    wire N__34118;
    wire N__34113;
    wire N__34104;
    wire N__34101;
    wire N__34100;
    wire N__34097;
    wire N__34096;
    wire N__34091;
    wire N__34088;
    wire N__34083;
    wire N__34080;
    wire N__34079;
    wire N__34074;
    wire N__34071;
    wire N__34070;
    wire N__34067;
    wire N__34064;
    wire N__34059;
    wire N__34058;
    wire N__34057;
    wire N__34056;
    wire N__34053;
    wire N__34050;
    wire N__34045;
    wire N__34042;
    wire N__34039;
    wire N__34032;
    wire N__34029;
    wire N__34026;
    wire N__34025;
    wire N__34022;
    wire N__34019;
    wire N__34014;
    wire N__34011;
    wire N__34010;
    wire N__34009;
    wire N__34002;
    wire N__33999;
    wire N__33996;
    wire N__33993;
    wire N__33990;
    wire N__33987;
    wire N__33984;
    wire N__33981;
    wire N__33980;
    wire N__33977;
    wire N__33974;
    wire N__33969;
    wire N__33966;
    wire N__33965;
    wire N__33962;
    wire N__33959;
    wire N__33954;
    wire N__33951;
    wire N__33948;
    wire N__33945;
    wire N__33942;
    wire N__33941;
    wire N__33940;
    wire N__33939;
    wire N__33936;
    wire N__33929;
    wire N__33924;
    wire N__33923;
    wire N__33918;
    wire N__33915;
    wire N__33912;
    wire N__33911;
    wire N__33910;
    wire N__33909;
    wire N__33906;
    wire N__33901;
    wire N__33898;
    wire N__33891;
    wire N__33890;
    wire N__33889;
    wire N__33886;
    wire N__33883;
    wire N__33880;
    wire N__33873;
    wire N__33872;
    wire N__33871;
    wire N__33870;
    wire N__33867;
    wire N__33864;
    wire N__33859;
    wire N__33852;
    wire N__33851;
    wire N__33848;
    wire N__33847;
    wire N__33846;
    wire N__33843;
    wire N__33838;
    wire N__33835;
    wire N__33828;
    wire N__33827;
    wire N__33826;
    wire N__33825;
    wire N__33822;
    wire N__33817;
    wire N__33814;
    wire N__33807;
    wire N__33806;
    wire N__33805;
    wire N__33802;
    wire N__33799;
    wire N__33796;
    wire N__33789;
    wire N__33788;
    wire N__33787;
    wire N__33784;
    wire N__33781;
    wire N__33778;
    wire N__33771;
    wire N__33770;
    wire N__33769;
    wire N__33766;
    wire N__33763;
    wire N__33760;
    wire N__33757;
    wire N__33754;
    wire N__33747;
    wire N__33746;
    wire N__33745;
    wire N__33742;
    wire N__33739;
    wire N__33736;
    wire N__33729;
    wire N__33726;
    wire N__33723;
    wire N__33720;
    wire N__33717;
    wire N__33714;
    wire N__33711;
    wire N__33708;
    wire N__33705;
    wire N__33702;
    wire N__33699;
    wire N__33696;
    wire N__33693;
    wire N__33690;
    wire N__33687;
    wire N__33684;
    wire N__33681;
    wire N__33678;
    wire N__33675;
    wire N__33672;
    wire N__33669;
    wire N__33666;
    wire N__33663;
    wire N__33660;
    wire N__33659;
    wire N__33656;
    wire N__33653;
    wire N__33650;
    wire N__33645;
    wire N__33644;
    wire N__33643;
    wire N__33642;
    wire N__33639;
    wire N__33630;
    wire N__33627;
    wire N__33626;
    wire N__33625;
    wire N__33622;
    wire N__33619;
    wire N__33616;
    wire N__33609;
    wire N__33608;
    wire N__33607;
    wire N__33604;
    wire N__33601;
    wire N__33598;
    wire N__33591;
    wire N__33588;
    wire N__33585;
    wire N__33582;
    wire N__33579;
    wire N__33578;
    wire N__33577;
    wire N__33574;
    wire N__33569;
    wire N__33564;
    wire N__33561;
    wire N__33558;
    wire N__33555;
    wire N__33552;
    wire N__33549;
    wire N__33546;
    wire N__33543;
    wire N__33540;
    wire N__33537;
    wire N__33536;
    wire N__33533;
    wire N__33530;
    wire N__33527;
    wire N__33524;
    wire N__33519;
    wire N__33516;
    wire N__33513;
    wire N__33510;
    wire N__33509;
    wire N__33508;
    wire N__33501;
    wire N__33498;
    wire N__33495;
    wire N__33492;
    wire N__33489;
    wire N__33486;
    wire N__33483;
    wire N__33482;
    wire N__33477;
    wire N__33474;
    wire N__33471;
    wire N__33468;
    wire N__33467;
    wire N__33466;
    wire N__33465;
    wire N__33464;
    wire N__33463;
    wire N__33462;
    wire N__33461;
    wire N__33460;
    wire N__33459;
    wire N__33458;
    wire N__33457;
    wire N__33456;
    wire N__33455;
    wire N__33454;
    wire N__33423;
    wire N__33420;
    wire N__33417;
    wire N__33414;
    wire N__33411;
    wire N__33408;
    wire N__33405;
    wire N__33404;
    wire N__33403;
    wire N__33400;
    wire N__33397;
    wire N__33394;
    wire N__33389;
    wire N__33386;
    wire N__33381;
    wire N__33378;
    wire N__33375;
    wire N__33374;
    wire N__33371;
    wire N__33368;
    wire N__33363;
    wire N__33362;
    wire N__33361;
    wire N__33358;
    wire N__33353;
    wire N__33350;
    wire N__33347;
    wire N__33342;
    wire N__33341;
    wire N__33340;
    wire N__33337;
    wire N__33332;
    wire N__33327;
    wire N__33324;
    wire N__33323;
    wire N__33320;
    wire N__33317;
    wire N__33316;
    wire N__33313;
    wire N__33310;
    wire N__33307;
    wire N__33304;
    wire N__33299;
    wire N__33296;
    wire N__33293;
    wire N__33290;
    wire N__33285;
    wire N__33284;
    wire N__33281;
    wire N__33278;
    wire N__33273;
    wire N__33270;
    wire N__33267;
    wire N__33264;
    wire N__33261;
    wire N__33258;
    wire N__33255;
    wire N__33252;
    wire N__33249;
    wire N__33246;
    wire N__33243;
    wire N__33240;
    wire N__33237;
    wire N__33234;
    wire N__33231;
    wire N__33228;
    wire N__33225;
    wire N__33222;
    wire N__33219;
    wire N__33216;
    wire N__33213;
    wire N__33210;
    wire N__33207;
    wire N__33204;
    wire N__33201;
    wire N__33198;
    wire N__33195;
    wire N__33192;
    wire N__33189;
    wire N__33186;
    wire N__33183;
    wire N__33180;
    wire N__33177;
    wire N__33174;
    wire N__33171;
    wire N__33168;
    wire N__33165;
    wire N__33162;
    wire N__33159;
    wire N__33156;
    wire N__33153;
    wire N__33150;
    wire N__33147;
    wire N__33144;
    wire N__33141;
    wire N__33138;
    wire N__33137;
    wire N__33132;
    wire N__33129;
    wire N__33126;
    wire N__33123;
    wire N__33120;
    wire N__33117;
    wire N__33114;
    wire N__33111;
    wire N__33108;
    wire N__33105;
    wire N__33102;
    wire N__33099;
    wire N__33096;
    wire N__33093;
    wire N__33090;
    wire N__33087;
    wire N__33084;
    wire N__33081;
    wire N__33078;
    wire N__33075;
    wire N__33072;
    wire N__33069;
    wire N__33066;
    wire N__33063;
    wire N__33060;
    wire N__33057;
    wire N__33054;
    wire N__33051;
    wire N__33048;
    wire N__33045;
    wire N__33042;
    wire N__33039;
    wire N__33036;
    wire N__33035;
    wire N__33034;
    wire N__33027;
    wire N__33024;
    wire N__33021;
    wire N__33018;
    wire N__33015;
    wire N__33012;
    wire N__33009;
    wire N__33006;
    wire N__33003;
    wire N__33000;
    wire N__32997;
    wire N__32994;
    wire N__32991;
    wire N__32988;
    wire N__32985;
    wire N__32982;
    wire N__32979;
    wire N__32976;
    wire N__32973;
    wire N__32970;
    wire N__32967;
    wire N__32964;
    wire N__32961;
    wire N__32958;
    wire N__32955;
    wire N__32952;
    wire N__32949;
    wire N__32946;
    wire N__32943;
    wire N__32942;
    wire N__32937;
    wire N__32934;
    wire N__32931;
    wire N__32928;
    wire N__32925;
    wire N__32924;
    wire N__32919;
    wire N__32916;
    wire N__32915;
    wire N__32914;
    wire N__32907;
    wire N__32904;
    wire N__32901;
    wire N__32898;
    wire N__32895;
    wire N__32892;
    wire N__32889;
    wire N__32888;
    wire N__32883;
    wire N__32880;
    wire N__32877;
    wire N__32874;
    wire N__32871;
    wire N__32868;
    wire N__32865;
    wire N__32862;
    wire N__32859;
    wire N__32856;
    wire N__32853;
    wire N__32850;
    wire N__32847;
    wire N__32844;
    wire N__32841;
    wire N__32838;
    wire N__32835;
    wire N__32832;
    wire N__32829;
    wire N__32826;
    wire N__32823;
    wire N__32820;
    wire N__32817;
    wire N__32814;
    wire N__32811;
    wire N__32808;
    wire N__32805;
    wire N__32802;
    wire N__32799;
    wire N__32796;
    wire N__32793;
    wire N__32790;
    wire N__32787;
    wire N__32784;
    wire N__32781;
    wire N__32778;
    wire N__32777;
    wire N__32776;
    wire N__32769;
    wire N__32766;
    wire N__32763;
    wire N__32760;
    wire N__32757;
    wire N__32754;
    wire N__32753;
    wire N__32748;
    wire N__32745;
    wire N__32742;
    wire N__32739;
    wire N__32738;
    wire N__32733;
    wire N__32730;
    wire N__32727;
    wire N__32726;
    wire N__32721;
    wire N__32718;
    wire N__32717;
    wire N__32712;
    wire N__32711;
    wire N__32708;
    wire N__32705;
    wire N__32700;
    wire N__32697;
    wire N__32694;
    wire N__32691;
    wire N__32688;
    wire N__32687;
    wire N__32684;
    wire N__32681;
    wire N__32678;
    wire N__32673;
    wire N__32670;
    wire N__32667;
    wire N__32664;
    wire N__32661;
    wire N__32658;
    wire N__32655;
    wire N__32654;
    wire N__32651;
    wire N__32648;
    wire N__32645;
    wire N__32642;
    wire N__32639;
    wire N__32634;
    wire N__32631;
    wire N__32628;
    wire N__32627;
    wire N__32626;
    wire N__32625;
    wire N__32616;
    wire N__32613;
    wire N__32610;
    wire N__32607;
    wire N__32606;
    wire N__32605;
    wire N__32602;
    wire N__32597;
    wire N__32592;
    wire N__32589;
    wire N__32588;
    wire N__32583;
    wire N__32580;
    wire N__32577;
    wire N__32576;
    wire N__32573;
    wire N__32570;
    wire N__32565;
    wire N__32564;
    wire N__32563;
    wire N__32558;
    wire N__32555;
    wire N__32552;
    wire N__32549;
    wire N__32546;
    wire N__32541;
    wire N__32538;
    wire N__32537;
    wire N__32534;
    wire N__32531;
    wire N__32526;
    wire N__32523;
    wire N__32520;
    wire N__32517;
    wire N__32514;
    wire N__32513;
    wire N__32510;
    wire N__32507;
    wire N__32504;
    wire N__32499;
    wire N__32498;
    wire N__32495;
    wire N__32492;
    wire N__32489;
    wire N__32486;
    wire N__32483;
    wire N__32478;
    wire N__32477;
    wire N__32476;
    wire N__32473;
    wire N__32470;
    wire N__32467;
    wire N__32464;
    wire N__32459;
    wire N__32456;
    wire N__32453;
    wire N__32450;
    wire N__32445;
    wire N__32444;
    wire N__32439;
    wire N__32436;
    wire N__32433;
    wire N__32430;
    wire N__32427;
    wire N__32426;
    wire N__32425;
    wire N__32418;
    wire N__32415;
    wire N__32412;
    wire N__32411;
    wire N__32406;
    wire N__32403;
    wire N__32400;
    wire N__32397;
    wire N__32394;
    wire N__32391;
    wire N__32388;
    wire N__32385;
    wire N__32382;
    wire N__32379;
    wire N__32378;
    wire N__32375;
    wire N__32372;
    wire N__32371;
    wire N__32368;
    wire N__32365;
    wire N__32362;
    wire N__32359;
    wire N__32356;
    wire N__32349;
    wire N__32346;
    wire N__32345;
    wire N__32340;
    wire N__32337;
    wire N__32334;
    wire N__32331;
    wire N__32328;
    wire N__32325;
    wire N__32322;
    wire N__32319;
    wire N__32316;
    wire N__32313;
    wire N__32310;
    wire N__32307;
    wire N__32304;
    wire N__32301;
    wire N__32298;
    wire N__32295;
    wire N__32292;
    wire N__32289;
    wire N__32286;
    wire N__32283;
    wire N__32280;
    wire N__32277;
    wire N__32274;
    wire N__32271;
    wire N__32268;
    wire N__32265;
    wire N__32262;
    wire N__32259;
    wire N__32256;
    wire N__32253;
    wire N__32250;
    wire N__32247;
    wire N__32244;
    wire N__32241;
    wire N__32238;
    wire N__32235;
    wire N__32232;
    wire N__32229;
    wire N__32226;
    wire N__32223;
    wire N__32220;
    wire N__32217;
    wire N__32214;
    wire N__32211;
    wire N__32208;
    wire N__32205;
    wire N__32202;
    wire N__32199;
    wire N__32196;
    wire N__32193;
    wire N__32190;
    wire N__32187;
    wire N__32184;
    wire N__32181;
    wire N__32178;
    wire N__32175;
    wire N__32172;
    wire N__32169;
    wire N__32166;
    wire N__32163;
    wire N__32160;
    wire N__32157;
    wire N__32154;
    wire N__32151;
    wire N__32148;
    wire N__32145;
    wire N__32142;
    wire N__32139;
    wire N__32136;
    wire N__32133;
    wire N__32130;
    wire N__32127;
    wire N__32124;
    wire N__32121;
    wire N__32118;
    wire N__32115;
    wire N__32112;
    wire N__32109;
    wire N__32106;
    wire N__32103;
    wire N__32100;
    wire N__32097;
    wire N__32094;
    wire N__32091;
    wire N__32088;
    wire N__32085;
    wire N__32082;
    wire N__32079;
    wire N__32076;
    wire N__32073;
    wire N__32070;
    wire N__32067;
    wire N__32064;
    wire N__32061;
    wire N__32058;
    wire N__32055;
    wire N__32052;
    wire N__32049;
    wire N__32046;
    wire N__32043;
    wire N__32040;
    wire N__32037;
    wire N__32034;
    wire N__32031;
    wire N__32028;
    wire N__32025;
    wire N__32024;
    wire N__32019;
    wire N__32016;
    wire N__32013;
    wire N__32010;
    wire N__32007;
    wire N__32004;
    wire N__32001;
    wire N__31998;
    wire N__31995;
    wire N__31992;
    wire N__31989;
    wire N__31986;
    wire N__31983;
    wire N__31980;
    wire N__31977;
    wire N__31976;
    wire N__31971;
    wire N__31968;
    wire N__31965;
    wire N__31962;
    wire N__31959;
    wire N__31956;
    wire N__31953;
    wire N__31950;
    wire N__31947;
    wire N__31944;
    wire N__31941;
    wire N__31938;
    wire N__31935;
    wire N__31932;
    wire N__31929;
    wire N__31926;
    wire N__31923;
    wire N__31920;
    wire N__31917;
    wire N__31914;
    wire N__31913;
    wire N__31908;
    wire N__31905;
    wire N__31902;
    wire N__31899;
    wire N__31896;
    wire N__31893;
    wire N__31892;
    wire N__31887;
    wire N__31884;
    wire N__31881;
    wire N__31878;
    wire N__31875;
    wire N__31872;
    wire N__31869;
    wire N__31866;
    wire N__31863;
    wire N__31860;
    wire N__31857;
    wire N__31854;
    wire N__31853;
    wire N__31848;
    wire N__31845;
    wire N__31844;
    wire N__31843;
    wire N__31840;
    wire N__31835;
    wire N__31830;
    wire N__31827;
    wire N__31824;
    wire N__31821;
    wire N__31818;
    wire N__31815;
    wire N__31812;
    wire N__31809;
    wire N__31806;
    wire N__31805;
    wire N__31800;
    wire N__31797;
    wire N__31796;
    wire N__31795;
    wire N__31788;
    wire N__31785;
    wire N__31782;
    wire N__31779;
    wire N__31776;
    wire N__31773;
    wire N__31770;
    wire N__31767;
    wire N__31764;
    wire N__31761;
    wire N__31758;
    wire N__31755;
    wire N__31752;
    wire N__31749;
    wire N__31746;
    wire N__31743;
    wire N__31742;
    wire N__31737;
    wire N__31734;
    wire N__31733;
    wire N__31732;
    wire N__31725;
    wire N__31722;
    wire N__31719;
    wire N__31716;
    wire N__31713;
    wire N__31710;
    wire N__31707;
    wire N__31704;
    wire N__31701;
    wire N__31698;
    wire N__31695;
    wire N__31692;
    wire N__31689;
    wire N__31686;
    wire N__31683;
    wire N__31680;
    wire N__31677;
    wire N__31674;
    wire N__31671;
    wire N__31668;
    wire N__31665;
    wire N__31662;
    wire N__31659;
    wire N__31656;
    wire N__31653;
    wire N__31650;
    wire N__31647;
    wire N__31644;
    wire N__31641;
    wire N__31638;
    wire N__31635;
    wire N__31632;
    wire N__31629;
    wire N__31626;
    wire N__31623;
    wire N__31620;
    wire N__31617;
    wire N__31614;
    wire N__31611;
    wire N__31608;
    wire N__31605;
    wire N__31602;
    wire N__31599;
    wire N__31596;
    wire N__31593;
    wire N__31590;
    wire N__31587;
    wire N__31584;
    wire N__31581;
    wire N__31578;
    wire N__31575;
    wire N__31572;
    wire N__31569;
    wire N__31566;
    wire N__31563;
    wire N__31560;
    wire N__31557;
    wire N__31554;
    wire N__31551;
    wire N__31548;
    wire N__31545;
    wire N__31542;
    wire N__31539;
    wire N__31536;
    wire N__31533;
    wire N__31530;
    wire N__31527;
    wire N__31524;
    wire N__31521;
    wire N__31518;
    wire N__31515;
    wire N__31512;
    wire N__31509;
    wire N__31506;
    wire N__31503;
    wire N__31500;
    wire N__31497;
    wire N__31494;
    wire N__31491;
    wire N__31488;
    wire N__31485;
    wire N__31482;
    wire N__31479;
    wire N__31476;
    wire N__31473;
    wire N__31470;
    wire N__31467;
    wire N__31464;
    wire N__31461;
    wire N__31458;
    wire N__31455;
    wire N__31452;
    wire N__31449;
    wire N__31446;
    wire N__31443;
    wire N__31440;
    wire N__31437;
    wire N__31434;
    wire N__31431;
    wire N__31428;
    wire N__31425;
    wire N__31422;
    wire N__31419;
    wire N__31416;
    wire N__31413;
    wire N__31410;
    wire N__31407;
    wire N__31404;
    wire N__31401;
    wire N__31398;
    wire N__31395;
    wire N__31392;
    wire N__31389;
    wire N__31386;
    wire N__31383;
    wire N__31380;
    wire N__31377;
    wire N__31374;
    wire N__31371;
    wire N__31368;
    wire N__31365;
    wire N__31362;
    wire N__31359;
    wire N__31356;
    wire N__31353;
    wire N__31350;
    wire N__31347;
    wire N__31344;
    wire N__31341;
    wire N__31338;
    wire N__31335;
    wire N__31332;
    wire N__31329;
    wire N__31326;
    wire N__31323;
    wire N__31320;
    wire N__31317;
    wire N__31314;
    wire N__31311;
    wire N__31308;
    wire N__31305;
    wire N__31302;
    wire N__31299;
    wire N__31296;
    wire N__31293;
    wire N__31290;
    wire N__31287;
    wire N__31284;
    wire N__31281;
    wire N__31278;
    wire N__31275;
    wire N__31272;
    wire N__31269;
    wire N__31266;
    wire N__31263;
    wire N__31260;
    wire N__31257;
    wire N__31254;
    wire N__31251;
    wire N__31248;
    wire N__31245;
    wire \Pc2drone_pll_inst.clk_system_pll ;
    wire GNDG0;
    wire VCCG0;
    wire \pid_alt.O_4_11 ;
    wire \pid_alt.O_3_21 ;
    wire \pid_alt.O_3_18 ;
    wire \pid_alt.O_3_11 ;
    wire \pid_alt.O_3_15 ;
    wire \pid_alt.O_3_17 ;
    wire \pid_alt.O_3_24 ;
    wire \pid_alt.O_3_20 ;
    wire \pid_alt.O_3_22 ;
    wire \pid_alt.O_3_23 ;
    wire \pid_alt.O_3_19 ;
    wire \pid_alt.O_3_8 ;
    wire \pid_alt.O_3_7 ;
    wire \pid_alt.O_3_10 ;
    wire \pid_alt.O_3_9 ;
    wire \pid_alt.O_3_14 ;
    wire \pid_alt.O_3_13 ;
    wire \pid_alt.O_3_6 ;
    wire \pid_alt.O_3_5 ;
    wire \pid_alt.O_3_12 ;
    wire \pid_alt.O_4_12 ;
    wire \pid_alt.O_4_13 ;
    wire \pid_alt.O_4_10 ;
    wire \pid_alt.O_4_15 ;
    wire \pid_alt.O_4_16 ;
    wire \pid_alt.O_4_17 ;
    wire \pid_alt.O_4_18 ;
    wire \pid_alt.O_4_19 ;
    wire \pid_alt.O_4_20 ;
    wire \pid_alt.O_4_21 ;
    wire \pid_alt.O_4_22 ;
    wire \pid_alt.O_4_23 ;
    wire \pid_alt.O_4_6 ;
    wire \pid_alt.O_4_24 ;
    wire \pid_alt.O_4_7 ;
    wire \pid_alt.O_4_8 ;
    wire \pid_alt.O_4_9 ;
    wire \pid_alt.O_4_14 ;
    wire \pid_alt.O_4_4 ;
    wire \pid_alt.O_5_4 ;
    wire \pid_alt.O_4_5 ;
    wire \pid_alt.O_3_4 ;
    wire \pid_front.O_0_14 ;
    wire \pid_front.O_0_15 ;
    wire \pid_front.O_0_16 ;
    wire \pid_front.O_0_17 ;
    wire \pid_front.O_0_18 ;
    wire \pid_front.O_0_19 ;
    wire \pid_front.O_0_10 ;
    wire \pid_front.O_0_21 ;
    wire \pid_front.O_0_22 ;
    wire \pid_front.O_0_5 ;
    wire \pid_front.O_0_23 ;
    wire \pid_front.O_0_24 ;
    wire \pid_front.O_0_11 ;
    wire \pid_front.O_0_7 ;
    wire \pid_front.O_0_8 ;
    wire \pid_front.O_0_9 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIGDHM_0Z0Z_11_cascade_ ;
    wire \pid_alt.error_d_reg_prev_esr_RNIDAHMZ0Z_10 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIGDHM_0Z0Z_11 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIDAHMZ0Z_10_cascade_ ;
    wire \pid_alt.error_d_reg_prevZ0Z_10 ;
    wire \pid_alt.error_d_regZ0Z_10 ;
    wire \pid_alt.error_d_reg_prevZ0Z_11 ;
    wire \pid_alt.error_d_regZ0Z_11 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI86IM_0Z0Z_19_cascade_ ;
    wire \pid_alt.error_d_reg_prev_esr_RNI53IMZ0Z_18 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI86IM_0Z0Z_19 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI53IMZ0Z_18_cascade_ ;
    wire \pid_alt.error_d_reg_prevZ0Z_18 ;
    wire \pid_alt.error_d_regZ0Z_18 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI53IM_0Z0Z_18 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI53IM_0Z0Z_18_cascade_ ;
    wire \pid_alt.error_d_reg_prev_esr_RNII5611Z0Z_8_cascade_ ;
    wire \pid_alt.error_d_reg_prev_esr_RNIL8611_0Z0Z_9 ;
    wire \pid_alt.error_d_reg_prev_esr_RNII5611Z0Z_8 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIL8611_0Z0Z_9_cascade_ ;
    wire \pid_alt.O_5_6 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI20IMZ0Z_17 ;
    wire \pid_alt.O_5_21 ;
    wire \pid_alt.O_5_8 ;
    wire \pid_alt.O_5_24 ;
    wire \pid_alt.O_5_16 ;
    wire \pid_alt.O_5_14 ;
    wire \pid_alt.error_p_regZ0Z_10 ;
    wire \pid_alt.O_5_15 ;
    wire \pid_alt.error_p_regZ0Z_11 ;
    wire \pid_alt.O_5_19 ;
    wire \pid_alt.O_5_13 ;
    wire \pid_alt.O_5_17 ;
    wire \pid_alt.O_5_18 ;
    wire \pid_alt.O_5_22 ;
    wire \pid_alt.error_p_regZ0Z_18 ;
    wire \pid_alt.O_5_9 ;
    wire \pid_alt.O_5_10 ;
    wire \pid_alt.O_5_11 ;
    wire \pid_alt.O_5_23 ;
    wire \pid_alt.O_5_20 ;
    wire \pid_alt.O_3_16 ;
    wire alt_kd_1;
    wire alt_kd_4;
    wire alt_kd_3;
    wire alt_kd_5;
    wire alt_kd_6;
    wire alt_kd_2;
    wire alt_kd_7;
    wire \Commands_frame_decoder.WDTZ0Z_0 ;
    wire bfn_2_9_0_;
    wire \Commands_frame_decoder.WDTZ0Z_1 ;
    wire \Commands_frame_decoder.un1_WDT_cry_0 ;
    wire \Commands_frame_decoder.WDTZ0Z_2 ;
    wire \Commands_frame_decoder.un1_WDT_cry_1 ;
    wire \Commands_frame_decoder.WDTZ0Z_3 ;
    wire \Commands_frame_decoder.un1_WDT_cry_2 ;
    wire \Commands_frame_decoder.un1_WDT_cry_3 ;
    wire \Commands_frame_decoder.un1_WDT_cry_4 ;
    wire \Commands_frame_decoder.un1_WDT_cry_5 ;
    wire \Commands_frame_decoder.un1_WDT_cry_6 ;
    wire \Commands_frame_decoder.un1_WDT_cry_7 ;
    wire bfn_2_10_0_;
    wire \Commands_frame_decoder.un1_WDT_cry_8 ;
    wire \Commands_frame_decoder.un1_WDT_cry_9 ;
    wire \Commands_frame_decoder.un1_WDT_cry_10 ;
    wire \Commands_frame_decoder.un1_WDT_cry_11 ;
    wire \Commands_frame_decoder.un1_WDT_cry_12 ;
    wire \Commands_frame_decoder.un1_WDT_cry_13 ;
    wire \Commands_frame_decoder.un1_WDT_cry_14 ;
    wire alt_ki_0;
    wire alt_ki_1;
    wire alt_ki_2;
    wire alt_ki_3;
    wire alt_ki_4;
    wire alt_ki_5;
    wire alt_ki_6;
    wire alt_ki_7;
    wire \Commands_frame_decoder.state_ns_0_a3_0_1_cascade_ ;
    wire \Commands_frame_decoder.state_ns_i_a2_2_1Z0Z_0_cascade_ ;
    wire \Commands_frame_decoder.N_410_cascade_ ;
    wire xy_kp_4;
    wire \Commands_frame_decoder.source_CH3data_1_sqmuxa_cascade_ ;
    wire \Commands_frame_decoder.stateZ0Z_5 ;
    wire \pid_alt.error_p_reg_esr_RNIOI4PZ0Z_0_cascade_ ;
    wire \pid_alt.error_d_reg_prevZ0Z_0 ;
    wire \pid_alt.error_d_regZ0Z_0 ;
    wire \pid_alt.error_p_regZ0Z_0 ;
    wire \pid_alt.error_d_reg_prev_esr_RNITF511Z0Z_1 ;
    wire \pid_alt.error_d_reg_prev_esr_RNITF511_0Z0Z_1_cascade_ ;
    wire \pid_alt.error_p_regZ0Z_2 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI0J511_0Z0Z_2 ;
    wire \pid_alt.error_d_regZ0Z_1 ;
    wire \pid_alt.error_d_reg_prevZ0Z_1 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI0J511_0Z0Z_2_cascade_ ;
    wire \pid_alt.error_p_reg_esr_RNIOI4PZ0Z_0 ;
    wire \pid_alt.un1_pid_prereg_16_0_cascade_ ;
    wire \pid_alt.error_d_reg_prev_esr_RNITF511_0Z0Z_1 ;
    wire \pid_alt.error_d_regZ0Z_2 ;
    wire \pid_alt.error_d_reg_prevZ0Z_2 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI3M511Z0Z_3 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI3M511Z0Z_3_cascade_ ;
    wire \pid_alt.error_p_regZ0Z_4 ;
    wire \pid_alt.error_d_reg_prevZ0Z_4 ;
    wire \pid_alt.error_d_regZ0Z_4 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI6P511_0Z0Z_4 ;
    wire \pid_alt.error_d_regZ0Z_3 ;
    wire \pid_alt.error_d_reg_prevZ0Z_3 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI3M511_0Z0Z_3 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI0J511Z0Z_2 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI3M511_0Z0Z_3_cascade_ ;
    wire \pid_alt.error_d_reg_prev_esr_RNII5LS3Z0Z_1 ;
    wire \pid_alt.error_d_regZ0Z_8 ;
    wire \pid_alt.error_d_reg_prevZ0Z_8 ;
    wire \pid_alt.error_d_reg_prev_esr_RNII5611_0Z0Z_8_cascade_ ;
    wire \pid_alt.error_d_reg_prev_esr_RNIF2611Z0Z_7 ;
    wire \pid_alt.error_d_reg_prev_esr_RNII5611_0Z0Z_8 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIF2611Z0Z_7_cascade_ ;
    wire \pid_alt.error_p_regZ0Z_7 ;
    wire \pid_alt.error_d_reg_prevZ0Z_7 ;
    wire \pid_alt.error_d_regZ0Z_7 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIF2611_0Z0Z_7 ;
    wire \pid_alt.error_d_reg_prev_esr_RNICV511Z0Z_6 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIF2611_0Z0Z_7_cascade_ ;
    wire bfn_2_18_0_;
    wire \pid_alt.error_i_regZ0Z_1 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_0 ;
    wire \pid_alt.error_i_regZ0Z_2 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_1 ;
    wire \pid_alt.error_i_regZ0Z_3 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_2 ;
    wire \pid_alt.error_i_regZ0Z_4 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_3 ;
    wire \pid_alt.error_i_regZ0Z_5 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_4 ;
    wire \pid_alt.error_i_regZ0Z_6 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_5 ;
    wire \pid_alt.error_i_regZ0Z_7 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_6 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_7 ;
    wire \pid_alt.error_i_regZ0Z_8 ;
    wire bfn_2_19_0_;
    wire \pid_alt.error_i_regZ0Z_9 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_8_c_RNI9POQ ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_8 ;
    wire \pid_alt.error_i_regZ0Z_10 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_9 ;
    wire \pid_alt.error_i_regZ0Z_11 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_10 ;
    wire \pid_alt.error_i_regZ0Z_12 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_11 ;
    wire \pid_alt.error_i_regZ0Z_13 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_12 ;
    wire \pid_alt.error_i_regZ0Z_14 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_13 ;
    wire \pid_alt.error_i_regZ0Z_15 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_14 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_15 ;
    wire \pid_alt.error_i_regZ0Z_16 ;
    wire bfn_2_20_0_;
    wire \pid_alt.error_i_regZ0Z_17 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_16 ;
    wire \pid_alt.error_i_regZ0Z_18 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_17 ;
    wire \pid_alt.error_i_regZ0Z_19 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_18 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_19 ;
    wire \pid_alt.error_i_regZ0Z_20 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_20 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_20_c_RNISVKK_cascade_ ;
    wire \pid_alt.error_p_regZ0Z_17 ;
    wire \pid_alt.error_i_reg_esr_RNI4NMPZ0Z_11 ;
    wire \pid_alt.error_i_reg_esr_RNI9HOJZ0Z_18 ;
    wire \pid_alt.error_d_regZ0Z_17 ;
    wire \pid_alt.error_d_reg_prevZ0Z_17 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_18 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_20 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_17 ;
    wire \pid_alt.m7_e_4_cascade_ ;
    wire \pid_alt.N_545_cascade_ ;
    wire \pid_alt.error_i_acumm_preregZ0Z_16 ;
    wire \pid_alt.error_i_reg_esr_RNIBKPJZ0Z_19 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_19 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_14 ;
    wire \pid_alt.O_5_12 ;
    wire \pid_alt.error_p_regZ0Z_8 ;
    wire \pid_alt.O_5_5 ;
    wire \pid_alt.error_p_regZ0Z_1 ;
    wire \pid_alt.O_5_7 ;
    wire \pid_alt.error_p_regZ0Z_3 ;
    wire \pid_alt.N_939_0_g ;
    wire alt_kd_0;
    wire \Commands_frame_decoder.state_RNIRSI31Z0Z_11 ;
    wire \Commands_frame_decoder.WDT8lto9_3_cascade_ ;
    wire \Commands_frame_decoder.state_0_sqmuxacf0_1 ;
    wire \Commands_frame_decoder.state_0_sqmuxacf1 ;
    wire \Commands_frame_decoder.state_0_sqmuxacf0_cascade_ ;
    wire \Commands_frame_decoder.WDT8lt12_0 ;
    wire \Commands_frame_decoder.state_0_sqmuxa ;
    wire \Commands_frame_decoder.preinitZ0 ;
    wire \Commands_frame_decoder.WDTZ0Z_8 ;
    wire \Commands_frame_decoder.WDTZ0Z_9 ;
    wire \Commands_frame_decoder.WDTZ0Z_10 ;
    wire \Commands_frame_decoder.WDTZ0Z_13 ;
    wire \Commands_frame_decoder.WDTZ0Z_12 ;
    wire \Commands_frame_decoder.WDTZ0Z_11 ;
    wire \Commands_frame_decoder.WDTZ0Z_6 ;
    wire \Commands_frame_decoder.WDTZ0Z_5 ;
    wire \Commands_frame_decoder.WDTZ0Z_7 ;
    wire \Commands_frame_decoder.WDTZ0Z_4 ;
    wire \Commands_frame_decoder.WDT_RNI2VDI1Z0Z_10 ;
    wire \Commands_frame_decoder.WDT_RNITK4LZ0Z_8 ;
    wire \Commands_frame_decoder.WDT_RNIET8A1Z0Z_4_cascade_ ;
    wire \Commands_frame_decoder.WDT_RNIHV6PZ0Z_11 ;
    wire \Commands_frame_decoder.WDT8lt14_0_cascade_ ;
    wire \Commands_frame_decoder.state_RNIQRI31Z0Z_10 ;
    wire \Commands_frame_decoder.count_1_sqmuxa ;
    wire \Commands_frame_decoder.un1_state57_iZ0 ;
    wire \Commands_frame_decoder.countZ0Z_0 ;
    wire \Commands_frame_decoder.N_370_2 ;
    wire \Commands_frame_decoder.N_371 ;
    wire \Commands_frame_decoder.N_370_2_cascade_ ;
    wire \Commands_frame_decoder.N_365_0 ;
    wire \Commands_frame_decoder.state_ns_i_0_0_cascade_ ;
    wire \Commands_frame_decoder.stateZ0Z_0 ;
    wire \Commands_frame_decoder.state_ns_0_a3_3_1 ;
    wire \Commands_frame_decoder.stateZ0Z_1 ;
    wire \Commands_frame_decoder.N_372 ;
    wire \Commands_frame_decoder.stateZ0Z_14 ;
    wire \Commands_frame_decoder.stateZ0Z_13 ;
    wire \Commands_frame_decoder.N_410 ;
    wire \Commands_frame_decoder.N_406 ;
    wire \Commands_frame_decoder.WDT8lt14_0 ;
    wire \Commands_frame_decoder.WDTZ0Z_14 ;
    wire \Commands_frame_decoder.WDTZ0Z_15 ;
    wire \Commands_frame_decoder.N_403_cascade_ ;
    wire \Commands_frame_decoder.stateZ0Z_11 ;
    wire \Commands_frame_decoder.stateZ0Z_8 ;
    wire \Commands_frame_decoder.stateZ0Z_9 ;
    wire \Commands_frame_decoder.stateZ0Z_7 ;
    wire \pid_alt.source_pid_1_sqmuxa_0_a2_2_5_cascade_ ;
    wire \pid_alt.N_539_cascade_ ;
    wire \pid_alt.source_pid_9_0_0_4_cascade_ ;
    wire \pid_alt.source_pid_1_sqmuxa_0_a2_2_6 ;
    wire \pid_alt.error_d_reg_prev_i_0 ;
    wire bfn_3_15_0_;
    wire \pid_alt.error_p_reg_esr_RNI3SMI1Z0Z_0 ;
    wire \pid_alt.un1_pid_prereg_0 ;
    wire \pid_alt.un1_pid_prereg_un1_pid_prereg_0_cry_0_c_THRU_CO ;
    wire \pid_alt.error_d_reg_prev_esr_RNIFPN33Z0Z_1 ;
    wire \pid_alt.un1_pid_prereg_0_cry_0 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIF0465Z0Z_1 ;
    wire \pid_alt.un1_pid_prereg_0_cry_1 ;
    wire \pid_alt.error_d_reg_prev_esr_RNILDG87Z0Z_2 ;
    wire \pid_alt.un1_pid_prereg_0_cry_2 ;
    wire \pid_alt.error_d_reg_prev_esr_RNILE0V5Z0Z_2 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI11TA9Z0Z_3 ;
    wire \pid_alt.un1_pid_prereg_0_cry_3 ;
    wire \pid_alt.un1_pid_prereg_0_cry_4 ;
    wire \pid_alt.un1_pid_prereg_0_cry_5 ;
    wire \pid_alt.un1_pid_prereg_0_cry_6 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIJR3Q5Z0Z_6 ;
    wire bfn_3_16_0_;
    wire \pid_alt.error_d_reg_prev_esr_RNI5G6Q5Z0Z_7 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIUI2T2Z0Z_6 ;
    wire \pid_alt.un1_pid_prereg_0_cry_7 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIN49Q5Z0Z_8 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI7T3T2Z0Z_7 ;
    wire \pid_alt.un1_pid_prereg_0_cry_8 ;
    wire \pid_alt.un1_pid_prereg_0_cry_9 ;
    wire \pid_alt.error_d_reg_prev_esr_RNITPKD4Z0Z_10 ;
    wire \pid_alt.un1_pid_prereg_0_cry_10 ;
    wire \pid_alt.un1_pid_prereg_0_cry_11 ;
    wire \pid_alt.un1_pid_prereg_0_cry_12 ;
    wire \pid_alt.pid_preregZ0Z_14 ;
    wire \pid_alt.un1_pid_prereg_0_cry_13 ;
    wire \pid_alt.un1_pid_prereg_0_cry_14 ;
    wire \pid_alt.pid_preregZ0Z_15 ;
    wire bfn_3_17_0_;
    wire \pid_alt.pid_preregZ0Z_16 ;
    wire \pid_alt.un1_pid_prereg_0_cry_15 ;
    wire \pid_alt.pid_preregZ0Z_17 ;
    wire \pid_alt.un1_pid_prereg_0_cry_16 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIOVN14Z0Z_17 ;
    wire \pid_alt.pid_preregZ0Z_18 ;
    wire \pid_alt.un1_pid_prereg_0_cry_17 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI8IQ14Z0Z_18 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIGKS02Z0Z_17 ;
    wire \pid_alt.pid_preregZ0Z_19 ;
    wire \pid_alt.un1_pid_prereg_0_cry_18 ;
    wire \pid_alt.pid_preregZ0Z_20 ;
    wire \pid_alt.un1_pid_prereg_0_cry_19 ;
    wire \pid_alt.pid_preregZ0Z_21 ;
    wire \pid_alt.un1_pid_prereg_0_cry_20 ;
    wire \pid_alt.pid_preregZ0Z_22 ;
    wire \pid_alt.un1_pid_prereg_0_cry_21 ;
    wire \pid_alt.un1_pid_prereg_0_cry_22 ;
    wire \pid_alt.pid_preregZ0Z_23 ;
    wire bfn_3_18_0_;
    wire \pid_alt.un1_pid_prereg_0_axb_24 ;
    wire \pid_alt.un1_pid_prereg_0_cry_23 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_6_c_RNI3HMQ ;
    wire \pid_alt.error_d_reg_prev_esr_RNICG9B1_0Z0Z_20 ;
    wire \pid_alt.error_p_regZ0Z_19 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIOTT02Z0Z_18 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI86IMZ0Z_19_cascade_ ;
    wire \pid_alt.error_d_reg_prev_esr_RNIK3024Z0Z_19 ;
    wire \pid_alt.un1_pid_prereg_236_1 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI86IMZ0Z_19 ;
    wire \pid_alt.un1_pid_prereg_236_1_cascade_ ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_19_c_RNI4FRJ ;
    wire \pid_alt.error_d_reg_prev_esr_RNIS5212Z0Z_19 ;
    wire \pid_alt.error_d_regZ0Z_19 ;
    wire \pid_alt.error_d_reg_prevZ0Z_19 ;
    wire \pid_alt.error_d_reg_prev_esr_RNICG9B1_1Z0Z_20 ;
    wire \pid_alt.error_d_reg_prev_esr_RNICG9B1Z0Z_20 ;
    wire \pid_alt.error_d_reg_prevZ0Z_20 ;
    wire \pid_alt.error_d_regZ0Z_20 ;
    wire \pid_alt.error_p_regZ0Z_20 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_20_c_RNISVKK ;
    wire \pid_alt.error_d_reg_prev_esr_RNICG9B1_2Z0Z_20 ;
    wire \pid_alt.error_p_regZ0Z_9 ;
    wire \pid_alt.error_d_reg_prevZ0Z_9 ;
    wire \pid_alt.error_d_regZ0Z_9 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIG75T2Z0Z_8 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIL8611Z0Z_9_cascade_ ;
    wire \pid_alt.error_d_reg_prev_esr_RNICI045Z0Z_9 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIL8611Z0Z_9 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIDAHM_0Z0Z_10 ;
    wire \pid_alt.error_d_reg_prev_esr_RNISAR62Z0Z_9 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI8BR02Z0Z_16 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIVSHMZ0Z_16 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI20IM_0Z0Z_17 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIVSHMZ0Z_16_cascade_ ;
    wire \pid_alt.error_i_reg_esr_RNI7ENJZ0Z_17 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI8DL14Z0Z_16 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI02Q02Z0Z_15 ;
    wire \pid_alt.error_p_regZ0Z_16 ;
    wire \pid_alt.error_d_reg_prevZ0Z_16 ;
    wire \pid_alt.error_d_regZ0Z_16 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIVSHM_0Z0Z_16 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIVSHM_0Z0Z_16_cascade_ ;
    wire \pid_alt.error_i_reg_esr_RNI5BMJZ0Z_16 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIOQI14Z0Z_15 ;
    wire \pid_alt.error_i_acumm_esr_RNI33H91Z0Z_4 ;
    wire \pid_alt.error_i_acumm_esr_RNITQE91Z0Z_2 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_15 ;
    wire \pid_alt.error_i_acumm_esr_RNI0VF91Z0Z_3 ;
    wire \pid_alt.un1_reset_0_i_cascade_ ;
    wire \pid_alt.source_pid_1_sqmuxa_0_o2_3_cascade_ ;
    wire \pid_alt.N_51_cascade_ ;
    wire \pid_alt.source_pid_1_sqmuxa_0_a2_0_3 ;
    wire \pid_alt.N_57_cascade_ ;
    wire \pid_alt.un1_reset_1 ;
    wire \pid_alt.source_pid_1_sqmuxa_0_a2_1_7 ;
    wire \pid_alt.N_51 ;
    wire \pid_alt.N_52 ;
    wire \pid_alt.pid_preregZ0Z_4 ;
    wire \pid_alt.N_52_cascade_ ;
    wire \pid_alt.N_54_cascade_ ;
    wire \pid_alt.N_54 ;
    wire \pid_alt.N_72_i_1 ;
    wire \pid_alt.pid_preregZ0Z_2 ;
    wire \pid_alt.pid_preregZ0Z_1 ;
    wire \pid_alt.pid_preregZ0Z_3 ;
    wire \pid_alt.pid_preregZ0Z_0 ;
    wire \pid_alt.source_pid_1_sqmuxa_0_a2_0_2 ;
    wire \Commands_frame_decoder.state_ns_0_a3_0_1Z0Z_2 ;
    wire \Commands_frame_decoder.source_CH4data_1_sqmuxa ;
    wire \pid_alt.pid_preregZ0Z_5 ;
    wire \pid_alt.N_154 ;
    wire \uart_pc.timer_Count_RNIMQ8T1Z0Z_2 ;
    wire \uart_pc.timer_Count_RNILR1B2Z0Z_2 ;
    wire \uart_pc.timer_Count_RNIMQ8T1Z0Z_2_cascade_ ;
    wire \Commands_frame_decoder.source_CH1data8lto7Z0Z_2_cascade_ ;
    wire \Commands_frame_decoder.source_CH1data8_cascade_ ;
    wire \Commands_frame_decoder.source_CH1data8 ;
    wire \Commands_frame_decoder.state_ns_i_a2_0_2_0 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI9S511Z0Z_5_cascade_ ;
    wire \pid_alt.error_d_reg_prev_esr_RNIL81T2Z0Z_5 ;
    wire \pid_alt.error_p_regZ0Z_6 ;
    wire \pid_alt.error_d_reg_prevZ0Z_6 ;
    wire \pid_alt.error_d_regZ0Z_6 ;
    wire \pid_alt.error_d_reg_prev_esr_RNICV511_0Z0Z_6 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI9S511Z0Z_5 ;
    wire \pid_alt.error_d_reg_prev_esr_RNICV511_0Z0Z_6_cascade_ ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_5_c_RNI0DLQ ;
    wire \pid_alt.error_d_reg_prev_esr_RNI171A6Z0Z_5 ;
    wire \pid_alt.error_d_reg_prev_esr_RNICUVC3Z0Z_4 ;
    wire \pid_alt.error_d_regZ0Z_5 ;
    wire \pid_alt.error_d_reg_prevZ0Z_5 ;
    wire \pid_alt.error_p_regZ0Z_5 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI9S511_0Z0Z_5 ;
    wire \pid_alt.error_d_reg_prev_esr_RNICISB3Z0Z_3 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI6P511Z0Z_4 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI9S511_0Z0Z_5_cascade_ ;
    wire \pid_alt.error_d_reg_prev_esr_RNIOGSO6Z0Z_4 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI88G14Z0Z_14 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIPMHMZ0Z_14 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIPMHMZ0Z_14_cascade_ ;
    wire \pid_alt.error_i_reg_esr_RNI38LJZ0Z_15 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIOOO02Z0Z_14 ;
    wire \pid_alt.error_d_reg_prev_esr_RNISPHM_0Z0Z_15 ;
    wire \pid_alt.error_p_regZ0Z_14 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIPMHM_0Z0Z_14_cascade_ ;
    wire \pid_alt.error_d_reg_prev_esr_RNICQF44Z0Z_13 ;
    wire \pid_alt.error_d_regZ0Z_14 ;
    wire \pid_alt.error_d_reg_prevZ0Z_14 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIPMHM_0Z0Z_14 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIMJHMZ0Z_13 ;
    wire \pid_alt.error_i_reg_esr_RNI15KJZ0Z_14 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIGFN02Z0Z_13 ;
    wire \uart_pc.N_126_li_cascade_ ;
    wire \uart_pc.N_143_cascade_ ;
    wire \uart_pc.timer_Count_RNO_0Z0Z_1 ;
    wire \pid_alt.drone_altitude_i_0 ;
    wire bfn_4_18_0_;
    wire \pid_alt.error_axbZ0Z_1 ;
    wire \pid_alt.error_1 ;
    wire \pid_alt.error_cry_0 ;
    wire \pid_alt.error_2 ;
    wire \pid_alt.error_cry_1 ;
    wire \pid_alt.error_3 ;
    wire \pid_alt.error_cry_2 ;
    wire alt_command_0;
    wire \pid_alt.error_4 ;
    wire \pid_alt.error_cry_3 ;
    wire alt_command_1;
    wire \pid_alt.error_5 ;
    wire \pid_alt.error_cry_4 ;
    wire alt_command_2;
    wire \pid_alt.error_6 ;
    wire \pid_alt.error_cry_5 ;
    wire alt_command_3;
    wire \pid_alt.error_7 ;
    wire \pid_alt.error_cry_6 ;
    wire \pid_alt.error_cry_7 ;
    wire \pid_alt.error_8 ;
    wire bfn_4_19_0_;
    wire \pid_alt.error_9 ;
    wire \pid_alt.error_cry_8 ;
    wire \pid_alt.error_10 ;
    wire \pid_alt.error_cry_9 ;
    wire \pid_alt.error_11 ;
    wire \pid_alt.error_cry_10 ;
    wire \pid_alt.error_12 ;
    wire \pid_alt.error_cry_11 ;
    wire \pid_alt.error_13 ;
    wire \pid_alt.error_cry_12 ;
    wire \pid_alt.error_14 ;
    wire \pid_alt.error_cry_13 ;
    wire \pid_alt.error_cry_14 ;
    wire \pid_alt.error_15 ;
    wire \pid_alt.m21_e_0 ;
    wire \pid_alt.error_i_acumm_esr_RNIQMD91Z0Z_1 ;
    wire \pid_alt.error_i_regZ0Z_0 ;
    wire \pid_alt.error_i_reg_esr_RNIT8KA1Z0Z_5 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_7_c_RNI6LNQ ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_9_c_RNIQN3F ;
    wire \pid_alt.m21_e_2_cascade_ ;
    wire \pid_alt.m21_e_8 ;
    wire \pid_alt.m21_e_9 ;
    wire \pid_alt.m21_e_10_cascade_ ;
    wire \pid_alt.N_111_cascade_ ;
    wire \pid_alt.m35_e_3 ;
    wire \pid_alt.m35_e_2 ;
    wire \pid_alt.N_9_0_cascade_ ;
    wire \pid_alt.error_i_acumm_preregZ0Z_1 ;
    wire \pid_alt.N_62_mux_cascade_ ;
    wire \pid_alt.error_i_acummZ0Z_1 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_2 ;
    wire \pid_alt.error_i_acummZ0Z_2 ;
    wire \pid_alt.N_159_cascade_ ;
    wire \pid_alt.error_i_acumm_preregZ0Z_0 ;
    wire \pid_alt.error_i_acummZ0Z_0 ;
    wire \pid_alt.error_i_acummZ0Z_4 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_3 ;
    wire \pid_alt.N_159 ;
    wire \pid_alt.error_i_acumm7lto4 ;
    wire \pid_alt.error_i_acummZ0Z_3 ;
    wire \uart_drone_sync.aux_1__0__0_0 ;
    wire \uart_drone_sync.aux_2__0__0_0 ;
    wire \uart_drone_sync.aux_3__0__0_0 ;
    wire bfn_5_9_0_;
    wire \uart_drone.timer_Count_RNO_0_0_2 ;
    wire \uart_drone.un4_timer_Count_1_cry_1 ;
    wire \uart_drone.un4_timer_Count_1_cry_2 ;
    wire \uart_drone.un4_timer_Count_1_cry_3 ;
    wire \uart_drone.timer_Count_RNO_0_0_4 ;
    wire \pid_alt.pid_preregZ0Z_13 ;
    wire \pid_alt.N_539 ;
    wire \pid_alt.pid_preregZ0Z_24 ;
    wire \pid_alt.pid_preregZ0Z_12 ;
    wire \uart_drone.timer_Count_RNO_0_0_1_cascade_ ;
    wire \uart_drone.timer_CountZ1Z_1 ;
    wire \pid_alt.pid_preregZ0Z_10 ;
    wire \pid_alt.source_pid_1_sqmuxa_0_a2_1_4_cascade_ ;
    wire \pid_alt.source_pid_1_sqmuxa_0_a2_1_5 ;
    wire \pid_alt.pid_preregZ0Z_11 ;
    wire \pid_alt.pid_preregZ0Z_6 ;
    wire \pid_alt.pid_preregZ0Z_7 ;
    wire \pid_alt.pid_preregZ0Z_8 ;
    wire \pid_alt.pid_preregZ0Z_9 ;
    wire \pid_alt.source_pid_9_0_tz_6 ;
    wire \pid_alt.un1_reset_0_i ;
    wire \uart_pc.data_Auxce_0_0_0 ;
    wire \uart_pc.data_AuxZ1Z_0 ;
    wire \uart_pc.data_Auxce_0_1 ;
    wire \uart_pc.data_AuxZ1Z_1 ;
    wire \uart_pc.data_Auxce_0_0_2 ;
    wire \uart_pc.data_AuxZ1Z_2 ;
    wire \uart_pc.data_Auxce_0_3 ;
    wire \uart_pc.data_AuxZ0Z_3 ;
    wire \uart_pc.data_Auxce_0_0_4 ;
    wire \uart_pc.data_AuxZ0Z_4 ;
    wire \uart_pc.data_Auxce_0_5 ;
    wire \uart_pc.data_AuxZ0Z_5 ;
    wire \uart_pc.data_Auxce_0_6 ;
    wire \uart_pc.data_AuxZ0Z_6 ;
    wire \uart_pc.data_AuxZ0Z_7 ;
    wire \uart_pc.N_145_cascade_ ;
    wire \uart_pc.N_144_1 ;
    wire \uart_pc.N_144_1_cascade_ ;
    wire \Commands_frame_decoder.stateZ0Z_12 ;
    wire \Commands_frame_decoder.stateZ0Z_6 ;
    wire alt_kp_4;
    wire \uart_pc.data_rdyc_1 ;
    wire \Commands_frame_decoder.stateZ0Z_2 ;
    wire \Commands_frame_decoder.un1_sink_data_valid_2_0_cascade_ ;
    wire \Commands_frame_decoder.un1_sink_data_valid_2_0 ;
    wire \Commands_frame_decoder.stateZ0Z_3 ;
    wire uart_pc_data_rdy;
    wire \Commands_frame_decoder.source_CH2data_1_sqmuxa ;
    wire \Commands_frame_decoder.source_CH2data_1_sqmuxa_cascade_ ;
    wire \Commands_frame_decoder.stateZ0Z_4 ;
    wire \pid_front.O_0_20 ;
    wire \pid_front.O_0_6 ;
    wire \pid_front.O_0_12 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI64JA4Z0Z_12 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIJGHMZ0Z_12 ;
    wire \pid_alt.error_i_acumm_esr_RNIJ6LMZ0Z_13 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIJGHMZ0Z_12_cascade_ ;
    wire \pid_alt.error_d_reg_prev_esr_RNISAO32Z0Z_12 ;
    wire \pid_alt.error_p_regZ0Z_13 ;
    wire \pid_alt.error_d_reg_prevZ0Z_13 ;
    wire \pid_alt.error_d_regZ0Z_13 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIMJHM_0Z0Z_13 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIAPQ62Z0Z_11 ;
    wire \pid_alt.error_d_reg_prevZ0Z_12 ;
    wire \pid_alt.error_p_regZ0Z_12 ;
    wire \pid_alt.error_d_regZ0Z_12 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIJGHM_0Z0Z_12 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI1FP62Z0Z_10 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIGDHMZ0Z_11 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIJGHM_0Z0Z_12_cascade_ ;
    wire \pid_alt.error_i_reg_esr_RNI7RNPZ0Z_12 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIB8KD4Z0Z_11 ;
    wire drone_altitude_0;
    wire drone_altitude_1;
    wire \dron_frame_decoder_1.drone_altitude_4 ;
    wire drone_altitude_i_4;
    wire \dron_frame_decoder_1.drone_altitude_5 ;
    wire drone_altitude_i_5;
    wire \dron_frame_decoder_1.drone_altitude_6 ;
    wire drone_altitude_i_6;
    wire \dron_frame_decoder_1.drone_altitude_7 ;
    wire drone_altitude_i_7;
    wire drone_altitude_i_8;
    wire drone_altitude_i_9;
    wire alt_kp_0;
    wire alt_kp_1;
    wire alt_kp_2;
    wire alt_kp_3;
    wire alt_kp_5;
    wire alt_kp_6;
    wire alt_kp_7;
    wire \Commands_frame_decoder.state_RNIF38SZ0Z_6 ;
    wire drone_altitude_i_10;
    wire alt_command_4;
    wire alt_command_5;
    wire alt_command_6;
    wire alt_command_7;
    wire \Commands_frame_decoder.un1_sink_data_valid_2_0_0 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_10 ;
    wire \pid_alt.error_i_acummZ0Z_10 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_11 ;
    wire \pid_alt.error_i_acummZ0Z_11 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_6 ;
    wire \pid_alt.error_i_acummZ0Z_6 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_7 ;
    wire \pid_alt.error_i_acummZ0Z_7 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_8 ;
    wire \pid_alt.error_i_acummZ0Z_8 ;
    wire \pid_alt.N_158 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_9 ;
    wire \pid_alt.error_i_acummZ0Z_9 ;
    wire \pid_alt.error_i_acumm7lto12 ;
    wire \pid_alt.N_9_0 ;
    wire \pid_alt.error_i_acummZ0Z_12 ;
    wire \Commands_frame_decoder.N_403 ;
    wire \Commands_frame_decoder.stateZ0Z_10 ;
    wire \reset_module_System.reset6_13 ;
    wire \reset_module_System.reset6_17_cascade_ ;
    wire \reset_module_System.reset6_11 ;
    wire \reset_module_System.reset6_19_cascade_ ;
    wire scaler_4_data_5;
    wire uart_input_pc_c;
    wire \uart_pc_sync.aux_0__0_Z0Z_0 ;
    wire \uart_pc_sync.aux_3__0_Z0Z_0 ;
    wire \uart_pc_sync.aux_1__0_Z0Z_0 ;
    wire \uart_pc_sync.aux_2__0_Z0Z_0 ;
    wire \uart_drone.state_srsts_0_0_0_cascade_ ;
    wire \uart_drone.stateZ0Z_0 ;
    wire \uart_drone.stateZ0Z_1 ;
    wire \uart_drone.state_srsts_i_0_2_cascade_ ;
    wire \uart_drone.timer_CountZ0Z_0 ;
    wire \uart_drone.timer_Count_RNO_0_0_3 ;
    wire \uart_drone.timer_CountZ1Z_2 ;
    wire \uart_drone.N_143 ;
    wire \uart_drone.timer_Count_0_sqmuxa ;
    wire \uart_pc.state_srsts_0_0_0_cascade_ ;
    wire \uart_drone.N_126_li ;
    wire \uart_drone.un1_state_2_0_a3_0 ;
    wire \uart_pc.stateZ0Z_0 ;
    wire \uart_pc.un1_state_7_0 ;
    wire \uart_pc.bit_CountZ0Z_1 ;
    wire \uart_pc.bit_CountZ0Z_2 ;
    wire \uart_pc.state_RNIEAGSZ0Z_4 ;
    wire \Commands_frame_decoder.source_xy_ki_1_sqmuxa ;
    wire \Commands_frame_decoder.source_offset4data_1_sqmuxa ;
    wire \uart_pc.un1_state_4_0_cascade_ ;
    wire \uart_pc.CO0 ;
    wire debug_CH2_18A_c;
    wire \uart_pc.stateZ0Z_1 ;
    wire \uart_pc.state_srsts_i_0_2_cascade_ ;
    wire \uart_pc.stateZ0Z_2 ;
    wire \uart_pc.timer_CountZ1Z_1 ;
    wire bfn_7_15_0_;
    wire \uart_pc.un4_timer_Count_1_cry_1 ;
    wire \uart_pc.un4_timer_Count_1_cry_2 ;
    wire \uart_pc.un4_timer_Count_1_cry_3 ;
    wire \uart_pc.N_126_li ;
    wire \uart_pc.stateZ0Z_4 ;
    wire \uart_pc.un1_state_2_0_a3_0 ;
    wire \uart_pc.un1_state_2_0 ;
    wire \uart_pc.timer_Count_RNO_0Z0Z_3 ;
    wire \uart_pc.timer_CountZ1Z_3 ;
    wire \uart_pc.timer_Count_RNO_0Z0Z_4 ;
    wire \uart_pc.timer_CountZ0Z_4 ;
    wire \uart_pc.timer_Count_RNO_0Z0Z_2 ;
    wire \uart_pc.timer_CountZ1Z_2 ;
    wire \pid_front.N_99_cascade_ ;
    wire \pid_alt.error_axbZ0Z_12 ;
    wire \pid_alt.error_axbZ0Z_13 ;
    wire \pid_alt.error_axbZ0Z_14 ;
    wire \dron_frame_decoder_1.drone_altitude_10 ;
    wire drone_altitude_12;
    wire drone_altitude_13;
    wire drone_altitude_14;
    wire drone_altitude_15;
    wire \dron_frame_decoder_1.drone_altitude_8 ;
    wire \dron_frame_decoder_1.drone_altitude_9 ;
    wire bfn_8_1_0_;
    wire \reset_module_System.countZ0Z_2 ;
    wire \reset_module_System.count_1_2 ;
    wire \reset_module_System.count_1_cry_1 ;
    wire \reset_module_System.countZ0Z_3 ;
    wire \reset_module_System.count_1_cry_2 ;
    wire \reset_module_System.countZ0Z_4 ;
    wire \reset_module_System.count_1_cry_3 ;
    wire \reset_module_System.countZ0Z_5 ;
    wire \reset_module_System.count_1_cry_4 ;
    wire \reset_module_System.countZ0Z_6 ;
    wire \reset_module_System.count_1_cry_5 ;
    wire \reset_module_System.countZ0Z_7 ;
    wire \reset_module_System.count_1_cry_6 ;
    wire \reset_module_System.countZ0Z_8 ;
    wire \reset_module_System.count_1_cry_7 ;
    wire \reset_module_System.count_1_cry_8 ;
    wire \reset_module_System.countZ0Z_9 ;
    wire bfn_8_2_0_;
    wire \reset_module_System.count_1_cry_9 ;
    wire \reset_module_System.count_1_cry_10 ;
    wire \reset_module_System.countZ0Z_12 ;
    wire \reset_module_System.count_1_cry_11 ;
    wire \reset_module_System.count_1_cry_12 ;
    wire \reset_module_System.countZ0Z_14 ;
    wire \reset_module_System.count_1_cry_13 ;
    wire \reset_module_System.count_1_cry_14 ;
    wire \reset_module_System.countZ0Z_16 ;
    wire \reset_module_System.count_1_cry_15 ;
    wire \reset_module_System.count_1_cry_16 ;
    wire \reset_module_System.countZ0Z_17 ;
    wire bfn_8_3_0_;
    wire \reset_module_System.countZ0Z_18 ;
    wire \reset_module_System.count_1_cry_17 ;
    wire \reset_module_System.count_1_cry_18 ;
    wire \reset_module_System.countZ0Z_20 ;
    wire \reset_module_System.count_1_cry_19 ;
    wire \reset_module_System.count_1_cry_20 ;
    wire \reset_module_System.countZ0Z_10 ;
    wire \reset_module_System.countZ0Z_11 ;
    wire \reset_module_System.reset6_3 ;
    wire \reset_module_System.countZ0Z_19 ;
    wire \reset_module_System.countZ0Z_15 ;
    wire \reset_module_System.countZ0Z_21 ;
    wire \reset_module_System.countZ0Z_13 ;
    wire uart_input_drone_c;
    wire \uart_drone_sync.aux_0__0__0_0 ;
    wire \reset_module_System.countZ0Z_0 ;
    wire \reset_module_System.reset6_15 ;
    wire \reset_module_System.reset6_19 ;
    wire \reset_module_System.count_1_1_cascade_ ;
    wire \reset_module_System.reset6_14 ;
    wire \reset_module_System.countZ0Z_1 ;
    wire bfn_8_8_0_;
    wire \ppm_encoder_1.un1_throttle_cry_0 ;
    wire \ppm_encoder_1.un1_throttle_cry_1 ;
    wire throttle_order_3;
    wire \ppm_encoder_1.un1_throttle_cry_2_THRU_CO ;
    wire \ppm_encoder_1.un1_throttle_cry_2 ;
    wire \ppm_encoder_1.un1_throttle_cry_3 ;
    wire throttle_order_5;
    wire \ppm_encoder_1.un1_throttle_cry_4_THRU_CO ;
    wire \ppm_encoder_1.un1_throttle_cry_4 ;
    wire \ppm_encoder_1.un1_throttle_cry_5 ;
    wire \ppm_encoder_1.un1_throttle_cry_6 ;
    wire \ppm_encoder_1.un1_throttle_cry_7 ;
    wire bfn_8_9_0_;
    wire throttle_order_9;
    wire \ppm_encoder_1.un1_throttle_cry_8_THRU_CO ;
    wire \ppm_encoder_1.un1_throttle_cry_8 ;
    wire \ppm_encoder_1.un1_throttle_cry_9 ;
    wire throttle_order_11;
    wire \ppm_encoder_1.un1_throttle_cry_10_THRU_CO ;
    wire \ppm_encoder_1.un1_throttle_cry_10 ;
    wire \ppm_encoder_1.un1_throttle_cry_11 ;
    wire \ppm_encoder_1.un1_throttle_cry_12 ;
    wire \ppm_encoder_1.un1_throttle_cry_13 ;
    wire \ppm_encoder_1.un1_throttle_cry_5_THRU_CO ;
    wire throttle_order_6;
    wire throttle_order_8;
    wire \ppm_encoder_1.un1_throttle_cry_7_THRU_CO ;
    wire debug_CH3_20A_c;
    wire \uart_drone.timer_Count_RNIES9Q1Z0Z_2_cascade_ ;
    wire \uart_pc.N_152 ;
    wire \uart_pc.un1_state_4_0 ;
    wire \uart_pc.stateZ0Z_3 ;
    wire \uart_pc.bit_CountZ0Z_0 ;
    wire \Commands_frame_decoder.source_CH4data_1_sqmuxa_0 ;
    wire \Commands_frame_decoder.source_offset4data_1_sqmuxa_0 ;
    wire \dron_frame_decoder_1.WDTZ0Z_0 ;
    wire bfn_8_13_0_;
    wire \dron_frame_decoder_1.WDTZ0Z_1 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_0 ;
    wire \dron_frame_decoder_1.WDTZ0Z_2 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_1 ;
    wire \dron_frame_decoder_1.WDTZ0Z_3 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_2 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_3 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_4 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_5 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_6 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_7 ;
    wire bfn_8_14_0_;
    wire \dron_frame_decoder_1.un1_WDT_cry_8 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_9 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_10 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_11 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_12 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_13 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_14 ;
    wire \dron_frame_decoder_1.source_data_valid_2_sqmuxa_iZ0 ;
    wire bfn_8_15_0_;
    wire \pid_front.un11lto30_i_a2 ;
    wire \pid_front.un11lto30_i_a2_0 ;
    wire \pid_front.un11lto30_i_a2_1 ;
    wire \pid_front.un11lto30_i_a2_2 ;
    wire \pid_front.un11lto30_i_a2_3 ;
    wire \pid_front.un11lto30_i_a2_4 ;
    wire \pid_front.un11lto30_i_a2_5 ;
    wire \pid_front.un11lto30_i_a2_6 ;
    wire bfn_8_16_0_;
    wire \uart_pc.N_143 ;
    wire \uart_pc.timer_Count_0_sqmuxa ;
    wire \uart_pc.timer_CountZ0Z_0 ;
    wire \pid_front.un11lto30_i_a2_3_and ;
    wire \pid_front.source_pid_1_sqmuxa_1_0_a2_1_4 ;
    wire \pid_front.N_11_i ;
    wire \pid_front.un11lto30_i_a2_0_and ;
    wire \pid_front.un11lto30_i_a2_2_and ;
    wire \pid_front.pid_preregZ0Z_14 ;
    wire \pid_front.un11lto30_i_a2_4_and ;
    wire \pid_front.un11lto30_i_a2_5_and ;
    wire \pid_front.un11lto30_i_a2_4_and_cascade_ ;
    wire \pid_front.source_pid_1_sqmuxa_1_0_a2_0_0 ;
    wire \pid_front.source_pid_1_sqmuxa_1_0_a4_3 ;
    wire \pid_front.N_98_cascade_ ;
    wire \pid_front.un1_pid_prereg_0_9_cascade_ ;
    wire \pid_front.un1_pid_prereg_0_10_cascade_ ;
    wire \pid_front.un1_pid_prereg_0_8 ;
    wire \pid_front.un1_pid_prereg_0_8_cascade_ ;
    wire \pid_front.un1_pid_prereg_0_9 ;
    wire \pid_front.un1_pid_prereg_0_22_cascade_ ;
    wire \pid_front.un1_pid_prereg_0_20 ;
    wire \pid_front.un1_pid_prereg_0_21 ;
    wire \pid_front.un1_pid_prereg_0_20_cascade_ ;
    wire \pid_front.un1_pid_prereg_0_22 ;
    wire \pid_front.un1_pid_prereg_0_25_cascade_ ;
    wire \pid_front.un1_pid_prereg_0_24 ;
    wire \pid_front.un1_pid_prereg_0_26 ;
    wire \pid_front.un1_pid_prereg_0_25 ;
    wire \pid_front.un1_pid_prereg_0_23 ;
    wire \ppm_encoder_1.throttleZ0Z_5 ;
    wire \ppm_encoder_1.elevator_RNIC96OZ0Z_5_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_0_0_5 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_1_5_cascade_ ;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_5_cascade_ ;
    wire \ppm_encoder_1.elevatorZ0Z_5 ;
    wire \ppm_encoder_1.elevator_RNIFC6OZ0Z_8_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_0_2_8_cascade_ ;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_8_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_0_1_8 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_2_3_cascade_ ;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_3_cascade_ ;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_4_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_0_1_4 ;
    wire \ppm_encoder_1.un1_throttle_cry_3_THRU_CO ;
    wire throttle_order_4;
    wire \ppm_encoder_1.throttleZ0Z_4 ;
    wire bfn_9_6_0_;
    wire \ppm_encoder_1.un1_rudder_cry_6 ;
    wire \ppm_encoder_1.un1_rudder_cry_7 ;
    wire \ppm_encoder_1.un1_rudder_cry_8 ;
    wire \ppm_encoder_1.un1_rudder_cry_9 ;
    wire \ppm_encoder_1.un1_rudder_cry_10 ;
    wire \ppm_encoder_1.un1_rudder_cry_11 ;
    wire \ppm_encoder_1.un1_rudder_cry_12 ;
    wire \ppm_encoder_1.un1_rudder_cry_13 ;
    wire bfn_9_7_0_;
    wire \scaler_4.un2_source_data_0_cry_1_c_RNOZ0 ;
    wire bfn_9_8_0_;
    wire scaler_4_data_6;
    wire \scaler_4.un2_source_data_0_cry_1 ;
    wire \scaler_4.un2_source_data_0_cry_2 ;
    wire \scaler_4.un2_source_data_0_cry_3 ;
    wire \scaler_4.un2_source_data_0_cry_4 ;
    wire \scaler_4.un2_source_data_0_cry_5 ;
    wire \scaler_4.un2_source_data_0_cry_6 ;
    wire \scaler_4.un2_source_data_0_cry_7 ;
    wire \scaler_4.un2_source_data_0_cry_8 ;
    wire bfn_9_9_0_;
    wire \scaler_4.un2_source_data_0_cry_9 ;
    wire scaler_4_data_14;
    wire \scaler_4.debug_CH3_20A_c_0 ;
    wire frame_decoder_CH4data_0;
    wire frame_decoder_OFF4data_0;
    wire bfn_9_11_0_;
    wire frame_decoder_CH4data_1;
    wire frame_decoder_OFF4data_1;
    wire \scaler_4.un2_source_data_0 ;
    wire \scaler_4.un3_source_data_0_cry_0 ;
    wire frame_decoder_CH4data_2;
    wire frame_decoder_OFF4data_2;
    wire \scaler_4.un3_source_data_0_cry_1_c_RNI74CL ;
    wire \scaler_4.un3_source_data_0_cry_1 ;
    wire frame_decoder_CH4data_3;
    wire frame_decoder_OFF4data_3;
    wire \scaler_4.un3_source_data_0_cry_2_c_RNIA8DL ;
    wire \scaler_4.un3_source_data_0_cry_2 ;
    wire frame_decoder_CH4data_4;
    wire frame_decoder_OFF4data_4;
    wire \scaler_4.un3_source_data_0_cry_3_c_RNIDCEL ;
    wire \scaler_4.un3_source_data_0_cry_3 ;
    wire frame_decoder_CH4data_5;
    wire frame_decoder_OFF4data_5;
    wire \scaler_4.un3_source_data_0_cry_4_c_RNIGGFL ;
    wire \scaler_4.un3_source_data_0_cry_4 ;
    wire frame_decoder_CH4data_6;
    wire frame_decoder_OFF4data_6;
    wire \scaler_4.un3_source_data_0_cry_5_c_RNIJKGL ;
    wire \scaler_4.un3_source_data_0_cry_5 ;
    wire \scaler_4.un3_source_data_0_axb_7 ;
    wire \scaler_4.un3_source_data_0_cry_6_c_RNIOUNN ;
    wire \scaler_4.un3_source_data_0_cry_6 ;
    wire \scaler_4.un3_source_data_0_cry_7 ;
    wire \scaler_4.un3_source_data_0_cry_7_c_RNIP0PN ;
    wire bfn_9_12_0_;
    wire \scaler_4.un3_source_data_0_cry_8 ;
    wire \scaler_4.un3_source_data_0_cry_8_c_RNIS918 ;
    wire \dron_frame_decoder_1.WDTZ0Z_8 ;
    wire \dron_frame_decoder_1.WDTZ0Z_5 ;
    wire \dron_frame_decoder_1.WDTZ0Z_9 ;
    wire \dron_frame_decoder_1.WDTZ0Z_4 ;
    wire \dron_frame_decoder_1.WDT10_0_i_1_cascade_ ;
    wire \dron_frame_decoder_1.WDT10_0_i ;
    wire \dron_frame_decoder_1.WDTZ0Z_6 ;
    wire \dron_frame_decoder_1.WDTZ0Z_7 ;
    wire \dron_frame_decoder_1.WDTZ0Z_10 ;
    wire \dron_frame_decoder_1.WDT10lto9_3 ;
    wire \dron_frame_decoder_1.WDT10lt12_0 ;
    wire \dron_frame_decoder_1.WDTZ0Z_11 ;
    wire \dron_frame_decoder_1.WDTZ0Z_13 ;
    wire \dron_frame_decoder_1.WDT10lt12_0_cascade_ ;
    wire \dron_frame_decoder_1.WDTZ0Z_12 ;
    wire \dron_frame_decoder_1.WDTZ0Z_14 ;
    wire \dron_frame_decoder_1.WDTZ0Z_15 ;
    wire \dron_frame_decoder_1.WDT10lt14_0_cascade_ ;
    wire \dron_frame_decoder_1.N_218_cascade_ ;
    wire \pid_front.un11lto30_i_a2_6_and ;
    wire \pid_front.source_pid_1_sqmuxa_1_0_o2_sx ;
    wire \pid_front.N_389 ;
    wire \pid_front.N_102_cascade_ ;
    wire \pid_front.un1_reset_0_i_cascade_ ;
    wire \pid_front.N_99 ;
    wire \pid_front.source_pid_1_sqmuxa_1_0_a4_4 ;
    wire \pid_front.source_pid10lt4_0 ;
    wire \pid_front.N_75 ;
    wire bfn_9_17_0_;
    wire \pid_front.pid_preregZ0Z_0 ;
    wire \pid_front.un1_pid_prereg_0_cry_0_c_THRU_CO ;
    wire \pid_front.pid_preregZ0Z_1 ;
    wire \pid_front.un1_pid_prereg_0_cry_0 ;
    wire \pid_front.pid_preregZ0Z_2 ;
    wire \pid_front.un1_pid_prereg_0_cry_1 ;
    wire \pid_front.pid_preregZ0Z_3 ;
    wire \pid_front.un1_pid_prereg_0_cry_2 ;
    wire \pid_front.pid_preregZ0Z_4 ;
    wire \pid_front.un1_pid_prereg_0_cry_3 ;
    wire \pid_front.pid_preregZ0Z_5 ;
    wire \pid_front.un1_pid_prereg_0_cry_4 ;
    wire \pid_front.pid_preregZ0Z_6 ;
    wire \pid_front.un1_pid_prereg_0_cry_5 ;
    wire \pid_front.un1_pid_prereg_0_cry_6 ;
    wire \pid_front.pid_preregZ0Z_7 ;
    wire bfn_9_18_0_;
    wire \pid_front.un1_pid_prereg_0_cry_7 ;
    wire \pid_front.error_p_reg_esr_RNIV7CQ2Z0Z_8 ;
    wire \pid_front.pid_preregZ0Z_9 ;
    wire \pid_front.un1_pid_prereg_0_cry_8 ;
    wire \pid_front.un1_pid_prereg_0_cry_9 ;
    wire \pid_front.un1_pid_prereg_0_cry_10 ;
    wire \pid_front.un1_pid_prereg_0_cry_11 ;
    wire \pid_front.un1_pid_prereg_0_cry_12 ;
    wire \pid_front.un1_pid_prereg_0_cry_13_THRU_CO ;
    wire \pid_front.un1_pid_prereg_0_cry_13 ;
    wire \pid_front.un1_pid_prereg_0_cry_14 ;
    wire \pid_front.pid_preregZ0Z_15 ;
    wire bfn_9_19_0_;
    wire \pid_front.pid_preregZ0Z_16 ;
    wire \pid_front.un1_pid_prereg_0_cry_15 ;
    wire \pid_front.pid_preregZ0Z_17 ;
    wire \pid_front.un1_pid_prereg_0_cry_16 ;
    wire \pid_front.pid_preregZ0Z_18 ;
    wire \pid_front.un1_pid_prereg_0_cry_17 ;
    wire \pid_front.pid_preregZ0Z_19 ;
    wire \pid_front.un1_pid_prereg_0_cry_18 ;
    wire \pid_front.error_p_reg_esr_RNI80EDDZ0Z_17 ;
    wire \pid_front.pid_preregZ0Z_20 ;
    wire \pid_front.un1_pid_prereg_0_cry_19 ;
    wire \pid_front.error_p_reg_esr_RNISOJEDZ0Z_18 ;
    wire \pid_front.error_p_reg_esr_RNIQOPM6Z0Z_18 ;
    wire \pid_front.pid_preregZ0Z_21 ;
    wire \pid_front.un1_pid_prereg_0_cry_20 ;
    wire \pid_front.error_p_reg_esr_RNI20QN6Z0Z_19 ;
    wire \pid_front.pid_preregZ0Z_22 ;
    wire \pid_front.un1_pid_prereg_0_cry_21 ;
    wire \pid_front.un1_pid_prereg_0_cry_22 ;
    wire \pid_front.pid_preregZ0Z_23 ;
    wire bfn_9_20_0_;
    wire \pid_front.pid_preregZ0Z_24 ;
    wire \pid_front.un1_pid_prereg_0_cry_23 ;
    wire \pid_front.pid_preregZ0Z_25 ;
    wire \pid_front.un1_pid_prereg_0_cry_24 ;
    wire \pid_front.error_d_reg_prev_esr_RNIKE2O8Z0Z_22 ;
    wire \pid_front.pid_preregZ0Z_26 ;
    wire \pid_front.un1_pid_prereg_0_cry_25 ;
    wire \pid_front.error_d_reg_prev_esr_RNISQ6O8Z0Z_22 ;
    wire \pid_front.error_d_reg_prev_esr_RNICA2C4Z0Z_22 ;
    wire \pid_front.pid_preregZ0Z_27 ;
    wire \pid_front.un1_pid_prereg_0_cry_26 ;
    wire \pid_front.error_d_reg_prev_esr_RNI36BO8Z0Z_22 ;
    wire \pid_front.error_d_reg_prev_esr_RNIGG4C4Z0Z_22 ;
    wire \pid_front.pid_preregZ0Z_28 ;
    wire \pid_front.un1_pid_prereg_0_cry_27 ;
    wire \pid_front.error_d_reg_prev_esr_RNI7DEO8Z0Z_22 ;
    wire \pid_front.error_d_reg_prev_esr_RNIJL6C4Z0Z_22 ;
    wire \pid_front.pid_preregZ0Z_29 ;
    wire \pid_front.un1_pid_prereg_0_cry_28 ;
    wire \pid_front.un1_pid_prereg_0_axb_30 ;
    wire \pid_front.un1_pid_prereg_0_cry_29 ;
    wire \pid_front.un1_pid_prereg_0_17_cascade_ ;
    wire \pid_front.error_d_reg_prev_esr_RNI4UTB4Z0Z_22 ;
    wire \pid_front.un1_pid_prereg_0_18_cascade_ ;
    wire \pid_front.error_d_reg_prev_esr_RNIC2UN8Z0Z_22 ;
    wire \pid_front.un1_pid_prereg_0_17 ;
    wire \pid_front.error_d_reg_prev_esr_RNIFJ8U9Z0Z_22 ;
    wire \pid_front.un1_pid_prereg_0_19 ;
    wire \pid_front.un1_pid_prereg_0_19_cascade_ ;
    wire \pid_front.un1_pid_prereg_0_18 ;
    wire \pid_front.error_d_reg_prev_esr_RNI840C4Z0Z_22 ;
    wire \pid_front.error_p_reg_esr_RNI1IK9EZ0Z_12 ;
    wire \pid_front.un1_pid_prereg_167_0_1_cascade_ ;
    wire \pid_front.un1_pid_prereg_153_0_cascade_ ;
    wire \pid_front.error_d_reg_prev_esr_RNIHM5CDZ0Z_10 ;
    wire \pid_front.N_2191_i ;
    wire \pid_front.N_2191_i_cascade_ ;
    wire \pid_front.error_p_reg_esr_RNILTVH2Z0Z_12 ;
    wire \pid_front.error_p_reg_esr_RNIJVCREZ0Z_13 ;
    wire \pid_front.error_p_reg_esr_RNIHFPHLZ0Z_13 ;
    wire \pid_front.un1_pid_prereg_0_1_cascade_ ;
    wire \pid_front.error_p_reg_esr_RNIUFCM6Z0Z_14 ;
    wire \pid_front.error_p_reg_esr_RNIH0C61Z0Z_14_cascade_ ;
    wire \pid_front.error_p_reg_esr_RNIH0C61Z0Z_14 ;
    wire \pid_front.error_d_reg_prev_esr_RNI5JRF4Z0Z_10 ;
    wire \pid_front.error_p_reg_esr_RNIK3C61_0Z0Z_15 ;
    wire \pid_front.error_p_regZ0Z_15 ;
    wire \pid_front.error_d_reg_prevZ0Z_15 ;
    wire \pid_front.error_p_regZ0Z_16 ;
    wire \pid_front.error_d_reg_prevZ0Z_16 ;
    wire \pid_front.un1_pid_prereg_0_0 ;
    wire \pid_front.un1_pid_prereg_0_1 ;
    wire \pid_front.error_p_reg_esr_RNICIRCDZ0Z_14 ;
    wire \pid_front.un1_pid_prereg_0_3_cascade_ ;
    wire \pid_front.error_p_reg_esr_RNIE2FM6Z0Z_15 ;
    wire \pid_front.error_p_reg_esr_RNIN6C61Z0Z_16 ;
    wire \pid_front.un1_pid_prereg_0_3 ;
    wire \pid_front.un1_pid_prereg_0_4_cascade_ ;
    wire \pid_front.error_p_reg_esr_RNICN0DDZ0Z_15 ;
    wire \pid_front.un1_pid_prereg_0_5_cascade_ ;
    wire \pid_front.error_p_reg_esr_RNIUKHM6Z0Z_16 ;
    wire \pid_front.error_p_reg_esr_RNIK3C61Z0Z_15 ;
    wire \pid_front.error_p_reg_esr_RNIN6C61_0Z0Z_16 ;
    wire \pid_front.un1_pid_prereg_0_2 ;
    wire scaler_4_data_11;
    wire \ppm_encoder_1.un1_rudder_cry_10_THRU_CO ;
    wire bfn_10_3_0_;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_0 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_1 ;
    wire \ppm_encoder_1.init_pulses_RNIALAI5Z0Z_3 ;
    wire \ppm_encoder_1.N_256_i_i ;
    wire \ppm_encoder_1.un1_init_pulses_10_3 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_2 ;
    wire \ppm_encoder_1.init_pulses_RNIMENT5Z0Z_4 ;
    wire \ppm_encoder_1.N_260_i_i ;
    wire \ppm_encoder_1.un1_init_pulses_10_4 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_3 ;
    wire \ppm_encoder_1.init_pulses_RNISKNT5Z0Z_5 ;
    wire \ppm_encoder_1.N_261_i_i ;
    wire \ppm_encoder_1.un1_init_pulses_10_5 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_4 ;
    wire \ppm_encoder_1.un1_init_pulses_10_6 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_5 ;
    wire \ppm_encoder_1.un1_init_pulses_10_7 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_6 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_7 ;
    wire \ppm_encoder_1.init_pulses_RNI85KU5Z0Z_8 ;
    wire \ppm_encoder_1.N_264_i_i ;
    wire \ppm_encoder_1.un1_init_pulses_10_8 ;
    wire bfn_10_4_0_;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_8 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_9 ;
    wire \ppm_encoder_1.un1_init_pulses_10_11 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_10 ;
    wire \ppm_encoder_1.un1_init_pulses_10_12 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_11 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_12 ;
    wire \ppm_encoder_1.un1_init_pulses_10_14 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_13 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_14 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_15 ;
    wire bfn_10_5_0_;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_16 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_17 ;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_16 ;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_17 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_1_3 ;
    wire \ppm_encoder_1.aileronZ0Z_5 ;
    wire \ppm_encoder_1.un1_rudder_cry_9_THRU_CO ;
    wire scaler_4_data_10;
    wire \ppm_encoder_1.un1_rudder_cry_11_THRU_CO ;
    wire scaler_4_data_12;
    wire \ppm_encoder_1.un1_rudder_cry_6_THRU_CO ;
    wire scaler_4_data_7;
    wire \ppm_encoder_1.un1_rudder_cry_7_THRU_CO ;
    wire scaler_4_data_8;
    wire scaler_4_data_9;
    wire \ppm_encoder_1.un1_rudder_cry_8_THRU_CO ;
    wire \ppm_encoder_1.counter24_0_I_57_c_RNIJMMDZ0_cascade_ ;
    wire ppm_output_c;
    wire \ppm_encoder_1.un1_throttle_cry_9_THRU_CO ;
    wire throttle_order_10;
    wire throttle_order_13;
    wire \ppm_encoder_1.un1_throttle_cry_12_THRU_CO ;
    wire \ppm_encoder_1.un1_throttle_cry_1_THRU_CO ;
    wire throttle_order_2;
    wire \ppm_encoder_1.aileronZ0Z_4 ;
    wire \uart_drone.stateZ0Z_2 ;
    wire \uart_drone.N_145_cascade_ ;
    wire \uart_drone.stateZ0Z_4 ;
    wire \uart_drone.un1_state_4_0_cascade_ ;
    wire \uart_drone.stateZ0Z_3 ;
    wire \uart_drone.N_152_cascade_ ;
    wire bfn_10_11_0_;
    wire front_order_1;
    wire \ppm_encoder_1.un1_elevator_cry_0_THRU_CO ;
    wire \ppm_encoder_1.un1_elevator_cry_0 ;
    wire front_order_2;
    wire \ppm_encoder_1.un1_elevator_cry_1_THRU_CO ;
    wire \ppm_encoder_1.un1_elevator_cry_1 ;
    wire front_order_3;
    wire \ppm_encoder_1.un1_elevator_cry_2_THRU_CO ;
    wire \ppm_encoder_1.un1_elevator_cry_2 ;
    wire front_order_4;
    wire \ppm_encoder_1.un1_elevator_cry_3_THRU_CO ;
    wire \ppm_encoder_1.un1_elevator_cry_3 ;
    wire front_order_5;
    wire \ppm_encoder_1.un1_elevator_cry_4_THRU_CO ;
    wire \ppm_encoder_1.un1_elevator_cry_4 ;
    wire \ppm_encoder_1.un1_elevator_cry_5 ;
    wire \ppm_encoder_1.un1_elevator_cry_6 ;
    wire \ppm_encoder_1.un1_elevator_cry_7 ;
    wire \ppm_encoder_1.un1_elevator_cry_7_THRU_CO ;
    wire bfn_10_12_0_;
    wire front_order_9;
    wire \ppm_encoder_1.un1_elevator_cry_8_THRU_CO ;
    wire \ppm_encoder_1.un1_elevator_cry_8 ;
    wire \ppm_encoder_1.un1_elevator_cry_9_THRU_CO ;
    wire \ppm_encoder_1.un1_elevator_cry_9 ;
    wire \ppm_encoder_1.un1_elevator_cry_10_THRU_CO ;
    wire \ppm_encoder_1.un1_elevator_cry_10 ;
    wire \ppm_encoder_1.un1_elevator_cry_11_THRU_CO ;
    wire \ppm_encoder_1.un1_elevator_cry_11 ;
    wire \ppm_encoder_1.un1_elevator_cry_12_THRU_CO ;
    wire \ppm_encoder_1.un1_elevator_cry_12 ;
    wire \ppm_encoder_1.un1_elevator_cry_13 ;
    wire front_order_13;
    wire \pid_front.N_98 ;
    wire \pid_front.pid_preregZ0Z_13 ;
    wire \pid_front.pid_preregZ0Z_12 ;
    wire front_order_12;
    wire \pid_front.pid_preregZ0Z_8 ;
    wire front_order_8;
    wire \pid_front.pid_preregZ0Z_11 ;
    wire front_order_11;
    wire \pid_front.N_76 ;
    wire \pid_front.pid_preregZ0Z_30 ;
    wire \pid_front.pid_preregZ0Z_10 ;
    wire front_order_10;
    wire \pid_front.state_0_1 ;
    wire \pid_front.un1_reset_0_i ;
    wire \pid_front.error_p_reg_esr_RNID8VU1Z0Z_3 ;
    wire \pid_front.error_p_reg_esr_RNIUAE8_0Z0Z_4 ;
    wire \pid_front.error_p_reg_esr_RNIUAE8_0Z0Z_4_cascade_ ;
    wire \pid_front.error_p_reg_esr_RNIMI772Z0Z_3 ;
    wire \pid_front.error_p_reg_esr_RNIB9N71_0Z0Z_5 ;
    wire \pid_front.error_p_regZ0Z_4 ;
    wire \pid_front.error_d_reg_prevZ0Z_4 ;
    wire \pid_front.error_p_reg_esr_RNIUAE8Z0Z_4_cascade_ ;
    wire \pid_front.error_p_reg_esr_RNIVOSG_0Z0Z_5_cascade_ ;
    wire \pid_front.error_p_reg_esr_RNIB9N71Z0Z_5 ;
    wire \pid_front.error_p_reg_esr_RNI6B6F_0Z0Z_6_cascade_ ;
    wire \pid_front.error_p_reg_esr_RNIVOSG_0Z0Z_5 ;
    wire \pid_front.un1_pid_prereg_66_0_cascade_ ;
    wire \pid_front.error_p_reg_esr_RNI8CGM2Z0Z_5 ;
    wire \pid_front.error_p_reg_esr_RNI6B6F_0Z0Z_6 ;
    wire \pid_front.error_p_reg_esr_RNIT2PE1Z0Z_5 ;
    wire \pid_front.error_p_regZ0Z_5 ;
    wire \pid_front.error_p_reg_esr_RNIUAE8Z0Z_4 ;
    wire \pid_front.error_p_reg_esr_RNIVOSGZ0Z_5 ;
    wire \pid_front.N_2155_i ;
    wire \pid_front.N_2155_i_cascade_ ;
    wire \pid_front.error_p_regZ0Z_6 ;
    wire \pid_front.N_2179_i_cascade_ ;
    wire \pid_front.error_p_reg_esr_RNIFM3D1Z0Z_10_cascade_ ;
    wire \pid_front.error_p_reg_esr_RNIS5CU3Z0Z_9 ;
    wire \pid_front.error_p_reg_esr_RNILQ6FZ0Z_9 ;
    wire \pid_front.error_p_reg_esr_RNIFM3D1Z0Z_10 ;
    wire \pid_front.error_p_reg_esr_RNILQ6FZ0Z_9_cascade_ ;
    wire \pid_front.error_p_reg_esr_RNIEB5T7Z0Z_9 ;
    wire \pid_front.error_p_regZ0Z_9 ;
    wire \pid_front.error_p_reg_esr_RNILQ6F_0Z0Z_9 ;
    wire \pid_front.error_p_reg_esr_RNILQ6F_0Z0Z_9_cascade_ ;
    wire \pid_front.error_p_reg_esr_RNI6R6D1Z0Z_8 ;
    wire \pid_front.un1_pid_prereg_0_15_cascade_ ;
    wire \pid_front.error_d_reg_prev_esr_RNIBLAI5Z0Z_22 ;
    wire \pid_front.un1_pid_prereg_0_10 ;
    wire \pid_front.un1_pid_prereg_0_11 ;
    wire \pid_front.error_p_reg_esr_RNIF7HGDZ0Z_19 ;
    wire \pid_front.un1_pid_prereg_0_14 ;
    wire \pid_front.un1_pid_prereg_0_14_cascade_ ;
    wire \pid_front.un1_pid_prereg_0_15 ;
    wire \pid_front.error_d_reg_prev_esr_RNIOS1BCZ0Z_22 ;
    wire \pid_front.un1_pid_prereg_370_1 ;
    wire \pid_front.un1_pid_prereg_370_1_cascade_ ;
    wire \pid_front.un1_pid_prereg_0_13 ;
    wire \pid_front.un1_pid_prereg_0_13_cascade_ ;
    wire \pid_front.error_p_reg_esr_RNID7NO6Z0Z_20 ;
    wire \pid_front.g1_1_cascade_ ;
    wire \pid_front.g0_3_2_cascade_ ;
    wire \pid_front.g0_1_0_1 ;
    wire \pid_front.N_4_1_1_1 ;
    wire \pid_front.g0_1_cascade_ ;
    wire \pid_front.g0_2_0 ;
    wire \pid_front.error_p_reg_esr_RNIU52U6Z0Z_12_cascade_ ;
    wire \pid_front.g1_3 ;
    wire \pid_front.g1_2_1 ;
    wire \pid_front.error_p_reg_esr_RNICU3D1_0Z0Z_6 ;
    wire \pid_front.error_p_reg_esr_RNI6B6FZ0Z_6 ;
    wire \pid_front.N_2198_0_0_0 ;
    wire \pid_front.error_d_reg_fast_esr_RNID6KB1Z0Z_12_cascade_ ;
    wire \pid_front.error_d_reg_fast_esr_RNIQSG63Z0Z_12_cascade_ ;
    wire \pid_front.error_p_reg_esr_RNIETB61_1Z0Z_13 ;
    wire \pid_front.un1_pid_prereg_97_cascade_ ;
    wire \pid_front.un1_pid_prereg_167_0 ;
    wire \pid_front.error_p_reg_esr_RNI8C7GBZ0Z_13 ;
    wire \pid_front.error_p_reg_esr_RNIT79QCZ0Z_12 ;
    wire \pid_front.error_p_reg_esr_RNI8C7GBZ0Z_13_cascade_ ;
    wire \pid_front.error_p_reg_esr_RNIBJ5B3_0Z0Z_14 ;
    wire \pid_front.error_p_reg_esr_RNIG7MLRZ0Z_12 ;
    wire \pid_front.error_d_reg_fast_esr_RNI5VGKZ0Z_12 ;
    wire \pid_front.error_d_reg_prevZ0Z_22 ;
    wire \pid_front.un1_pid_prereg_0_16 ;
    wire \pid_front.O_12 ;
    wire \pid_front.O_13 ;
    wire \pid_front.O_11 ;
    wire \pid_front.error_d_reg_fastZ0Z_12 ;
    wire \pid_front.O_15 ;
    wire \pid_front.error_p_reg_esr_RNIKG5U_0Z0Z_10_cascade_ ;
    wire \pid_front.error_p_reg_esr_RNIKG5UZ0Z_10 ;
    wire \pid_front.error_d_reg_prev_esr_RNI379B2Z0Z_10 ;
    wire \pid_front.error_d_reg_prevZ0Z_10 ;
    wire \pid_front.error_d_regZ0Z_10 ;
    wire \pid_front.error_d_reg_prev_esr_RNI379B2Z0Z_10_cascade_ ;
    wire \pid_front.error_p_reg_esr_RNI8NB61_1Z0Z_11 ;
    wire \pid_front.error_d_reg_prev_esr_RNI5JRF4_0Z0Z_10_cascade_ ;
    wire \pid_front.error_d_reg_prev_esr_RNIO00C5_0Z0Z_10 ;
    wire \pid_front.error_d_reg_prev_esr_RNI5JRF4_0Z0Z_10 ;
    wire \pid_front.error_d_reg_prev_esr_RNIO00C5Z0Z_10 ;
    wire \pid_front.error_d_regZ0Z_9 ;
    wire \pid_front.error_d_reg_prevZ0Z_9 ;
    wire \pid_front.N_2173_i ;
    wire \pid_front.state_RNIPKTDZ0Z_0 ;
    wire \ppm_encoder_1.N_39_i ;
    wire bfn_11_1_0_;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_0 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_1 ;
    wire \ppm_encoder_1.un1_init_pulses_11_3 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_2 ;
    wire \ppm_encoder_1.un1_init_pulses_11_4 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_3 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_5 ;
    wire \ppm_encoder_1.un1_init_pulses_11_5 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_4 ;
    wire \ppm_encoder_1.un1_init_pulses_11_6 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_5 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_7 ;
    wire \ppm_encoder_1.un1_init_pulses_11_7 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_6 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_7 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_8 ;
    wire \ppm_encoder_1.un1_init_pulses_11_8 ;
    wire bfn_11_2_0_;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_8 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_9 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_11 ;
    wire \ppm_encoder_1.un1_init_pulses_11_11 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_10 ;
    wire \ppm_encoder_1.un1_init_pulses_11_12 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_11 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_12 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_14 ;
    wire \ppm_encoder_1.un1_init_pulses_11_14 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_13 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_14 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_15 ;
    wire bfn_11_3_0_;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_16 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_17 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_15 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_16 ;
    wire \ppm_encoder_1.un1_init_pulses_11_15 ;
    wire \ppm_encoder_1.un1_init_pulses_10_15 ;
    wire \ppm_encoder_1.un1_init_pulses_10_16 ;
    wire \ppm_encoder_1.un1_init_pulses_11_16 ;
    wire \ppm_encoder_1.un1_init_pulses_11_17 ;
    wire \ppm_encoder_1.un1_init_pulses_10_17 ;
    wire \ppm_encoder_1.un1_init_pulses_11_18 ;
    wire \ppm_encoder_1.un1_init_pulses_10_18 ;
    wire \ppm_encoder_1.un1_init_pulses_10_1 ;
    wire \ppm_encoder_1.un1_init_pulses_11_1 ;
    wire \ppm_encoder_1.un1_init_pulses_10_10 ;
    wire \ppm_encoder_1.un1_init_pulses_11_10 ;
    wire \ppm_encoder_1.un1_init_pulses_11_9 ;
    wire \ppm_encoder_1.un1_init_pulses_10_9 ;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_9_cascade_ ;
    wire \ppm_encoder_1.init_pulses_RNIEBKU5Z0Z_9 ;
    wire \ppm_encoder_1.N_265_i_i ;
    wire \ppm_encoder_1.throttleZ0Z_9 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_1_9 ;
    wire \ppm_encoder_1.elevatorZ0Z_4 ;
    wire \ppm_encoder_1.rudder_RNIM1KQZ0Z_12_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_0_2_12_cascade_ ;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_12_cascade_ ;
    wire \ppm_encoder_1.N_267_i_i ;
    wire \ppm_encoder_1.init_pulses_RNI7OHF5Z0Z_12 ;
    wire \ppm_encoder_1.elevatorZ0Z_12 ;
    wire throttle_order_12;
    wire \ppm_encoder_1.un1_throttle_cry_11_THRU_CO ;
    wire \ppm_encoder_1.throttleZ0Z_12 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_1_12 ;
    wire \ppm_encoder_1.un1_throttle_cry_6_THRU_CO ;
    wire throttle_order_7;
    wire \ppm_encoder_1.elevatorZ0Z_8 ;
    wire \ppm_encoder_1.aileronZ0Z_8 ;
    wire \ppm_encoder_1.aileronZ0Z_9 ;
    wire \ppm_encoder_1.elevatorZ0Z_9 ;
    wire bfn_11_9_0_;
    wire \ppm_encoder_1.un1_aileron_cry_0 ;
    wire \ppm_encoder_1.un1_aileron_cry_1_THRU_CO ;
    wire \ppm_encoder_1.un1_aileron_cry_1 ;
    wire \ppm_encoder_1.un1_aileron_cry_2 ;
    wire \ppm_encoder_1.un1_aileron_cry_3_THRU_CO ;
    wire \ppm_encoder_1.un1_aileron_cry_3 ;
    wire \ppm_encoder_1.un1_aileron_cry_4_THRU_CO ;
    wire \ppm_encoder_1.un1_aileron_cry_4 ;
    wire \ppm_encoder_1.un1_aileron_cry_5 ;
    wire \ppm_encoder_1.un1_aileron_cry_6 ;
    wire \ppm_encoder_1.un1_aileron_cry_7 ;
    wire \ppm_encoder_1.un1_aileron_cry_7_THRU_CO ;
    wire bfn_11_10_0_;
    wire \ppm_encoder_1.un1_aileron_cry_8_THRU_CO ;
    wire \ppm_encoder_1.un1_aileron_cry_8 ;
    wire \ppm_encoder_1.un1_aileron_cry_9_THRU_CO ;
    wire \ppm_encoder_1.un1_aileron_cry_9 ;
    wire \ppm_encoder_1.un1_aileron_cry_10_THRU_CO ;
    wire \ppm_encoder_1.un1_aileron_cry_10 ;
    wire \ppm_encoder_1.un1_aileron_cry_11 ;
    wire \ppm_encoder_1.un1_aileron_cry_12_THRU_CO ;
    wire \ppm_encoder_1.un1_aileron_cry_12 ;
    wire \ppm_encoder_1.un1_aileron_cry_13 ;
    wire \uart_drone.data_Auxce_0_3 ;
    wire \uart_drone.un1_state_2_0 ;
    wire \uart_drone.state_RNIOU0NZ0Z_4 ;
    wire \uart_drone.data_AuxZ0Z_0 ;
    wire \uart_drone.data_AuxZ0Z_1 ;
    wire \uart_drone.data_AuxZ0Z_2 ;
    wire \uart_drone.data_AuxZ0Z_3 ;
    wire \uart_drone.data_AuxZ0Z_4 ;
    wire \uart_drone.data_AuxZ0Z_5 ;
    wire \uart_drone.data_AuxZ0Z_6 ;
    wire \uart_drone.data_AuxZ0Z_7 ;
    wire \uart_drone.data_rdyc_1_0 ;
    wire \uart_drone.timer_Count_RNIES9Q1Z0Z_2 ;
    wire \dron_frame_decoder_1.N_230_5_cascade_ ;
    wire \dron_frame_decoder_1.N_224_cascade_ ;
    wire \dron_frame_decoder_1.state_ns_i_a2_1_1Z0Z_0_cascade_ ;
    wire \dron_frame_decoder_1.N_220 ;
    wire \dron_frame_decoder_1.N_224 ;
    wire \dron_frame_decoder_1.N_220_cascade_ ;
    wire \dron_frame_decoder_1.N_198 ;
    wire \dron_frame_decoder_1.state_ns_i_a2_0_2_0 ;
    wire \dron_frame_decoder_1.un1_sink_data_valid_5_i_0 ;
    wire \dron_frame_decoder_1.un1_sink_data_valid_5_i_0_cascade_ ;
    wire \dron_frame_decoder_1.state_RNI3T3K1Z0Z_7_cascade_ ;
    wire \dron_frame_decoder_1.N_732_0 ;
    wire debug_CH0_16A_c;
    wire \uart_drone.data_rdyc_1 ;
    wire \dron_frame_decoder_1.stateZ0Z_5 ;
    wire \dron_frame_decoder_1.stateZ0Z_4 ;
    wire \dron_frame_decoder_1.state_RNI6P6KZ0Z_4_cascade_ ;
    wire \pid_front.N_2167_i_cascade_ ;
    wire \dron_frame_decoder_1.stateZ0Z_2 ;
    wire \pid_front.error_p_reg_esr_RNIPC5D1Z0Z_7 ;
    wire \pid_front.error_p_reg_esr_RNIBG6FZ0Z_7 ;
    wire \pid_front.error_p_reg_esr_RNIGL6F_0Z0Z_8 ;
    wire \pid_front.error_p_reg_esr_RNICU3D1Z0Z_6 ;
    wire \pid_front.error_p_reg_esr_RNIBG6FZ0Z_7_cascade_ ;
    wire \pid_front.error_p_reg_esr_RNI5B9Q2Z0Z_7 ;
    wire \pid_front.N_2161_i ;
    wire \pid_front.error_p_regZ0Z_7 ;
    wire \pid_front.error_d_reg_prevZ0Z_6 ;
    wire \pid_front.N_2161_i_cascade_ ;
    wire \pid_front.error_p_reg_esr_RNIBG6F_0Z0Z_7 ;
    wire \pid_front.error_p_regZ0Z_8 ;
    wire \pid_front.error_d_reg_prevZ0Z_7 ;
    wire \pid_front.N_2167_i ;
    wire \pid_front.error_p_reg_esr_RNIGL6FZ0Z_8 ;
    wire \dron_frame_decoder_1.drone_H_disp_side_10 ;
    wire \dron_frame_decoder_1.drone_H_disp_side_8 ;
    wire \dron_frame_decoder_1.drone_H_disp_side_9 ;
    wire \dron_frame_decoder_1.N_716_0 ;
    wire \pid_alt.error_i_acumm7lto5 ;
    wire \pid_alt.N_62_mux ;
    wire \pid_alt.error_i_acummZ0Z_5 ;
    wire \pid_front.error_d_reg_prev_esr_RNIBTE61_0Z0Z_21 ;
    wire \pid_front.error_d_reg_prev_esr_RNIBTE61_0Z0Z_21_cascade_ ;
    wire \pid_front.un1_pid_prereg_0_12 ;
    wire \pid_front.error_p_reg_esr_RNI8QE61Z0Z_20 ;
    wire \pid_front.error_p_regZ0Z_21 ;
    wire \pid_front.error_d_reg_prev_esr_RNIBTE61Z0Z_21 ;
    wire \pid_front.error_p_regZ0Z_20 ;
    wire \pid_front.error_p_reg_esr_RNI8QE61_0Z0Z_20 ;
    wire \pid_front.error_d_reg_fast_esr_RNIQSG63Z0Z_12 ;
    wire \pid_front.N_5 ;
    wire \pid_front.error_d_reg_prevZ0Z_20 ;
    wire \pid_front.error_d_reg_prevZ0Z_21 ;
    wire \pid_front.error_d_reg_prevZ0Z_5 ;
    wire \pid_front.error_d_reg_prevZ0Z_8 ;
    wire \pid_front.error_d_reg_prev_fastZ0Z_12 ;
    wire \pid_front.error_p_regZ0Z_12 ;
    wire \pid_front.N_3_i_1_1_cascade_ ;
    wire \pid_front.un1_pid_prereg_79 ;
    wire \pid_front.error_p_regZ0Z_13 ;
    wire \pid_front.error_d_reg_prevZ0Z_13 ;
    wire \pid_front.error_d_regZ0Z_13 ;
    wire \pid_front.N_2198_0_cascade_ ;
    wire \pid_front.N_5_0 ;
    wire \pid_front.N_5_0_0 ;
    wire \pid_front.g0_2_cascade_ ;
    wire \pid_front.N_3_i_1 ;
    wire \pid_front.error_p_reg_esr_RNI6D5L7Z0Z_12_cascade_ ;
    wire \pid_front.error_d_reg_prev_esr_RNI6J3B5Z0Z_12 ;
    wire \pid_front.un1_pid_prereg_0_axb_14 ;
    wire \pid_front.error_d_reg_prevZ0Z_12 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_21 ;
    wire \pid_alt.error_i_acumm7lto13 ;
    wire \pid_alt.N_545 ;
    wire \pid_alt.error_i_acummZ0Z_13 ;
    wire \pid_alt.N_72_i_0 ;
    wire \pid_alt.un1_reset_1_0_i ;
    wire \pid_front.error_d_reg_prevZ0Z_19 ;
    wire \pid_front.error_p_regZ0Z_19 ;
    wire \pid_front.error_p_reg_esr_RNI0GC61Z0Z_19 ;
    wire \pid_front.un1_pid_prereg_135_0 ;
    wire \pid_front.error_d_reg_prevZ0Z_11 ;
    wire \pid_front.error_d_regZ0Z_11 ;
    wire \pid_front.error_p_regZ0Z_11 ;
    wire \pid_front.g0_1_0 ;
    wire \pid_front.O_6 ;
    wire \pid_front.error_d_regZ0Z_4 ;
    wire \pid_front.O_7 ;
    wire \pid_front.error_d_regZ0Z_5 ;
    wire \pid_front.O_8 ;
    wire \pid_front.error_d_regZ0Z_6 ;
    wire \pid_front.O_9 ;
    wire \pid_front.error_d_regZ0Z_7 ;
    wire \pid_front.O_10 ;
    wire \pid_front.error_d_regZ0Z_8 ;
    wire \pid_front.O_14 ;
    wire \pid_front.error_d_regZ0Z_12 ;
    wire \pid_front.O_0_3 ;
    wire \pid_front.error_p_regZ0Z_0 ;
    wire \pid_front.O_0_13 ;
    wire \pid_front.error_p_regZ0Z_10 ;
    wire \pid_front.un10lt9_1_cascade_ ;
    wire \pid_front.un10lt9_cascade_ ;
    wire \pid_front.un10lt9_1 ;
    wire \pid_front.error_i_acumm16lt9_0_cascade_ ;
    wire \pid_front.error_i_acumm_prereg_esr_RNISDO3Z0Z_7 ;
    wire \pid_front.O_0_4 ;
    wire \pid_front.un1_pid_prereg_9_0_cascade_ ;
    wire \pid_front.error_d_reg_prev_esr_RNIMRLTZ0Z_0 ;
    wire \pid_front.O_3 ;
    wire \pid_front.error_d_reg_prev_esr_RNIAHDKZ0Z_0 ;
    wire \pid_front.error_i_acumm_prereg_esr_RNIRU7IZ0Z_10_cascade_ ;
    wire \pid_front.un10lt11_0 ;
    wire \pid_front.O_2 ;
    wire \pid_front.un10lto27_9_cascade_ ;
    wire \pid_front.error_i_acumm_prereg_esr_RNI18694_0Z0Z_14 ;
    wire \pid_front.un10lto27_10 ;
    wire \pid_front.error_i_acumm_preregZ0Z_19 ;
    wire \pid_front.error_i_acumm_preregZ0Z_18 ;
    wire \pid_front.error_i_acumm_preregZ0Z_14 ;
    wire \pid_front.error_i_acumm_preregZ0Z_15 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_1 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_3 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_10 ;
    wire \ppm_encoder_1.elevatorZ0Z_14 ;
    wire \ppm_encoder_1.rudderZ0Z_14 ;
    wire \ppm_encoder_1.N_56_cascade_ ;
    wire \ppm_encoder_1.init_pulses_RNIV9203Z0Z_6 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_12 ;
    wire \ppm_encoder_1.N_254_i_i ;
    wire \ppm_encoder_1.N_254_i_i_cascade_ ;
    wire \ppm_encoder_1.init_pulses_RNI82G01Z0Z_15 ;
    wire \ppm_encoder_1.N_268_i_i_cascade_ ;
    wire \ppm_encoder_1.init_pulses_RNITIRP2Z0Z_13 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_0_6 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_1_6_cascade_ ;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_6_cascade_ ;
    wire \ppm_encoder_1.N_262_i_i ;
    wire \ppm_encoder_1.init_pulses_RNIPOJU5Z0Z_6 ;
    wire \ppm_encoder_1.elevator_RNIB86OZ0Z_4 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_2_4 ;
    wire scaler_4_data_4;
    wire \ppm_encoder_1.pid_altitude_dv_0 ;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_10_cascade_ ;
    wire \ppm_encoder_1.init_pulses_RNIUCPF5Z0Z_10 ;
    wire \ppm_encoder_1.elevator_RNIGD6OZ0Z_9 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_2_9 ;
    wire \ppm_encoder_1.elevator_RNIOEGEZ0Z_10 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_2_10 ;
    wire \ppm_encoder_1.N_255_i_i ;
    wire \ppm_encoder_1.un1_aileron_cry_0_THRU_CO ;
    wire \ppm_encoder_1.un1_throttle_cry_0_THRU_CO ;
    wire throttle_order_1;
    wire \ppm_encoder_1.un1_elevator_cry_6_THRU_CO ;
    wire front_order_7;
    wire \ppm_encoder_1.elevatorZ0Z_7 ;
    wire \ppm_encoder_1.pulses2count_9_0_3_1_11_cascade_ ;
    wire \ppm_encoder_1.elevatorZ0Z_13 ;
    wire \ppm_encoder_1.rudderZ0Z_12 ;
    wire \ppm_encoder_1.pulses2count_9_0_3_1_12 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_12_cascade_ ;
    wire \ppm_encoder_1.init_pulsesZ0Z_12 ;
    wire \uart_drone.data_Auxce_0_1 ;
    wire \uart_drone.data_Auxce_0_0_2 ;
    wire \uart_drone.data_Auxce_0_0_4 ;
    wire \uart_drone.data_Auxce_0_5 ;
    wire \uart_drone.data_Auxce_0_6 ;
    wire \ppm_encoder_1.un1_aileron_cry_2_THRU_CO ;
    wire \ppm_encoder_1.un1_aileron_cry_11_THRU_CO ;
    wire \ppm_encoder_1.un1_elevator_cry_5_THRU_CO ;
    wire front_order_6;
    wire \ppm_encoder_1.elevatorZ0Z_6 ;
    wire \ppm_encoder_1.un1_aileron_cry_5_THRU_CO ;
    wire \ppm_encoder_1.un1_aileron_cry_6_THRU_CO ;
    wire \uart_drone.un1_state_4_0 ;
    wire \uart_drone.CO0 ;
    wire \uart_drone.un1_state_7_0 ;
    wire \uart_drone.N_152 ;
    wire \uart_drone.timer_CountZ1Z_3 ;
    wire \uart_drone.timer_CountZ0Z_4 ;
    wire \uart_drone.N_144_1 ;
    wire xy_kp_5;
    wire xy_kp_6;
    wire \pid_side.state_RNIL5IFZ0Z_0 ;
    wire \dron_frame_decoder_1.state_ns_0_i_a2_0_2_3_cascade_ ;
    wire \dron_frame_decoder_1.stateZ0Z_3 ;
    wire \dron_frame_decoder_1.N_230_5 ;
    wire \dron_frame_decoder_1.state_ns_0_i_a2_0_3_3 ;
    wire \dron_frame_decoder_1.stateZ0Z_1 ;
    wire \dron_frame_decoder_1.N_200 ;
    wire \dron_frame_decoder_1.stateZ0Z_0 ;
    wire \dron_frame_decoder_1.state_ns_i_a2_0_1_0 ;
    wire \dron_frame_decoder_1.stateZ0Z_6 ;
    wire uart_drone_data_rdy;
    wire \Commands_frame_decoder.source_CH3data_1_sqmuxa ;
    wire xy_kp_0;
    wire xy_kp_2;
    wire xy_kp_3;
    wire xy_kp_7;
    wire \dron_frame_decoder_1.state_RNI4N6KZ0Z_2 ;
    wire \dron_frame_decoder_1.N_218 ;
    wire \dron_frame_decoder_1.state_RNI6P6KZ0Z_4 ;
    wire \dron_frame_decoder_1.stateZ0Z_7 ;
    wire \pid_front.error_i_acumm_prereg_esr_RNIRU7I_0Z0Z_10 ;
    wire \pid_front.state_RNIM14NZ0Z_0 ;
    wire \pid_front.state_RNIVIRQZ0Z_0 ;
    wire \pid_front.error_p_reg_esr_RNI3I672Z0Z_2 ;
    wire \pid_front.error_p_reg_esr_RNIO4E8Z0Z_2 ;
    wire \pid_front.error_p_reg_esr_RNIO4E8Z0Z_2_cascade_ ;
    wire \pid_front.error_p_reg_esr_RNI2VEVZ0Z_2 ;
    wire \pid_front.error_p_reg_esr_RNIR7E8_0Z0Z_3 ;
    wire \pid_front.error_p_regZ0Z_2 ;
    wire \pid_front.error_d_reg_prevZ0Z_2 ;
    wire \pid_front.error_p_regZ0Z_3 ;
    wire \pid_front.error_d_reg_prevZ0Z_3 ;
    wire \pid_front.error_p_reg_esr_RNIR7E8Z0Z_3 ;
    wire \pid_alt.error_p_regZ0Z_15 ;
    wire \pid_alt.error_d_reg_prev_esr_RNISPHMZ0Z_15 ;
    wire \pid_alt.error_d_regZ0Z_15 ;
    wire \pid_alt.error_d_reg_prevZ0Z_15 ;
    wire \pid_alt.state_0_g_0 ;
    wire \pid_front.error_p_reg_esr_RNIETB61_4Z0Z_13 ;
    wire \pid_front.error_d_reg_prev_esr_RNIOLN44Z0Z_12 ;
    wire \pid_front.error_d_reg_prev_esr_RNI8SE96Z0Z_12 ;
    wire \pid_front.error_p_reg_esr_RNIQ9C61Z0Z_17 ;
    wire \pid_front.error_p_reg_esr_RNIQ9C61Z0Z_17_cascade_ ;
    wire \pid_front.error_p_reg_esr_RNITCC61_0Z0Z_18 ;
    wire \pid_front.un1_pid_prereg_0_4 ;
    wire \pid_front.un1_pid_prereg_0_5 ;
    wire \pid_front.un1_pid_prereg_0_6_cascade_ ;
    wire \pid_front.error_p_reg_esr_RNICS5DDZ0Z_16 ;
    wire \pid_front.error_p_regZ0Z_17 ;
    wire \pid_front.error_d_reg_prevZ0Z_17 ;
    wire \pid_front.error_p_reg_esr_RNIQ9C61_0Z0Z_17 ;
    wire \pid_front.error_p_reg_esr_RNI0GC61_0Z0Z_19 ;
    wire \pid_front.un1_pid_prereg_0_7 ;
    wire \pid_front.un1_pid_prereg_0_7_cascade_ ;
    wire \pid_front.un1_pid_prereg_0_6 ;
    wire \pid_front.error_p_reg_esr_RNIE7KM6Z0Z_17 ;
    wire \Commands_frame_decoder.source_CH3data_1_sqmuxa_0 ;
    wire \dron_frame_decoder_1.N_700_0 ;
    wire \dron_frame_decoder_1.drone_H_disp_front_8 ;
    wire \dron_frame_decoder_1.drone_H_disp_front_10 ;
    wire \pid_front.N_3_cascade_ ;
    wire \pid_front.m2_0_03_3_i_0_cascade_ ;
    wire \dron_frame_decoder_1.drone_H_disp_front_9 ;
    wire \pid_front.error_i_acumm_preregZ0Z_7 ;
    wire \pid_front.error_i_acumm_3_sqmuxa ;
    wire \pid_front.error_i_acumm_preregZ0Z_9 ;
    wire \pid_front.error_i_acumm_preregZ0Z_1 ;
    wire \pid_front.error_i_acumm_preregZ0Z_2 ;
    wire \pid_front.error_i_acumm16lto3 ;
    wire \pid_front.error_i_acumm_prereg_esr_RNIV9S71Z0Z_12 ;
    wire \pid_front.error_i_acumm_2_sqmuxa_1_cascade_ ;
    wire \pid_front.error_i_acumm_prereg_esr_RNI0I2H5Z0Z_12 ;
    wire \pid_front.error_i_acumm_2_sqmuxa_cascade_ ;
    wire \pid_front.error_i_acumm_preregZ0Z_10 ;
    wire \pid_front.error_i_acumm_preregZ0Z_4 ;
    wire \pid_front.error_i_acumm_preregZ0Z_5 ;
    wire \pid_front.error_i_acumm_preregZ0Z_6 ;
    wire \pid_front.error_i_acumm_preregZ0Z_11 ;
    wire \pid_front.error_i_acumm_2_sqmuxa_1 ;
    wire \pid_front.error_i_acumm_2_sqmuxa ;
    wire \pid_front.error_p_reg_esr_RNI2BC9_0Z0Z_1_cascade_ ;
    wire \pid_front.error_d_reg_prev_esr_RNIFSHOZ0Z_1_cascade_ ;
    wire \pid_front.error_d_reg_prev_esr_RNID19M1Z0Z_1 ;
    wire \pid_front.error_p_reg_esr_RNIO4E8_0Z0Z_2 ;
    wire \pid_front.error_d_reg_prev_esr_RNIFSHOZ0Z_1 ;
    wire \pid_front.error_d_reg_prev_esr_RNI1JN71Z0Z_1 ;
    wire \pid_front.error_p_regZ0Z_1 ;
    wire \pid_front.error_p_reg_esr_RNI2BC9Z0Z_1 ;
    wire \pid_front.error_d_regZ0Z_0 ;
    wire \pid_front.error_d_reg_prevZ0Z_0 ;
    wire \pid_front.error_d_reg_prev_esr_RNIQHN6Z0Z_1 ;
    wire \pid_front.error_d_regZ0Z_1 ;
    wire \pid_front.error_d_reg_prevZ0Z_1 ;
    wire \pid_front.error_i_acumm_preregZ0Z_21 ;
    wire \pid_front.error_i_acumm_preregZ0Z_8 ;
    wire \pid_front.error_i_acumm_preregZ0Z_16 ;
    wire \pid_front.error_i_acumm_preregZ0Z_20 ;
    wire \pid_front.un10lto12 ;
    wire \pid_front.error_i_acumm16lto27_10 ;
    wire \pid_front.error_i_acumm16lto27_9 ;
    wire \pid_front.error_i_acumm16lto27_7_cascade_ ;
    wire \pid_front.error_i_acumm16lto27_8 ;
    wire \pid_front.error_i_acumm16lto27_13 ;
    wire \pid_front.error_i_acumm_preregZ0Z_22 ;
    wire \pid_front.error_i_acumm_preregZ0Z_24 ;
    wire \pid_front.error_i_acumm_preregZ0Z_13 ;
    wire \pid_front.un10lto27_8_cascade_ ;
    wire \pid_front.un10lto27_11 ;
    wire \pid_front.error_i_acumm_preregZ0Z_26 ;
    wire \ppm_encoder_1.elevatorZ0Z_11 ;
    wire \ppm_encoder_1.elevator_RNIPFGEZ0Z_11_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_0_2_11_cascade_ ;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_11_cascade_ ;
    wire \ppm_encoder_1.init_pulses_RNI4JPF5Z0Z_11 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_11 ;
    wire \ppm_encoder_1.N_266_i_i ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_4 ;
    wire \ppm_encoder_1.un1_init_pulses_11_13 ;
    wire \ppm_encoder_1.un1_init_pulses_10_13 ;
    wire \ppm_encoder_1.un1_init_pulses_11_2 ;
    wire \ppm_encoder_1.un1_init_pulses_10_2 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1 ;
    wire \ppm_encoder_1.elevatorZ0Z_3 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1 ;
    wire \ppm_encoder_1.pulses2count_9_0_0_0_3_cascade_ ;
    wire \ppm_encoder_1.init_pulsesZ0Z_3 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_0_0_cascade_ ;
    wire \ppm_encoder_1.throttle_RNI25564Z0Z_0 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_1_0 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_0_0 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_1_0_cascade_ ;
    wire throttle_order_0;
    wire \ppm_encoder_1.aileronZ0Z_0 ;
    wire \ppm_encoder_1.throttleZ0Z_0 ;
    wire front_order_0;
    wire \ppm_encoder_1.un2_throttle_iv_i_i_0_14_cascade_ ;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_14_cascade_ ;
    wire \ppm_encoder_1.init_pulses_RNIE8336Z0Z_14 ;
    wire \ppm_encoder_1.PPM_STATE_RNIV4V5Z0Z_1_cascade_ ;
    wire \ppm_encoder_1.N_269_i_i ;
    wire \ppm_encoder_1.N_269_i ;
    wire \ppm_encoder_1.counter24_0_I_57_c_RNIJMMDZ0 ;
    wire \ppm_encoder_1.aileronZ0Z_1 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIHO7DZ0Z_0_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_0_1_10 ;
    wire \ppm_encoder_1.throttleZ0Z_2 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIJQ7DZ0Z_1_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_0_0_1_7_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_0_0_0_7 ;
    wire \ppm_encoder_1.N_263_i_i ;
    wire \ppm_encoder_1.N_263_i_i_cascade_ ;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_7 ;
    wire \ppm_encoder_1.init_pulses_RNI2VJU5Z0Z_7 ;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_13_cascade_ ;
    wire \ppm_encoder_1.N_268_i_i ;
    wire \ppm_encoder_1.init_pulses_RNIFVPF5Z0Z_13 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_1_13 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_0_13 ;
    wire \ppm_encoder_1.elevator_RNIRHGEZ0Z_13 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_13 ;
    wire scaler_4_data_13;
    wire \ppm_encoder_1.un1_rudder_cry_12_THRU_CO ;
    wire \ppm_encoder_1.aileronZ0Z_7 ;
    wire \ppm_encoder_1.throttleZ0Z_7 ;
    wire \ppm_encoder_1.rudderZ0Z_11 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_11 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_3 ;
    wire \ppm_encoder_1.rudderZ0Z_13 ;
    wire \ppm_encoder_1.rudder_RNIN2KQZ0Z_13 ;
    wire side_order_5;
    wire side_order_7;
    wire side_order_3;
    wire side_order_11;
    wire side_order_1;
    wire side_order_0;
    wire side_order_10;
    wire side_order_4;
    wire side_order_8;
    wire side_order_9;
    wire \ppm_encoder_1.N_257_i_i ;
    wire frame_decoder_OFF4data_7;
    wire frame_decoder_CH4data_7;
    wire \scaler_4.N_2725_i_l_ofxZ0 ;
    wire \pid_side.error_p_reg_esr_RNISPTC1Z0Z_8_cascade_ ;
    wire \pid_side.error_p_reg_esr_RNISPTC1Z0Z_8 ;
    wire \pid_side.error_p_reg_esr_RNI1VTC1_0Z0Z_9 ;
    wire \pid_side.N_2374_i ;
    wire \pid_side.error_d_reg_prevZ0Z_7 ;
    wire \pid_side.N_2374_i_cascade_ ;
    wire \pid_side.error_d_reg_prevZ0Z_8 ;
    wire \pid_side.error_i_reg_esr_RNO_0Z0Z_22_cascade_ ;
    wire \pid_side.m36_1_ns_1 ;
    wire \pid_side.N_37_1_cascade_ ;
    wire \pid_side.N_39_1_cascade_ ;
    wire \pid_side.N_126_0_cascade_ ;
    wire \pid_side.m2_0_03_3_i_0_cascade_ ;
    wire \pid_side.N_41_0 ;
    wire \pid_side.N_41_0_cascade_ ;
    wire \pid_side.error_i_reg_9_rn_0_26_cascade_ ;
    wire \pid_side.m6_2_03_cascade_ ;
    wire \pid_side.N_39_1 ;
    wire \pid_side.error_i_reg_9_rn_0_18_cascade_ ;
    wire drone_H_disp_side_2;
    wire drone_H_disp_side_3;
    wire \dron_frame_decoder_1.N_724_0 ;
    wire \pid_alt.error_axbZ0Z_2 ;
    wire drone_altitude_2;
    wire \pid_alt.error_axbZ0Z_3 ;
    wire drone_altitude_3;
    wire \dron_frame_decoder_1.N_740_0 ;
    wire drone_H_disp_side_1;
    wire xy_kd_2;
    wire xy_kd_6;
    wire \dron_frame_decoder_1.drone_altitude_11 ;
    wire drone_altitude_i_11;
    wire \pid_front.error_d_reg_prevZ0Z_14 ;
    wire \pid_front.error_p_regZ0Z_14 ;
    wire \pid_front.error_p_reg_esr_RNIH0C61_0Z0Z_14 ;
    wire front_command_7;
    wire drone_H_disp_front_11;
    wire \pid_front.error_axb_0 ;
    wire bfn_13_21_0_;
    wire \pid_front.error_axbZ0Z_1 ;
    wire \pid_front.error_cry_0 ;
    wire \pid_front.error_axbZ0Z_2 ;
    wire \pid_front.error_cry_1 ;
    wire \pid_front.error_axbZ0Z_3 ;
    wire \pid_front.error_cry_2 ;
    wire drone_H_disp_front_i_4;
    wire front_command_0;
    wire \pid_front.error_cry_3 ;
    wire drone_H_disp_front_i_5;
    wire front_command_1;
    wire \pid_front.error_cry_0_0 ;
    wire drone_H_disp_front_i_6;
    wire front_command_2;
    wire \pid_front.error_cry_1_0 ;
    wire drone_H_disp_front_i_7;
    wire front_command_3;
    wire \pid_front.error_cry_2_0 ;
    wire \pid_front.error_cry_3_0 ;
    wire drone_H_disp_front_i_8;
    wire front_command_4;
    wire bfn_13_22_0_;
    wire drone_H_disp_front_i_9;
    wire front_command_5;
    wire \pid_front.error_cry_4 ;
    wire front_command_6;
    wire drone_H_disp_front_i_10;
    wire \pid_front.error_cry_5 ;
    wire \pid_front.error_axbZ0Z_7 ;
    wire \pid_front.error_cry_6 ;
    wire \pid_front.error_axb_8_l_ofx_0 ;
    wire drone_H_disp_front_12;
    wire \pid_front.error_cry_7 ;
    wire drone_H_disp_front_i_12;
    wire drone_H_disp_front_13;
    wire \pid_front.error_cry_8 ;
    wire drone_H_disp_front_i_13;
    wire \pid_front.error_cry_9 ;
    wire drone_H_disp_front_15;
    wire drone_H_disp_front_14;
    wire \pid_front.error_cry_10 ;
    wire \pid_front.un1_pid_prereg_0 ;
    wire bfn_13_23_0_;
    wire \pid_front.error_i_acummZ0Z_1 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_0_c_RNI9AGE ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_0 ;
    wire \pid_front.error_i_acummZ0Z_2 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_1_c_RNICEHE ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_1 ;
    wire \pid_front.error_i_acummZ0Z_3 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_2_c_RNIFIIE ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_2 ;
    wire \pid_front.error_i_acummZ0Z_4 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_3_c_RNIIMJE ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_3 ;
    wire \pid_front.error_i_acummZ0Z_5 ;
    wire \pid_front.error_i_regZ0Z_5 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_4_c_RNICGQM ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_4 ;
    wire \pid_front.error_i_acummZ0Z_6 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_5_c_RNIOULE ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_5 ;
    wire \pid_front.error_i_acummZ0Z_7 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_6_c_RNIR2NE ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_6 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_7 ;
    wire \pid_front.error_i_acummZ0Z_8 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_7_c_RNIU6OE ;
    wire bfn_13_24_0_;
    wire \pid_front.error_i_acummZ0Z_9 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_8_c_RNI1BPE ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_8 ;
    wire \pid_front.error_i_acummZ0Z_10 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_9_c_RNIIPQK ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_9 ;
    wire \pid_front.error_i_acummZ0Z_11 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_10_c_RNIJD4S ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_10 ;
    wire \pid_front.error_i_acummZ0Z_12 ;
    wire \pid_front.error_i_reg_esr_RNIV4AUZ0Z_12 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_11 ;
    wire \pid_front.error_i_reg_esr_RNI29BUZ0Z_13 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_12 ;
    wire \pid_front.error_i_reg_esr_RNI4CCUZ0Z_14 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_13 ;
    wire \pid_front.error_i_reg_esr_RNI6FDUZ0Z_15 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_14 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_15 ;
    wire \pid_front.error_i_reg_esr_RNI8IEUZ0Z_16 ;
    wire bfn_13_25_0_;
    wire \pid_front.un1_error_i_acumm_prereg_cry_16 ;
    wire \pid_front.error_i_reg_esr_RNICOGUZ0Z_18 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_17 ;
    wire \pid_front.error_i_reg_esr_RNIERHUZ0Z_19 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_18 ;
    wire \pid_front.error_i_reg_esr_RNI7MJUZ0Z_20 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_19 ;
    wire \pid_front.error_i_reg_esr_RNI08DVZ0Z_21 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_20 ;
    wire \pid_front.error_i_reg_esr_RNI2BEVZ0Z_22 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_21 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_22 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_23 ;
    wire \pid_front.error_i_reg_esr_RNI6HGVZ0Z_24 ;
    wire bfn_13_26_0_;
    wire \pid_front.un1_error_i_acumm_prereg_cry_24 ;
    wire \pid_front.error_i_reg_esr_RNIANIVZ0Z_26 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_25 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_26 ;
    wire \pid_front.error_i_acummZ0Z_13 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_27 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_27_c_RNIDSKV ;
    wire \pid_front.error_i_acumm_preregZ0Z_28 ;
    wire \pid_front.error_i_reg_esr_RNI8KHVZ0Z_25 ;
    wire \pid_front.error_i_acumm_preregZ0Z_25 ;
    wire \pid_front.error_i_reg_esr_RNI4EFVZ0Z_23 ;
    wire \pid_front.error_i_acumm_preregZ0Z_23 ;
    wire \pid_front.un1_error_i_acumm_prereg_cry_26_c_RNICQJV ;
    wire \pid_front.error_i_acumm_preregZ0Z_27 ;
    wire \pid_front.error_i_reg_esr_RNIALFUZ0Z_17 ;
    wire \pid_front.error_i_acumm_preregZ0Z_17 ;
    wire \pid_front.error_i_acummZ0Z_0 ;
    wire \pid_front.error_i_acumm_preregZ0Z_0 ;
    wire \pid_front.N_764_g ;
    wire \pid_alt.stateZ0Z_0 ;
    wire \pid_alt.state_0_0 ;
    wire \ppm_encoder_1.un1_init_pulses_11_0 ;
    wire \ppm_encoder_1.un1_init_pulses_10_0 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_RNIB7481Z0Z_3 ;
    wire \ppm_encoder_1.counter24_0_I_57_c_RNIV9SJZ0Z1 ;
    wire bfn_14_2_0_;
    wire \ppm_encoder_1.counter24_0_data_tmp_0 ;
    wire \ppm_encoder_1.counter24_0_data_tmp_1 ;
    wire \ppm_encoder_1.counter24_0_data_tmp_2 ;
    wire \ppm_encoder_1.counter24_0_data_tmp_3 ;
    wire \ppm_encoder_1.counter24_0_data_tmp_4 ;
    wire \ppm_encoder_1.counter24_0_data_tmp_5 ;
    wire \ppm_encoder_1.counter24_0_data_tmp_6 ;
    wire \ppm_encoder_1.counter24_0_data_tmp_7 ;
    wire bfn_14_3_0_;
    wire CONSTANT_ONE_NET;
    wire \ppm_encoder_1.counter24_0_data_tmp_8 ;
    wire \ppm_encoder_1.counter24_0_N_2 ;
    wire \ppm_encoder_1.aileronZ0Z_10 ;
    wire \ppm_encoder_1.elevatorZ0Z_10 ;
    wire \ppm_encoder_1.counter24_0_I_57_c_RNOZ0 ;
    wire \ppm_encoder_1.N_258_i_i ;
    wire \ppm_encoder_1.N_258_i_i_cascade_ ;
    wire \ppm_encoder_1.init_pulses_RNI40GS4Z0Z_1 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_7 ;
    wire \ppm_encoder_1.PPM_STATE_RNI5C4LZ0Z_1_cascade_ ;
    wire \ppm_encoder_1.aileron_RNIFUAPZ0Z_1 ;
    wire \ppm_encoder_1.init_pulses_RNI7A1R_0Z0Z_1_cascade_ ;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_1 ;
    wire \ppm_encoder_1.N_56 ;
    wire \ppm_encoder_1.throttleZ0Z_11 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_1_11 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIM4C21Z0Z_2 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIM4C21Z0Z_2_cascade_ ;
    wire \ppm_encoder_1.init_pulses_RNIN1203Z0Z_2 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIIP7DZ0Z_0 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI5QE01Z0Z_3 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_1_2 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_2_2_cascade_ ;
    wire \ppm_encoder_1.PPM_STATE_RNI5C4LZ0Z_1 ;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_2_cascade_ ;
    wire \ppm_encoder_1.init_pulses_RNI5GAI5Z0Z_2 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_3_repZ0Z1 ;
    wire \ppm_encoder_1.N_259_i_i ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_1 ;
    wire \ppm_encoder_1.throttleZ0Z_14 ;
    wire \ppm_encoder_1.aileronZ0Z_14 ;
    wire \ppm_encoder_1.pulses2count_9_i_0_14_cascade_ ;
    wire \ppm_encoder_1.init_pulsesZ0Z_14 ;
    wire \ppm_encoder_1.pulses2count_9_i_1_14_cascade_ ;
    wire \ppm_encoder_1.elevator_esr_RNI6C0M1Z0Z_14 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_ns_0 ;
    wire \ppm_encoder_1.elevatorZ0Z_2 ;
    wire \ppm_encoder_1.elevatorZ0Z_1 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIJQ7DZ0Z_1 ;
    wire \ppm_encoder_1.throttleZ0Z_1 ;
    wire \ppm_encoder_1.throttle_RNI2JJC1Z0Z_1 ;
    wire \ppm_encoder_1.counter24_0_I_21_c_RNOZ0 ;
    wire \ppm_encoder_1.rudderZ0Z_7 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_2Z0Z_7 ;
    wire \ppm_encoder_1.elevator_RNIEB6OZ0Z_7 ;
    wire \ppm_encoder_1.pulses2count_9_i_0_7 ;
    wire \ppm_encoder_1.pulses2count_9_i_2_7_cascade_ ;
    wire \ppm_encoder_1.pulses2countZ0Z_7 ;
    wire \ppm_encoder_1.rudderZ0Z_6 ;
    wire \ppm_encoder_1.elevator_RNIDA6OZ0Z_6 ;
    wire \ppm_encoder_1.pulses2count_9_0_2_6_cascade_ ;
    wire \ppm_encoder_1.pulses2countZ0Z_6 ;
    wire \ppm_encoder_1.pulses2count_9_0_2_13 ;
    wire side_order_6;
    wire side_order_2;
    wire \pid_side.un1_reset_0_i_cascade_ ;
    wire \pid_side.N_75 ;
    wire \pid_side.N_75_cascade_ ;
    wire \pid_side.N_102 ;
    wire \pid_side.N_76 ;
    wire side_order_12;
    wire side_order_13;
    wire \pid_side.state_0_1 ;
    wire \pid_side.un1_reset_0_i ;
    wire \pid_side.state_ns_0_cascade_ ;
    wire \pid_side.error_i_acumm_prereg_esr_RNIGSJVZ0Z_7_cascade_ ;
    wire \pid_side.error_i_acumm_prereg_esr_RNIJ04N_0Z0Z_10 ;
    wire \pid_side.error_p_reg_esr_RNINKTC1_0Z0Z_7_cascade_ ;
    wire \pid_side.N_2362_i_cascade_ ;
    wire \pid_side.error_p_reg_esr_RNIIFTC1Z0Z_6 ;
    wire \pid_side.error_p_reg_esr_RNIIFTC1Z0Z_6_cascade_ ;
    wire \pid_side.error_p_reg_esr_RNINKTC1_0Z0Z_7 ;
    wire \pid_side.N_2368_i ;
    wire \pid_side.error_d_reg_prevZ0Z_6 ;
    wire \pid_side.error_p_reg_esr_RNINKTC1Z0Z_7_cascade_ ;
    wire \pid_side.error_i_reg_9_rn_0_19_cascade_ ;
    wire \pid_side.m2_2_03_cascade_ ;
    wire \pid_side.g1 ;
    wire \pid_side.g3_cascade_ ;
    wire \pid_side.m37_1_ns_1_cascade_ ;
    wire \pid_side.N_38_1_cascade_ ;
    wire \pid_side.error_i_reg_esr_RNO_3Z0Z_22_cascade_ ;
    wire \pid_side.error_i_reg_esr_RNO_2Z0Z_22 ;
    wire \pid_side.error_i_reg_esr_RNO_1Z0Z_22 ;
    wire \pid_side.N_37_1 ;
    wire \pid_side.m136_ns_1_cascade_ ;
    wire \pid_side.m18_2_03_4 ;
    wire \pid_side.error_cry_1_0_c_RNIEAJZ0Z82 ;
    wire \pid_side.error_cry_1_0_c_RNIEAJ82Z0Z_0_cascade_ ;
    wire \pid_side.N_39_0_cascade_ ;
    wire \pid_side.m7_2_03 ;
    wire \pid_side.m134_0_ns_1_cascade_ ;
    wire \pid_side.m19_2_03_0_cascade_ ;
    wire \pid_side.error_cry_5_c_RNIN1DBZ0Z2_cascade_ ;
    wire \pid_side.error_cry_5_c_RNIN1DB2Z0Z_0 ;
    wire \pid_side.N_103_0_cascade_ ;
    wire \pid_side.N_53_0 ;
    wire \pid_side.N_50_1_cascade_ ;
    wire \pid_side.N_50_1 ;
    wire \pid_side.error_i_reg_9_rn_0_27 ;
    wire \dron_frame_decoder_1.drone_H_disp_side_4 ;
    wire \dron_frame_decoder_1.drone_H_disp_side_5 ;
    wire \dron_frame_decoder_1.drone_H_disp_side_6 ;
    wire \dron_frame_decoder_1.drone_H_disp_side_7 ;
    wire \pid_side.N_88_0_0 ;
    wire uart_drone_data_1;
    wire drone_H_disp_front_1;
    wire uart_drone_data_2;
    wire drone_H_disp_front_2;
    wire uart_drone_data_3;
    wire drone_H_disp_front_3;
    wire uart_drone_data_4;
    wire \dron_frame_decoder_1.drone_H_disp_front_4 ;
    wire uart_drone_data_5;
    wire \dron_frame_decoder_1.drone_H_disp_front_5 ;
    wire uart_drone_data_6;
    wire \dron_frame_decoder_1.drone_H_disp_front_6 ;
    wire uart_drone_data_7;
    wire \dron_frame_decoder_1.drone_H_disp_front_7 ;
    wire \pid_front.m0_0_03_cascade_ ;
    wire uart_drone_data_0;
    wire dron_frame_decoder_1_source_H_disp_front_fast_0;
    wire \dron_frame_decoder_1.N_708_0 ;
    wire \pid_side.un4_error_i_reg_31_ns_1_0 ;
    wire \pid_front.m11_0_ns_1 ;
    wire \pid_front.N_48_1_cascade_ ;
    wire \pid_front.error_cry_1_0_c_RNIOOIF3Z0Z_0_cascade_ ;
    wire \pid_front.N_116_0_cascade_ ;
    wire \pid_front.error_cry_1_0_c_RNIOOIFZ0Z3 ;
    wire \pid_front.N_21_1 ;
    wire \pid_front.error_cry_6_c_RNI1ADU1Z0Z_0_cascade_ ;
    wire \pid_front.error_cry_6_c_RNI1ADUZ0Z1 ;
    wire \pid_front.m4_2_03 ;
    wire \pid_front.error_i_reg_9_rn_0_16_cascade_ ;
    wire \pid_front.error_i_regZ0Z_16 ;
    wire \pid_front.error_i_reg_esr_RNO_0Z0Z_16 ;
    wire \pid_front.N_36_0_cascade_ ;
    wire \pid_front.N_37_1_cascade_ ;
    wire \pid_front.N_18_1 ;
    wire \pid_front.error_i_reg_esr_RNO_2_0_16 ;
    wire \pid_front.error_i_reg_esr_RNO_4Z0Z_21_cascade_ ;
    wire \pid_front.g0_5_1 ;
    wire \pid_front.N_126_0_cascade_ ;
    wire \pid_front.N_88_0_0 ;
    wire \pid_front.m25_2_03_0_cascade_ ;
    wire \pid_front.m9_2_03_3_i_0 ;
    wire \pid_front.error_i_regZ0Z_21 ;
    wire \pid_front.error_i_regZ0Z_12 ;
    wire \pid_front.error_i_regZ0Z_18 ;
    wire \pid_front.error_9 ;
    wire \pid_front.N_25_0 ;
    wire \pid_front.error_cry_4_c_RNI81RMZ0Z1_cascade_ ;
    wire \pid_front.error_cry_4_c_RNI81RM1Z0Z_0 ;
    wire \pid_front.N_38_1_cascade_ ;
    wire \pid_front.N_37_1 ;
    wire \pid_front.N_39_1_cascade_ ;
    wire \pid_front.error_i_regZ0Z_10 ;
    wire \pid_front.N_38_1 ;
    wire \pid_front.N_110_cascade_ ;
    wire \pid_front.m2_2_03 ;
    wire \pid_front.error_i_reg_9_rn_1_14_cascade_ ;
    wire \pid_front.N_136 ;
    wire \pid_front.error_i_regZ0Z_14 ;
    wire \pid_front.m10_2_03_3_i_0_cascade_ ;
    wire \pid_front.m26_2_03_0 ;
    wire \pid_front.error_i_regZ0Z_22 ;
    wire \pid_front.stateZ0Z_0 ;
    wire \pid_front.stateZ0Z_1 ;
    wire \pid_front.N_196_mux_cascade_ ;
    wire \pid_front.error_i_acumm_1_sqmuxa_1_i ;
    wire pid_side_m153_e_5;
    wire debug_CH1_0A_c;
    wire pid_side_m153_e_5_cascade_;
    wire \pid_side.stateZ0Z_0 ;
    wire \pid_side.N_196_mux ;
    wire \ppm_encoder_1.counter24_0_I_15_c_RNOZ0 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_2Z0Z_4 ;
    wire \ppm_encoder_1.rudderZ0Z_4 ;
    wire \ppm_encoder_1.pulses2count_9_i_1_4 ;
    wire \ppm_encoder_1.pulses2count_9_i_2_4_cascade_ ;
    wire \ppm_encoder_1.init_pulsesZ0Z_4 ;
    wire \ppm_encoder_1.pulses2countZ0Z_4 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_5 ;
    wire \ppm_encoder_1.elevator_RNIC96OZ0Z_5 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_2Z0Z_5_cascade_ ;
    wire \ppm_encoder_1.rudderZ0Z_5 ;
    wire \ppm_encoder_1.pulses2count_9_i_0_5 ;
    wire \ppm_encoder_1.pulses2count_9_i_2_5_cascade_ ;
    wire \ppm_encoder_1.pulses2countZ0Z_5 ;
    wire \ppm_encoder_1.pulses2count_9_0_0_0 ;
    wire \ppm_encoder_1.pulses2countZ0Z_13 ;
    wire \ppm_encoder_1.counter24_0_I_39_c_RNOZ0 ;
    wire \ppm_encoder_1.aileronZ0Z_12 ;
    wire \ppm_encoder_1.pulses2count_9_0_3_12 ;
    wire \ppm_encoder_1.pulses2countZ0Z_12 ;
    wire \ppm_encoder_1.pulses2count_9_0_3_11 ;
    wire \ppm_encoder_1.aileronZ0Z_11 ;
    wire \ppm_encoder_1.counter24_0_I_9_c_RNOZ0 ;
    wire \ppm_encoder_1.counter24_0_I_27_c_RNOZ0 ;
    wire \ppm_encoder_1.pulses2count_9_i_1_8 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_8 ;
    wire \ppm_encoder_1.pulses2countZ0Z_8 ;
    wire \ppm_encoder_1.pulses2count_9_i_1_9 ;
    wire \ppm_encoder_1.pulses2countZ0Z_9 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_18 ;
    wire \ppm_encoder_1.pulses2countZ0Z_18 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_10 ;
    wire \ppm_encoder_1.pulses2count_9_i_0_1_10 ;
    wire \ppm_encoder_1.pulses2countZ0Z_10 ;
    wire \ppm_encoder_1.pulses2countZ0Z_11 ;
    wire \ppm_encoder_1.counter24_0_I_33_c_RNOZ0 ;
    wire \ppm_encoder_1.ppm_output_reg_RNOZ0Z_0 ;
    wire \ppm_encoder_1.un1_PPM_STATE_0_sqmuxa_0_i_a2_18_10 ;
    wire \ppm_encoder_1.un1_PPM_STATE_0_sqmuxa_0_i_a2_18_11_cascade_ ;
    wire \ppm_encoder_1.un1_PPM_STATE_0_sqmuxa_0_i_a2_18_8 ;
    wire \ppm_encoder_1.N_486_18 ;
    wire \ppm_encoder_1.N_486_9 ;
    wire \ppm_encoder_1.N_486_18_cascade_ ;
    wire \ppm_encoder_1.PPM_STATEZ0Z_1 ;
    wire \ppm_encoder_1.counter_RNI09RH2Z0Z_18 ;
    wire \ppm_encoder_1.PPM_STATEZ0Z_0 ;
    wire \ppm_encoder_1.counter24_0_N_2_THRU_CO ;
    wire \ppm_encoder_1.counter_RNI09RH2Z0Z_18_cascade_ ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_17 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_3_repZ0Z2 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z2 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_3_rep2_RNIAZ0Z6041_cascade_ ;
    wire \ppm_encoder_1.rudderZ0Z_10 ;
    wire \ppm_encoder_1.pulses2count_9_i_0_2_10 ;
    wire \ppm_encoder_1.throttleZ0Z_10 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_2Z0Z_10 ;
    wire \ppm_encoder_1.throttleZ0Z_8 ;
    wire \ppm_encoder_1.rudderZ0Z_8 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_2Z0Z_8_cascade_ ;
    wire \ppm_encoder_1.pulses2count_9_i_2_8 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_2Z0Z_9 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_3_rep2_RNIAZ0Z6041 ;
    wire \ppm_encoder_1.rudderZ0Z_9 ;
    wire \ppm_encoder_1.pulses2count_9_i_2_9 ;
    wire \ppm_encoder_1.throttleZ0Z_6 ;
    wire \ppm_encoder_1.aileronZ0Z_6 ;
    wire \ppm_encoder_1.pulses2count_9_0_0_6 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_6 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_2Z0Z_6 ;
    wire \ppm_encoder_1.CHOOSE_CHANNELZ0Z_0 ;
    wire \ppm_encoder_1.throttleZ0Z_13 ;
    wire \ppm_encoder_1.CHOOSE_CHANNELZ0Z_1 ;
    wire \ppm_encoder_1.aileronZ0Z_13 ;
    wire \ppm_encoder_1.pulses2count_9_0_0_13 ;
    wire \pid_side.source_pid10lt4_0 ;
    wire bfn_15_8_0_;
    wire \pid_side.un11lto30_i_a2_0_and ;
    wire \pid_side.un11lto30_i_a2 ;
    wire \pid_side.N_11_i ;
    wire \pid_side.un11lto30_i_a2_0 ;
    wire \pid_side.un11lto30_i_a2_2_and ;
    wire \pid_side.un11lto30_i_a2_1 ;
    wire \pid_side.un11lto30_i_a2_2 ;
    wire \pid_side.un11lto30_i_a2_3 ;
    wire \pid_side.un11lto30_i_a2_4 ;
    wire \pid_side.un11lto30_i_a2_5 ;
    wire \pid_side.un11lto30_i_a2_6 ;
    wire bfn_15_9_0_;
    wire \pid_side.source_pid_1_sqmuxa_1_0_o2_sx ;
    wire \pid_side.N_389 ;
    wire \pid_side.source_pid_1_sqmuxa_1_0_a4_3 ;
    wire \pid_side.un11lto30_i_a2_5_and ;
    wire \pid_side.un11lto30_i_a2_6_and ;
    wire \pid_side.un11lto30_i_a2_5_and_cascade_ ;
    wire \pid_side.un11lto30_i_a2_4_and ;
    wire \pid_side.N_98 ;
    wire \pid_side.error_i_acumm_preregZ0Z_10 ;
    wire \pid_side.un10lt9_1_cascade_ ;
    wire \pid_side.error_i_acumm16lt9_0 ;
    wire \pid_side.un10lt9_1 ;
    wire \pid_side.un10lt9_cascade_ ;
    wire \pid_side.error_i_acumm_prereg_esr_RNIJ04NZ0Z_10 ;
    wire \pid_side.un10lt11_0_cascade_ ;
    wire \pid_side.error_i_acumm_preregZ0Z_7 ;
    wire \pid_side.error_i_acumm_preregZ0Z_8 ;
    wire \pid_side.error_i_acumm_preregZ0Z_0 ;
    wire \pid_side.error_p_reg_esr_RNISPTC1_0Z0Z_8 ;
    wire \pid_side.error_p_reg_esr_RNINKTC1Z0Z_7 ;
    wire \uart_drone.bit_CountZ0Z_2 ;
    wire \uart_drone.bit_CountZ0Z_1 ;
    wire \uart_drone.bit_CountZ0Z_0 ;
    wire \uart_drone.data_Auxce_0_0_0 ;
    wire \pid_side.N_15_0_cascade_ ;
    wire \pid_side.m4_2_03_cascade_ ;
    wire \pid_side.N_30_1 ;
    wire \pid_side.N_30_1_cascade_ ;
    wire \pid_side.N_63_cascade_ ;
    wire \pid_side.m2_0_03_3_i_0 ;
    wire \pid_side.un1_pid_prereg_0_23_cascade_ ;
    wire \pid_side.un1_pid_prereg_0_22_cascade_ ;
    wire \pid_side.un1_pid_prereg_0_23 ;
    wire \pid_side.un1_pid_prereg_0_22 ;
    wire \pid_side.un1_pid_prereg_0_24_cascade_ ;
    wire \pid_side.N_11_0_cascade_ ;
    wire \pid_side.N_15_1_cascade_ ;
    wire \pid_side.m3_2_03 ;
    wire \pid_side.N_15_1 ;
    wire \pid_side.N_63 ;
    wire \pid_side.N_38_1 ;
    wire \pid_side.N_55_0 ;
    wire \pid_side.N_110_cascade_ ;
    wire \pid_side.N_3 ;
    wire \pid_side.N_14_1 ;
    wire \pid_side.N_104 ;
    wire \pid_side.N_104_cascade_ ;
    wire \pid_side.N_49_0 ;
    wire \pid_side.un4_error_i_reg_33_bm_1_cascade_ ;
    wire \pid_side.N_39_0 ;
    wire \pid_side.error_i_reg_esr_RNO_1Z0Z_23_cascade_ ;
    wire \pid_side.error_cry_9_c_RNIL6R82Z0Z_0_cascade_ ;
    wire \pid_side.N_46_1 ;
    wire \pid_side.N_46_1_cascade_ ;
    wire \pid_side.error_i_reg_esr_RNO_0Z0Z_23 ;
    wire \pid_side.error_cry_9_c_RNIL6RZ0Z82 ;
    wire \pid_side.N_27_1 ;
    wire \pid_side.error_cry_3_0_c_RNIJIPSZ0Z1_cascade_ ;
    wire \pid_side.error_cry_3_0_c_RNIJIPS1Z0Z_0 ;
    wire \pid_side.N_28_1_cascade_ ;
    wire \pid_side.error_cry_0_c_RNI94FZ0Z58_cascade_ ;
    wire \pid_side.m8_2_03_3_i_0_cascade_ ;
    wire \pid_side.m24_2_03_0 ;
    wire \pid_side.G_5_0_a5_0_1_cascade_ ;
    wire \pid_side.N_9_cascade_ ;
    wire \pid_side.G_5_0_1 ;
    wire \pid_side.G_5_0_a5_2_0 ;
    wire \pid_side.N_45_1 ;
    wire \pid_side.m87_0_ns_1_0 ;
    wire GB_BUFFER_reset_system_g_THRU_CO;
    wire \pid_side.N_6_0 ;
    wire \pid_side.g2_cascade_ ;
    wire \pid_side.N_117_0 ;
    wire \pid_front.error_i_regZ0Z_2 ;
    wire \pid_front.error_i_regZ0Z_3 ;
    wire \pid_side.m1_0_03_cascade_ ;
    wire \pid_side.error_i_reg_esr_RNO_5Z0Z_17 ;
    wire \pid_side.error_i_reg_esr_RNO_4Z0Z_17 ;
    wire \pid_side.N_131_cascade_ ;
    wire \pid_side.m5_2_03 ;
    wire \pid_front.N_63_cascade_ ;
    wire \pid_front.m6_2_03_cascade_ ;
    wire \pid_front.error_i_reg_9_rn_0_18 ;
    wire \pid_front.m2_0_03_3_i_0 ;
    wire \pid_front.N_63 ;
    wire \pid_front.N_41_0 ;
    wire \pid_front.N_41_0_cascade_ ;
    wire \pid_front.m129_0_ns_1_cascade_ ;
    wire \pid_front.m16_2_03_4 ;
    wire \pid_front.error_8 ;
    wire \pid_front.N_29_1_cascade_ ;
    wire \pid_front.error_cry_3_0_c_RNI76FZ0Z08_cascade_ ;
    wire \pid_front.N_27_1 ;
    wire \pid_front.error_cry_3_0_c_RNIJZ0Z5832 ;
    wire \pid_front.error_cry_3_0_c_RNIJ5832Z0Z_0 ;
    wire \pid_front.N_28_1 ;
    wire \pid_front.error_i_regZ0Z_0 ;
    wire \pid_front.N_36_0 ;
    wire \pid_front.N_57_0_cascade_ ;
    wire \pid_front.N_59_0_cascade_ ;
    wire \pid_front.N_89_i ;
    wire \pid_front.error_i_regZ0Z_24 ;
    wire \pid_front.N_3 ;
    wire \pid_front.N_30_1 ;
    wire \pid_front.N_15_0 ;
    wire \pid_front.N_15_0_cascade_ ;
    wire \pid_front.N_57_0 ;
    wire \pid_front.m138_0_1_cascade_ ;
    wire \pid_front.N_22_0 ;
    wire \pid_front.m0_0_03 ;
    wire \pid_front.m0_2_03 ;
    wire \pid_front.m24_2_03_0 ;
    wire \pid_front.m8_2_03_3_i_0 ;
    wire \pid_front.error_i_regZ0Z_20 ;
    wire \pid_front.N_39_1 ;
    wire \pid_front.error_i_reg_9_rn_0_26 ;
    wire \pid_front.error_i_regZ0Z_26 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_16 ;
    wire \ppm_encoder_1.m9_0_i ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIHO7DZ0Z_0 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z1 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNISSERZ0_cascade_ ;
    wire \ppm_encoder_1.init_pulsesZ0Z_1 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_0 ;
    wire \ppm_encoder_1.elevatorZ0Z_0 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_2Z0Z_0_cascade_ ;
    wire \ppm_encoder_1.m9_0_i_o2 ;
    wire \ppm_encoder_1.pulses2count_9_0_2_0 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_9 ;
    wire \ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_9 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_2 ;
    wire \ppm_encoder_1.pulses2count_9_i_0_2 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_2 ;
    wire \ppm_encoder_1.pulses2countZ0Z_0 ;
    wire \ppm_encoder_1.counter24_0_I_1_c_RNOZ0 ;
    wire \ppm_encoder_1.pulses2count_9_0_3_1 ;
    wire \ppm_encoder_1.pulses2count_9_0_0_1 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_1 ;
    wire \ppm_encoder_1.pulses2countZ0Z_1 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_15 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_17 ;
    wire \ppm_encoder_1.CHOOSE_CHANNELZ0Z_3 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNISSERZ0 ;
    wire \ppm_encoder_1.pulses2countZ0Z_16 ;
    wire \ppm_encoder_1.pulses2countZ0Z_17 ;
    wire \ppm_encoder_1.counter24_0_I_51_c_RNOZ0 ;
    wire \ppm_encoder_1.PPM_STATE_RNIV4V5Z0Z_1 ;
    wire \ppm_encoder_1.counterZ0Z_0 ;
    wire bfn_16_4_0_;
    wire \ppm_encoder_1.counterZ0Z_1 ;
    wire \ppm_encoder_1.un1_counter_13_cry_0 ;
    wire \ppm_encoder_1.un1_counter_13_cry_1 ;
    wire \ppm_encoder_1.un1_counter_13_cry_2 ;
    wire \ppm_encoder_1.counterZ0Z_4 ;
    wire \ppm_encoder_1.un1_counter_13_cry_3 ;
    wire \ppm_encoder_1.counterZ0Z_5 ;
    wire \ppm_encoder_1.un1_counter_13_cry_4 ;
    wire \ppm_encoder_1.counterZ0Z_6 ;
    wire \ppm_encoder_1.un1_counter_13_cry_5 ;
    wire \ppm_encoder_1.counterZ0Z_7 ;
    wire \ppm_encoder_1.un1_counter_13_cry_6 ;
    wire \ppm_encoder_1.un1_counter_13_cry_7 ;
    wire \ppm_encoder_1.counterZ0Z_8 ;
    wire bfn_16_5_0_;
    wire \ppm_encoder_1.counterZ0Z_9 ;
    wire \ppm_encoder_1.un1_counter_13_cry_8 ;
    wire \ppm_encoder_1.counterZ0Z_10 ;
    wire \ppm_encoder_1.un1_counter_13_cry_9 ;
    wire \ppm_encoder_1.counterZ0Z_11 ;
    wire \ppm_encoder_1.un1_counter_13_cry_10 ;
    wire \ppm_encoder_1.counterZ0Z_12 ;
    wire \ppm_encoder_1.un1_counter_13_cry_11 ;
    wire \ppm_encoder_1.counterZ0Z_13 ;
    wire \ppm_encoder_1.un1_counter_13_cry_12 ;
    wire \ppm_encoder_1.un1_counter_13_cry_13 ;
    wire \ppm_encoder_1.un1_counter_13_cry_14 ;
    wire \ppm_encoder_1.un1_counter_13_cry_15 ;
    wire bfn_16_6_0_;
    wire \ppm_encoder_1.un1_counter_13_cry_16 ;
    wire \ppm_encoder_1.un1_counter_13_cry_17 ;
    wire \ppm_encoder_1.counterZ0Z_18 ;
    wire \ppm_encoder_1.counter24_0_I_57_c_RNIGCOZ0Z83 ;
    wire \pid_alt.N_72_i ;
    wire pid_altitude_dv;
    wire \pid_alt.state_1_0_0 ;
    wire \pid_side.un10lto27_10_cascade_ ;
    wire \pid_side.error_i_acumm_prereg_esr_RNI5LOD5_0Z0Z_14 ;
    wire \pid_side.un10lto27_9 ;
    wire \pid_side.error_i_acumm_preregZ0Z_20 ;
    wire \pid_side.error_i_acumm_preregZ0Z_19 ;
    wire \pid_side.error_i_acumm_preregZ0Z_18 ;
    wire \pid_side.error_i_acumm16lto27_9 ;
    wire \pid_side.error_i_acumm16lto27_8_cascade_ ;
    wire \pid_side.error_i_acumm16lto27_7 ;
    wire \pid_side.error_i_acumm_preregZ0Z_15 ;
    wire \pid_side.error_i_acumm_preregZ0Z_14 ;
    wire \pid_side.error_i_acumm16lto27_10 ;
    wire \pid_side.un10lto27_8_cascade_ ;
    wire \pid_side.un10lto27_11 ;
    wire \pid_side.error_i_acumm_preregZ0Z_26 ;
    wire \pid_side.error_i_acumm_preregZ0Z_1 ;
    wire \pid_side.error_i_acumm_preregZ0Z_2 ;
    wire \pid_side.error_i_acumm16lto3 ;
    wire \pid_side.error_i_acumm_preregZ0Z_16 ;
    wire \pid_side.error_i_acumm_preregZ0Z_9 ;
    wire \pid_side.error_i_acumm_preregZ0Z_27 ;
    wire \pid_side.error_i_acumm_preregZ0Z_11 ;
    wire \pid_side.error_i_acumm_preregZ0Z_4 ;
    wire \pid_side.error_i_acumm_preregZ0Z_6 ;
    wire \pid_side.error_i_acumm_1_sqmuxa_1_i ;
    wire \pid_side.error_i_acumm16lto27_13 ;
    wire \pid_side.error_i_acumm_prereg_esr_RNIBT1C4Z0Z_12 ;
    wire reset_system;
    wire \pid_side.error_i_acumm_2_sqmuxa_1 ;
    wire \pid_side.error_i_acumm_2_sqmuxa_1_cascade_ ;
    wire \pid_side.error_i_acumm_prereg_esr_RNIGIQP9Z0Z_12 ;
    wire \pid_side.error_i_acumm_2_sqmuxa ;
    wire \pid_side.un1_pid_prereg_370_1_cascade_ ;
    wire \pid_side.un1_pid_prereg_0_14_cascade_ ;
    wire \pid_side.un1_pid_prereg_0_15_cascade_ ;
    wire \pid_side.un1_pid_prereg_0_24 ;
    wire \pid_side.un1_pid_prereg_0_26 ;
    wire \pid_side.un1_pid_prereg_0_25 ;
    wire \pid_side.error_i_acummZ0Z_0 ;
    wire \pid_side.error_i_regZ0Z_0 ;
    wire bfn_16_13_0_;
    wire \pid_side.error_i_acummZ0Z_1 ;
    wire \pid_side.error_i_regZ0Z_1 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_0 ;
    wire \pid_side.error_i_acummZ0Z_2 ;
    wire \pid_side.error_i_regZ0Z_2 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_1 ;
    wire \pid_side.error_i_acummZ0Z_3 ;
    wire \pid_side.error_i_regZ0Z_3 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_2 ;
    wire \pid_side.error_i_acummZ0Z_4 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_3 ;
    wire \pid_side.error_i_acummZ0Z_5 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_4 ;
    wire \pid_side.error_i_acummZ0Z_6 ;
    wire \pid_side.error_i_regZ0Z_6 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_5 ;
    wire \pid_side.error_i_acummZ0Z_7 ;
    wire \pid_side.error_i_regZ0Z_7 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_6_c_RNIF9RN ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_6 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_7 ;
    wire \pid_side.error_i_acummZ0Z_8 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_7_c_RNI9JMJ ;
    wire bfn_16_14_0_;
    wire \pid_side.error_i_acummZ0Z_9 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_8_c_RNILHTN ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_8 ;
    wire \pid_side.error_i_acummZ0Z_10 ;
    wire \pid_side.error_i_regZ0Z_10 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_9 ;
    wire \pid_side.error_i_acummZ0Z_11 ;
    wire \pid_side.error_i_regZ0Z_11 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_10 ;
    wire \pid_side.error_i_acummZ0Z_12 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_11 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_12 ;
    wire \pid_side.error_i_regZ0Z_14 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_13 ;
    wire \pid_side.error_i_regZ0Z_15 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_14 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_15 ;
    wire \pid_side.error_i_regZ0Z_16 ;
    wire bfn_16_15_0_;
    wire \pid_side.un1_error_i_acumm_prereg_cry_16 ;
    wire \pid_side.error_i_regZ0Z_18 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_17 ;
    wire \pid_side.error_i_regZ0Z_19 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_18 ;
    wire \pid_side.error_i_regZ0Z_20 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_19 ;
    wire \pid_side.error_i_regZ0Z_21 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_20 ;
    wire \pid_side.error_i_regZ0Z_22 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_21 ;
    wire \pid_side.error_i_regZ0Z_23 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_22 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_23 ;
    wire bfn_16_16_0_;
    wire \pid_side.un1_error_i_acumm_prereg_cry_24 ;
    wire \pid_side.error_i_regZ0Z_26 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_25 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_26_c_RNI0LUS ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_26 ;
    wire \pid_side.error_i_regZ0Z_27 ;
    wire \pid_side.error_i_acummZ0Z_13 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_27 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_27_c_RNI1NVS ;
    wire \pid_side.error_i_acumm_preregZ0Z_25 ;
    wire \pid_side.m32_0_ns_1_cascade_ ;
    wire \pid_side.N_89_i_cascade_ ;
    wire \pid_side.state_ns_0 ;
    wire \pid_side.error_i_regZ0Z_8 ;
    wire \pid_side.N_22_0_cascade_ ;
    wire \pid_side.N_22_0 ;
    wire \pid_side.error_i_reg_esr_RNO_4Z0Z_16_cascade_ ;
    wire \pid_side.error_i_reg_esr_RNO_3Z0Z_16 ;
    wire \pid_side.m20_2_03_0 ;
    wire \pid_side.N_11_0 ;
    wire \pid_side.N_12_1 ;
    wire \pid_side.N_12_1_cascade_ ;
    wire \pid_side.N_93_0_cascade_ ;
    wire \pid_side.un4_error_i_reg_35_am_1_cascade_ ;
    wire \pid_side.error_i_reg_esr_RNO_2_0_25 ;
    wire \pid_side.N_93_0 ;
    wire \pid_side.error_i_regZ0Z_9 ;
    wire pid_side_N_166_cascade_;
    wire \pid_side.error_cry_0_c_RNI94FZ0Z58 ;
    wire \pid_side.error_i_regZ0Z_4 ;
    wire \pid_side.error_i_reg_9_rn_1_17 ;
    wire \pid_side.error_i_regZ0Z_17 ;
    wire \pid_side.error_i_reg_9_rn_1_25 ;
    wire \pid_side.error_i_regZ0Z_25 ;
    wire \pid_side.m61_0_bmZ0 ;
    wire \pid_front.error_11 ;
    wire \pid_front.error_10 ;
    wire \pid_front.error_13 ;
    wire \pid_front.g0_15_1_cascade_ ;
    wire \pid_front.error_12 ;
    wire \pid_side.N_9_1_0 ;
    wire \pid_side.N_15_0 ;
    wire \pid_side.N_28_1 ;
    wire \pid_side.N_60_0_cascade_ ;
    wire \pid_side.error_i_reg_9_rn_1_12_cascade_ ;
    wire \pid_side.N_129 ;
    wire \pid_side.error_i_regZ0Z_12 ;
    wire \pid_front.error_4 ;
    wire \pid_front.error_5 ;
    wire \pid_front.error_6 ;
    wire \pid_front.error_7 ;
    wire \pid_front.N_9_1 ;
    wire \pid_front.error_cry_1_0_c_RNIDPRQ1Z0Z_0_cascade_ ;
    wire \pid_front.error_cry_1_0_c_RNIDPRQZ0Z1 ;
    wire xy_ki_fast_3;
    wire \pid_front.N_39_0_cascade_ ;
    wire \pid_front.m53_0_ns_1_cascade_ ;
    wire \pid_front.state_ns_0 ;
    wire \pid_front.N_54_0_cascade_ ;
    wire \pid_front.error_i_regZ0Z_11 ;
    wire \pid_front.N_54_0 ;
    wire \pid_front.error_i_regZ0Z_27 ;
    wire \pid_front.m7_2_03_cascade_ ;
    wire \pid_front.error_i_reg_9_rn_0_19_cascade_ ;
    wire \pid_front.error_i_regZ0Z_19 ;
    wire pid_front_error_i_reg_9_sn_19_cascade_;
    wire \pid_front.error_i_reg_esr_RNO_2Z0Z_19 ;
    wire \pid_front.N_55_0 ;
    wire \pid_front.N_110 ;
    wire \pid_front.error_i_regZ0Z_6 ;
    wire \pid_front.N_103_0 ;
    wire \pid_front.error_i_regZ0Z_7 ;
    wire \pid_front.error_i_regZ0Z_9 ;
    wire \pid_front.error_i_reg_esr_RNO_2Z0Z_25 ;
    wire \pid_front.error_i_reg_esr_RNO_1Z0Z_25_cascade_ ;
    wire \pid_front.N_93_0 ;
    wire \pid_front.error_i_reg_9_rn_1_25_cascade_ ;
    wire \pid_front.error_i_regZ0Z_25 ;
    wire \pid_front.N_29_1 ;
    wire \pid_front.N_32_0 ;
    wire \pid_front.error_i_regZ0Z_8 ;
    wire \pid_front.N_88_0_1 ;
    wire \pid_front.N_126_1 ;
    wire \pid_front.N_116_0 ;
    wire \pid_front.error_i_reg_9_rn_1_13_cascade_ ;
    wire \pid_front.N_127 ;
    wire \pid_front.error_i_regZ0Z_13 ;
    wire \pid_front.m1_0_03_cascade_ ;
    wire \pid_front.m1_2_03 ;
    wire pid_side_error_i_reg_9_sn_27;
    wire \pid_front.m61_0_bm_0 ;
    wire \pid_front.error_cry_3_0_c_RNI76FZ0Z08 ;
    wire \pid_front.error_i_regZ0Z_4 ;
    wire \pid_side.error_i_reg_9_sn_17 ;
    wire \pid_side.error_i_reg_9_sn_25 ;
    wire \ppm_encoder_1.aileronZ0Z_3 ;
    wire \ppm_encoder_1.pulses2countZ0Z_3 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_RNIUCMNZ0Z_1 ;
    wire \ppm_encoder_1.pulses2count_9_i_3_2 ;
    wire \ppm_encoder_1.aileronZ0Z_2 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_RNIC2521Z0Z_3 ;
    wire \ppm_encoder_1.pulses2countZ0Z_2 ;
    wire \ppm_encoder_1.N_295_i_0 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNIUTMRZ0 ;
    wire \ppm_encoder_1.pulses2count_9_0_0_1_3 ;
    wire \ppm_encoder_1.throttleZ0Z_3 ;
    wire \ppm_encoder_1.pulses2count_9_0_0_3_3 ;
    wire \ppm_encoder_1.counterZ0Z_14 ;
    wire \ppm_encoder_1.pulses2countZ0Z_14 ;
    wire \ppm_encoder_1.pulses2countZ0Z_15 ;
    wire \ppm_encoder_1.counterZ0Z_15 ;
    wire \ppm_encoder_1.counter24_0_I_45_c_RNOZ0 ;
    wire \ppm_encoder_1.counterZ0Z_16 ;
    wire \ppm_encoder_1.counterZ0Z_3 ;
    wire \ppm_encoder_1.counterZ0Z_17 ;
    wire \ppm_encoder_1.counterZ0Z_2 ;
    wire \ppm_encoder_1.un1_PPM_STATE_0_sqmuxa_0_i_a2_18_9 ;
    wire \pid_side.source_pid_1_sqmuxa_1_0_a4_4 ;
    wire \pid_side.un10lto12 ;
    wire \pid_side.error_i_acumm_preregZ0Z_21 ;
    wire \pid_side.error_i_acumm_preregZ0Z_13 ;
    wire \pid_side.error_i_acumm_preregZ0Z_22 ;
    wire \pid_side.error_i_acumm_preregZ0Z_23 ;
    wire \pid_side.error_i_acumm_preregZ0Z_24 ;
    wire \pid_side.error_i_acumm_preregZ0Z_17 ;
    wire \pid_side.error_i_acumm_preregZ0Z_5 ;
    wire \pid_side.un1_pid_prereg_0_17_cascade_ ;
    wire \pid_side.un1_pid_prereg_0_14 ;
    wire \pid_side.un1_pid_prereg_0_15 ;
    wire \pid_side.error_i_reg_esr_RNIQBRSZ0Z_24 ;
    wire \pid_side.un1_pid_prereg_0_17 ;
    wire \pid_side.un1_pid_prereg_0_18_cascade_ ;
    wire \pid_side.error_i_reg_esr_RNIO8QSZ0Z_23 ;
    wire \pid_side.un1_pid_prereg_0_16 ;
    wire \pid_side.un1_pid_prereg_0_19_cascade_ ;
    wire bfn_17_11_0_;
    wire \pid_side.pid_preregZ0Z_0 ;
    wire \pid_side.un1_pid_prereg_0_cry_0_c_THRU_CO ;
    wire \pid_side.pid_preregZ0Z_1 ;
    wire \pid_side.un1_pid_prereg_0_cry_0 ;
    wire \pid_side.pid_preregZ0Z_2 ;
    wire \pid_side.un1_pid_prereg_0_cry_1 ;
    wire \pid_side.pid_preregZ0Z_3 ;
    wire \pid_side.un1_pid_prereg_0_cry_2 ;
    wire \pid_side.pid_preregZ0Z_4 ;
    wire \pid_side.un1_pid_prereg_0_cry_3 ;
    wire \pid_side.pid_preregZ0Z_5 ;
    wire \pid_side.un1_pid_prereg_0_cry_4 ;
    wire \pid_side.un1_pid_prereg_0_cry_5 ;
    wire \pid_side.un1_pid_prereg_0_cry_6 ;
    wire \pid_side.error_p_reg_esr_RNIODMH3_0Z0Z_6 ;
    wire bfn_17_12_0_;
    wire \pid_side.error_p_reg_esr_RNIKF8V6Z0Z_7 ;
    wire \pid_side.error_p_reg_esr_RNIODMH3Z0Z_6 ;
    wire \pid_side.un1_pid_prereg_0_cry_7 ;
    wire \pid_side.error_p_reg_esr_RNIECBV6Z0Z_8 ;
    wire \pid_side.error_p_reg_esr_RNIS1ID3Z0Z_7 ;
    wire \pid_side.un1_pid_prereg_0_cry_8 ;
    wire \pid_side.un1_pid_prereg_0_cry_9 ;
    wire \pid_side.un1_pid_prereg_0_cry_10 ;
    wire \pid_side.error_d_reg_prev_esr_RNITU3P4Z0Z_10 ;
    wire \pid_side.pid_preregZ0Z_12 ;
    wire \pid_side.un1_pid_prereg_0_cry_11 ;
    wire \pid_side.un1_pid_prereg_0_cry_12 ;
    wire \pid_side.un1_pid_prereg_0_cry_13_THRU_CO ;
    wire \pid_side.un1_pid_prereg_0_cry_13 ;
    wire \pid_side.un1_pid_prereg_0_cry_14 ;
    wire bfn_17_13_0_;
    wire \pid_side.un1_pid_prereg_0_cry_15 ;
    wire \pid_side.un1_pid_prereg_0_cry_16 ;
    wire \pid_side.un1_pid_prereg_0_cry_17 ;
    wire \pid_side.un1_pid_prereg_0_cry_18 ;
    wire \pid_side.pid_preregZ0Z_20 ;
    wire \pid_side.un1_pid_prereg_0_cry_19 ;
    wire \pid_side.pid_preregZ0Z_21 ;
    wire \pid_side.un1_pid_prereg_0_cry_20 ;
    wire \pid_side.pid_preregZ0Z_22 ;
    wire \pid_side.un1_pid_prereg_0_cry_21 ;
    wire \pid_side.un1_pid_prereg_0_cry_22 ;
    wire \pid_side.error_d_reg_prev_esr_RNIK1TV8Z0Z_22 ;
    wire \pid_side.pid_preregZ0Z_23 ;
    wire bfn_17_14_0_;
    wire \pid_side.error_d_reg_prev_esr_RNIFQK34Z0Z_22 ;
    wire \pid_side.error_d_reg_prev_esr_RNI33ME7Z0Z_22 ;
    wire \pid_side.pid_preregZ0Z_24 ;
    wire \pid_side.un1_pid_prereg_0_cry_23 ;
    wire \pid_side.error_d_reg_prev_esr_RNICN4M6Z0Z_22 ;
    wire \pid_side.error_d_reg_prev_esr_RNIK81B3Z0Z_22 ;
    wire \pid_side.pid_preregZ0Z_25 ;
    wire \pid_side.un1_pid_prereg_0_cry_24 ;
    wire \pid_side.error_d_reg_prev_esr_RNIOE3B3Z0Z_22 ;
    wire \pid_side.pid_preregZ0Z_26 ;
    wire \pid_side.un1_pid_prereg_0_cry_25 ;
    wire \pid_side.error_d_reg_prev_esr_RNISFDM6Z0Z_22 ;
    wire \pid_side.pid_preregZ0Z_27 ;
    wire \pid_side.un1_pid_prereg_0_cry_26 ;
    wire \pid_side.error_d_reg_prev_esr_RNI3RHM6Z0Z_22 ;
    wire \pid_side.error_d_reg_prev_esr_RNI0R7B3Z0Z_22 ;
    wire \pid_side.pid_preregZ0Z_28 ;
    wire \pid_side.un1_pid_prereg_0_cry_27 ;
    wire \pid_side.error_d_reg_prev_esr_RNI72LM6Z0Z_22 ;
    wire \pid_side.error_d_reg_prev_esr_RNI30AB3Z0Z_22 ;
    wire \pid_side.pid_preregZ0Z_29 ;
    wire \pid_side.un1_pid_prereg_0_cry_28 ;
    wire \pid_side.un1_pid_prereg_0_axb_30 ;
    wire \pid_side.un1_pid_prereg_0_cry_29 ;
    wire \pid_side.pid_preregZ0Z_30 ;
    wire \pid_side.N_838_g ;
    wire \pid_side.un1_pid_prereg_370_1 ;
    wire \pid_side.error_i_reg_esr_RNIM5PSZ0Z_22 ;
    wire \pid_side.un1_pid_prereg_0_1_cascade_ ;
    wire \pid_side.error_d_reg_prev_esr_RNIMFTP4Z0Z_14 ;
    wire \pid_side.error_i_reg_esr_RNISCPRZ0Z_16 ;
    wire \pid_side.un1_pid_prereg_0_2_cascade_ ;
    wire \pid_side.error_d_reg_prev_esr_RNISHTJ9Z0Z_14 ;
    wire \pid_side.error_d_reg_prev_esr_RNISM2K9Z0Z_15 ;
    wire \pid_side.un1_pid_prereg_0_5_cascade_ ;
    wire \pid_side.error_d_reg_prev_esr_RNIMK2Q4Z0Z_16 ;
    wire \pid_side.error_i_reg_esr_RNI0JRRZ0Z_18 ;
    wire \pid_side.un1_pid_prereg_0_5 ;
    wire \pid_side.un1_pid_prereg_0_6_cascade_ ;
    wire \pid_side.error_d_reg_prev_esr_RNISR7K9Z0Z_16 ;
    wire \pid_side.un1_pid_prereg_0_7_cascade_ ;
    wire \pid_side.error_d_reg_prev_esr_RNI675Q4Z0Z_17 ;
    wire \pid_side.error_i_reg_esr_RNIUFQRZ0Z_17 ;
    wire \pid_side.un1_pid_prereg_0_4 ;
    wire \pid_side.m21_ns_1 ;
    wire \pid_side.g0_i_m4_1_cascade_ ;
    wire \pid_side.N_8_0 ;
    wire \pid_side.N_36_0_cascade_ ;
    wire \pid_side.error_i_reg_esr_RNO_2Z0Z_16 ;
    wire \pid_side.N_36_0 ;
    wire \pid_side.N_57_0_cascade_ ;
    wire \pid_side.N_59_0_cascade_ ;
    wire \pid_side.N_89_i ;
    wire \pid_side.error_i_regZ0Z_24 ;
    wire \pid_front.error_p_regZ0Z_18 ;
    wire \pid_front.error_p_reg_esr_RNITCC61Z0Z_18 ;
    wire \pid_front.error_d_reg_prevZ0Z_18 ;
    wire \pid_front.N_764_0 ;
    wire \pid_front.N_1705_g ;
    wire drone_H_disp_side_11;
    wire \pid_side.N_9_1 ;
    wire \pid_side.m87_0_ns_1_cascade_ ;
    wire \pid_side.N_88_0_cascade_ ;
    wire \pid_side.N_90_0 ;
    wire \pid_side.N_48_1 ;
    wire \pid_side.N_48_1_cascade_ ;
    wire \pid_side.N_89_0 ;
    wire \pid_side.N_126 ;
    wire \pid_side.N_88_0 ;
    wire \pid_side.error_i_reg_9_sn_13 ;
    wire \pid_side.N_127_cascade_ ;
    wire \pid_side.error_i_regZ0Z_13 ;
    wire xy_ki_6;
    wire xy_ki_5;
    wire xy_ki_7;
    wire pid_side_m153_e_4;
    wire \pid_side.m1_0_03 ;
    wire \pid_side.N_89_0_1_cascade_ ;
    wire \pid_side.error_i_reg_9_rn_2_13 ;
    wire pid_side_N_166_mux_cascade_;
    wire pid_front_error_i_reg_9_rn_sn_15;
    wire pid_front_error_i_reg_9_rn_sn_15_cascade_;
    wire \pid_front.m1_0_03 ;
    wire pid_side_N_166_mux;
    wire \pid_front.N_12_1 ;
    wire \pid_front.error_i_regZ0Z_1 ;
    wire \pid_side.m1_2_03 ;
    wire \pid_side.error_i_reg_9_rn_rn_2_13 ;
    wire \pid_front.error_i_reg_esr_RNO_1Z0Z_15 ;
    wire \pid_front.error_i_reg_esr_RNO_2Z0Z_15 ;
    wire \pid_front.error_i_regZ0Z_15 ;
    wire \pid_front.N_134 ;
    wire xy_ki_2;
    wire \pid_front.error_i_reg_esr_RNO_0_0_23_cascade_ ;
    wire \pid_front.error_i_regZ0Z_23 ;
    wire \pid_front.error_cry_9_c_RNICELJ1Z0Z_0_cascade_ ;
    wire \pid_front.error_cry_9_c_RNICELJZ0Z1 ;
    wire \pid_front.N_46_1 ;
    wire pid_front_error_i_reg_9_sn_19;
    wire \pid_front.N_46_1_cascade_ ;
    wire \pid_front.error_i_reg_esr_RNO_1Z0Z_19 ;
    wire \pid_front.O_5 ;
    wire \pid_front.error_d_regZ0Z_3 ;
    wire \pid_front.error_15 ;
    wire \pid_front.N_131_cascade_ ;
    wire \pid_front.m5_2_03 ;
    wire \pid_front.error_i_reg_9_sn_17 ;
    wire \pid_front.error_i_reg_9_rn_1_17_cascade_ ;
    wire \pid_front.error_i_regZ0Z_17 ;
    wire \pid_front.state_ns_0_0 ;
    wire \pid_front.error_i_reg_esr_RNO_4_0_17 ;
    wire \pid_front.N_51_1 ;
    wire \pid_front.N_48_1 ;
    wire \pid_front.N_47_1 ;
    wire \pid_front.m89_0_ns_1_cascade_ ;
    wire \pid_front.N_45_1 ;
    wire \pid_front.N_90_0 ;
    wire \pid_front.error_14 ;
    wire xy_ki_1;
    wire \pid_front.error_i_reg_esr_RNO_5_0_17 ;
    wire \pid_alt.state_RNIFCSD1Z0Z_0 ;
    wire \pid_alt.N_939_0 ;
    wire \pid_side.pid_preregZ0Z_10 ;
    wire \pid_side.pid_preregZ0Z_7 ;
    wire \pid_side.pid_preregZ0Z_11 ;
    wire \pid_side.pid_preregZ0Z_6 ;
    wire \pid_side.pid_preregZ0Z_13 ;
    wire \pid_side.pid_preregZ0Z_9 ;
    wire \pid_side.source_pid_1_sqmuxa_1_0_a2_1_4_cascade_ ;
    wire \pid_side.pid_preregZ0Z_8 ;
    wire \pid_side.N_99 ;
    wire \pid_side.pid_preregZ0Z_17 ;
    wire \pid_side.pid_preregZ0Z_18 ;
    wire \pid_side.pid_preregZ0Z_19 ;
    wire \pid_side.pid_preregZ0Z_16 ;
    wire \pid_side.un11lto30_i_a2_3_and ;
    wire \pid_side.pid_preregZ0Z_15 ;
    wire \pid_side.un11lto30_i_a2_3_and_cascade_ ;
    wire \pid_side.pid_preregZ0Z_14 ;
    wire \pid_side.source_pid_1_sqmuxa_1_0_a2_0_0 ;
    wire \pid_side.stateZ0Z_1 ;
    wire \pid_side.error_i_acumm_preregZ0Z_28 ;
    wire \pid_side.error_i_acumm_3_sqmuxa ;
    wire \pid_side.error_p_reg_esr_RNI5RKP3Z0Z_5 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_0_c_RNITGKN ;
    wire \pid_side.error_d_reg_prev_esr_RNIM6H42Z0Z_0 ;
    wire \pid_side.N_2380_i ;
    wire \pid_side.error_p_reg_esr_RNIIAPH3Z0Z_8 ;
    wire \pid_side.error_p_reg_esr_RNIKGHS6Z0Z_10 ;
    wire \pid_side.N_2386_i_cascade_ ;
    wire \pid_side.error_p_reg_esr_RNIRE1B1Z0Z_10 ;
    wire \pid_side.error_d_reg_prev_esr_RNITU3P4_0Z0Z_10 ;
    wire \pid_side.error_p_reg_esr_RNI1VTC1Z0Z_9 ;
    wire \pid_side.error_p_reg_esr_RNIRE1B1Z0Z_10_cascade_ ;
    wire \pid_side.error_i_reg_esr_RNI6OOIZ0Z_10 ;
    wire \pid_side.error_p_reg_esr_RNIV4S38Z0Z_10 ;
    wire \pid_side.error_i_reg_esr_RNISESSZ0Z_25 ;
    wire \pid_side.un1_pid_prereg_0_18 ;
    wire \pid_side.un1_pid_prereg_0_19 ;
    wire \pid_side.un1_pid_prereg_0_20_cascade_ ;
    wire \pid_side.error_d_reg_prev_esr_RNIK39M6Z0Z_22 ;
    wire \pid_side.error_i_reg_esr_RNIUHTSZ0Z_26 ;
    wire \pid_side.un1_pid_prereg_0_21 ;
    wire \pid_side.un1_pid_prereg_0_21_cascade_ ;
    wire \pid_side.un1_pid_prereg_0_20 ;
    wire \pid_side.error_d_reg_prev_esr_RNISK5B3Z0Z_22 ;
    wire \pid_side.error_d_reg_prevZ0Z_22 ;
    wire \pid_side.error_d_reg_prevZ0Z_21 ;
    wire \pid_side.error_d_reg_prev_esr_RNIVNLOZ0Z_21 ;
    wire \pid_side.error_d_reg_prev_esr_RNICOLL9Z0Z_18 ;
    wire \pid_side.un1_pid_prereg_0_10_cascade_ ;
    wire \pid_side.error_d_reg_prev_esr_RNIQVAR4Z0Z_19 ;
    wire \pid_side.error_d_reg_prev_esr_RNIVNLO_0Z0Z_21 ;
    wire \pid_side.error_i_reg_esr_RNIK2OSZ0Z_21 ;
    wire \pid_side.un1_pid_prereg_0_11 ;
    wire \pid_side.un1_pid_prereg_0_10 ;
    wire \pid_side.un1_pid_prereg_0_12_cascade_ ;
    wire \pid_side.error_d_reg_prev_esr_RNIV6JN9Z0Z_19 ;
    wire \pid_side.un1_pid_prereg_0_2 ;
    wire \pid_side.un1_pid_prereg_0_3 ;
    wire \pid_side.error_d_reg_prev_esr_RNI620Q4Z0Z_15 ;
    wire \pid_side.un1_pid_prereg_0_12 ;
    wire \pid_side.un1_pid_prereg_0_13 ;
    wire \pid_side.error_d_reg_prev_esr_RNI578S4Z0Z_20 ;
    wire \pid_side.un1_pid_prereg_0_1 ;
    wire \pid_side.un1_pid_prereg_0_0 ;
    wire \pid_side.error_d_reg_prev_esr_RNI1OK5FZ0Z_12 ;
    wire \pid_side.error_i_reg_esr_RNI2MSRZ0Z_19 ;
    wire \pid_side.un1_pid_prereg_0_7 ;
    wire \pid_side.un1_pid_prereg_0_6 ;
    wire \pid_side.un1_pid_prereg_0_8_cascade_ ;
    wire \pid_side.error_d_reg_prev_esr_RNIOVFK9Z0Z_17 ;
    wire \pid_side.error_i_reg_esr_RNIRGURZ0Z_20 ;
    wire \pid_side.un1_pid_prereg_0_9 ;
    wire \pid_side.un1_pid_prereg_0_9_cascade_ ;
    wire \pid_side.un1_pid_prereg_0_8 ;
    wire \pid_side.error_d_reg_prev_esr_RNIIOAQ4Z0Z_18 ;
    wire \pid_side.un1_pid_prereg_0 ;
    wire \pid_side.error_d_reg_prev_esr_RNIQ8P41Z0Z_0 ;
    wire uart_pc_data_6;
    wire side_command_7;
    wire \Commands_frame_decoder.source_CH2data_1_sqmuxa_0 ;
    wire dron_frame_decoder_1_source_H_disp_side_fast_0;
    wire \pid_side.error_axb_0 ;
    wire bfn_18_17_0_;
    wire \pid_side.error_axbZ0Z_1 ;
    wire \pid_side.error_1 ;
    wire \pid_side.error_cry_0 ;
    wire \pid_side.error_axbZ0Z_2 ;
    wire \pid_side.error_cry_1 ;
    wire \pid_side.error_axbZ0Z_3 ;
    wire \pid_side.error_cry_2 ;
    wire drone_H_disp_side_i_4;
    wire side_command_0;
    wire \pid_side.error_cry_3 ;
    wire drone_H_disp_side_i_5;
    wire side_command_1;
    wire \pid_side.error_cry_0_0 ;
    wire side_command_2;
    wire drone_H_disp_side_i_6;
    wire \pid_side.error_cry_1_0 ;
    wire side_command_3;
    wire drone_H_disp_side_i_7;
    wire \pid_side.error_cry_2_0 ;
    wire \pid_side.error_cry_3_0 ;
    wire drone_H_disp_side_i_8;
    wire side_command_4;
    wire bfn_18_18_0_;
    wire drone_H_disp_side_i_9;
    wire side_command_5;
    wire \pid_side.error_cry_4 ;
    wire drone_H_disp_side_i_10;
    wire side_command_6;
    wire \pid_side.error_cry_5 ;
    wire \pid_side.error_axbZ0Z_7 ;
    wire \pid_side.error_11 ;
    wire \pid_side.error_cry_6 ;
    wire \pid_side.error_axb_8_l_ofxZ0 ;
    wire drone_H_disp_side_12;
    wire \pid_side.error_12 ;
    wire \pid_side.error_cry_7 ;
    wire drone_H_disp_side_i_12;
    wire drone_H_disp_side_13;
    wire \pid_side.error_cry_8 ;
    wire drone_H_disp_side_i_13;
    wire \pid_side.error_cry_9 ;
    wire drone_H_disp_side_15;
    wire drone_H_disp_side_14;
    wire \pid_side.error_cry_10 ;
    wire \pid_side.error_15 ;
    wire \pid_side.error_8 ;
    wire \pid_side.N_48_1_0_cascade_ ;
    wire \pid_side.N_51_1_0 ;
    wire \pid_side.N_48_1_0 ;
    wire \pid_side.error_i_reg_esr_RNO_9Z0Z_21_cascade_ ;
    wire \pid_side.error_i_reg_esr_RNO_10Z0Z_21 ;
    wire \pid_side.N_116_0_0 ;
    wire \pid_side.N_51_1 ;
    wire \pid_side.error_9 ;
    wire \pid_side.error_10 ;
    wire \pid_side.error_13 ;
    wire \pid_side.G_5_0_m4_1_cascade_ ;
    wire \pid_side.error_14 ;
    wire \pid_side.N_7 ;
    wire \pid_side.error_6 ;
    wire \pid_side.error_7 ;
    wire \pid_side.g0_7_1 ;
    wire xy_ki_3;
    wire \pid_side.N_117 ;
    wire pid_side_N_166;
    wire \pid_side.error_i_regZ0Z_5 ;
    wire \pid_side.state_ns_0_0 ;
    wire \pid_side.g0_6_1_cascade_ ;
    wire \pid_side.N_12_1_1 ;
    wire \pid_side.N_12_1_1_cascade_ ;
    wire \pid_side.N_89_0_1 ;
    wire \pid_side.N_116_0 ;
    wire \pid_side.error_3 ;
    wire \pid_side.error_2 ;
    wire \pid_side.error_5 ;
    wire \pid_side.error_4 ;
    wire \pid_side.g0_10_1_cascade_ ;
    wire \pid_side.N_12_1_0 ;
    wire drone_H_disp_front_0;
    wire \pid_front.error_1 ;
    wire \pid_front.error_2 ;
    wire \pid_front.m14_0_ns_1_cascade_ ;
    wire \pid_front.error_3 ;
    wire \pid_front.N_15_1_cascade_ ;
    wire xy_ki_4;
    wire pid_front_N_331;
    wire \pid_front.m3_2_03_cascade_ ;
    wire \pid_front.error_i_reg_9_rn_rn_2_15 ;
    wire \pid_front.N_15_1 ;
    wire \pid_front.N_104 ;
    wire xy_ki_3_rep2;
    wire \pid_front.N_104_cascade_ ;
    wire \pid_front.N_39_0 ;
    wire \pid_front.N_49_0 ;
    wire \pid_front.error_i_reg_esr_RNO_2Z0Z_23_cascade_ ;
    wire \pid_front.error_i_reg_esr_RNO_3Z0Z_23 ;
    wire \pid_front.error_i_reg_esr_RNO_1_0_23 ;
    wire xy_ki_0_rep1;
    wire xy_ki_0_rep2;
    wire xy_ki_fast_0;
    wire xy_ki_1_rep1;
    wire xy_ki_fast_1;
    wire xy_ki_2_rep1;
    wire uart_pc_data_2;
    wire xy_ki_fast_2;
    wire \pid_side.O_2_9 ;
    wire \pid_side.error_p_reg_esr_RNI76TK1_0Z0Z_5_cascade_ ;
    wire \pid_side.error_p_reg_esr_RNIG7MC2Z0Z_5 ;
    wire \pid_side.error_p_reg_esr_RNIIHEQZ0Z_4 ;
    wire \pid_side.error_p_reg_esr_RNIIHEQZ0Z_4_cascade_ ;
    wire \pid_side.error_d_reg_prevZ0Z_5 ;
    wire \pid_side.error_p_regZ0Z_6 ;
    wire \pid_side.N_2362_i ;
    wire \pid_side.error_p_reg_esr_RNIIFTC1_0Z0Z_6 ;
    wire \pid_side.error_p_reg_esr_RNIIFTC1_0Z0Z_6_cascade_ ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_5_c_RNIC5QN ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_4_c_RNI91PN ;
    wire \pid_side.error_p_reg_esr_RNI76TK1_0Z0Z_5 ;
    wire \pid_side.un1_pid_prereg_66_0_cascade_ ;
    wire \pid_side.error_p_reg_esr_RNI76TK1Z0Z_5 ;
    wire \pid_side.error_p_reg_esr_RNIL2B66Z0Z_5 ;
    wire \pid_side.error_d_reg_prevZ0Z_9 ;
    wire \pid_side.error_p_reg_esr_RNI4O091_0Z0Z_10_cascade_ ;
    wire \pid_side.error_p_reg_esr_RNI4O091Z0Z_10 ;
    wire \pid_side.error_d_reg_prev_esr_RNIV62K2Z0Z_10_cascade_ ;
    wire \pid_side.error_d_reg_prev_esr_RNID3GT3_0Z0Z_10 ;
    wire \pid_side.error_i_reg_esr_RNIGRJRZ0Z_11 ;
    wire \pid_side.un1_pid_prereg_153_0_cascade_ ;
    wire \pid_side.error_d_reg_prev_esr_RNII28CBZ0Z_10 ;
    wire \pid_side.error_d_reg_prevZ0Z_10 ;
    wire \pid_side.error_d_reg_prev_esr_RNIV62K2Z0Z_10 ;
    wire \pid_side.error_d_reg_prev_esr_RNID3GT3Z0Z_10 ;
    wire \pid_side.error_i_reg_esr_RNIJVKRZ0Z_12 ;
    wire \pid_side.error_d_reg_prev_esr_RNISSNM4Z0Z_12 ;
    wire \pid_side.error_d_reg_prev_esr_RNID3GT3Z0Z_10_cascade_ ;
    wire \pid_side.error_d_reg_prev_esr_RNIH0S9BZ0Z_10 ;
    wire \pid_side.O_1_6 ;
    wire \Commands_frame_decoder.source_xy_ki_1_sqmuxa_0 ;
    wire reset_system_g;
    wire \pid_side.error_d_reg_prev_esr_RNI5RIOZ0Z_14 ;
    wire \pid_side.error_d_reg_prev_esr_RNI5RIOZ0Z_14_cascade_ ;
    wire \pid_side.error_i_reg_esr_RNIQ9ORZ0Z_15 ;
    wire \pid_side.error_d_reg_prev_esr_RNI8UIO_0Z0Z_15 ;
    wire \pid_side.error_d_reg_prevZ0Z_15 ;
    wire \pid_side.error_d_reg_prev_esr_RNI8UIOZ0Z_15 ;
    wire \pid_side.error_d_reg_prev_esr_RNIB8NBAZ0Z_12 ;
    wire \pid_side.error_d_reg_prev_esr_RNI73UC2_0Z0Z_14 ;
    wire \pid_side.error_d_reg_prev_esr_RNI0UI8JZ0Z_12 ;
    wire \pid_side.error_d_reg_prev_esr_RNI5RIO_0Z0Z_14 ;
    wire \pid_side.un1_pid_prereg_97_cascade_ ;
    wire \pid_side.error_d_reg_prev_esr_RNI45PU7Z0Z_12 ;
    wire \pid_side.error_d_reg_fast_esr_RNIPHKNZ0Z_12 ;
    wire \pid_side.error_d_reg_fast_esr_RNIPEC11Z0Z_12 ;
    wire \pid_side.error_d_reg_fast_esr_RNIEIJH2Z0Z_12_cascade_ ;
    wire \pid_side.g1_2_1_cascade_ ;
    wire \pid_side.g1_3_cascade_ ;
    wire \pid_side.error_p_reg_esr_RNILLRS8Z0Z_12 ;
    wire \pid_side.N_2405_0_0_0_cascade_ ;
    wire \pid_side.g0_2_0_cascade_ ;
    wire \pid_side.error_d_reg_prev_esr_RNIQ0PB4Z0Z_12 ;
    wire \pid_side.N_4_1_0_1 ;
    wire drone_H_disp_side_0;
    wire xy_ki_1_rep2;
    wire xy_ki_0;
    wire xy_ki_2_rep2;
    wire xy_ki_3_rep1;
    wire \pid_side.m0_0_03 ;
    wire \pid_side.m0_2_03 ;
    wire \pid_side.O_2_7 ;
    wire \pid_side.O_2_12 ;
    wire \pid_side.error_p_regZ0Z_9 ;
    wire \pid_side.O_2_8 ;
    wire \pid_side.error_p_regZ0Z_5 ;
    wire \pid_side.O_1_7 ;
    wire \pid_side.error_d_regZ0Z_5 ;
    wire \pid_side.O_2_6 ;
    wire \pid_side.O_1_4 ;
    wire \pid_side.O_1_12 ;
    wire \pid_side.error_d_regZ0Z_10 ;
    wire \pid_side.O_1_8 ;
    wire \pid_side.error_d_regZ0Z_6 ;
    wire \pid_side.O_1_9 ;
    wire \pid_side.error_d_regZ0Z_7 ;
    wire \pid_side.O_1_10 ;
    wire \pid_side.error_d_regZ0Z_8 ;
    wire \pid_side.O_1_11 ;
    wire \pid_side.error_d_regZ0Z_9 ;
    wire \pid_side.O_2_4 ;
    wire \pid_side.O_2_13 ;
    wire \pid_side.error_p_regZ0Z_10 ;
    wire \pid_side.error_p_reg_esr_RNIG7MC2_0Z0Z_5 ;
    wire \pid_side.error_p_reg_esr_RNIFEEQZ0Z_3_cascade_ ;
    wire \pid_side.error_p_reg_esr_RNIN4BP4Z0Z_3 ;
    wire \pid_side.error_p_regZ0Z_4 ;
    wire \pid_side.error_d_reg_prevZ0Z_4 ;
    wire \pid_side.error_d_regZ0Z_4 ;
    wire \pid_side.error_p_reg_esr_RNIIHEQ_0Z0Z_4 ;
    wire \pid_side.error_p_reg_esr_RNIFEEQZ0Z_3 ;
    wire \pid_side.error_p_reg_esr_RNIIHEQ_0Z0Z_4_cascade_ ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_3_c_RNI6TNN ;
    wire \pid_side.error_p_reg_esr_RNI5G8P4Z0Z_3 ;
    wire \pid_side.error_p_reg_esr_RNIUIJC2Z0Z_2 ;
    wire \pid_side.error_d_reg_prevZ0Z_3 ;
    wire \pid_side.error_p_regZ0Z_3 ;
    wire \pid_side.error_p_reg_esr_RNIFEEQ_0Z0Z_3 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_2_c_RNI3PMN ;
    wire \pid_side.error_p_reg_esr_RNIFEEQ_0Z0Z_3_cascade_ ;
    wire \pid_side.error_p_reg_esr_RNI7U286Z0Z_2 ;
    wire \pid_side.error_d_reg_prev_esr_RNIKAJO_0Z0Z_19 ;
    wire \pid_side.error_d_reg_prevZ0Z_19 ;
    wire \pid_side.error_d_reg_prev_esr_RNIKAJOZ0Z_19 ;
    wire \pid_side.g0_1_0 ;
    wire \pid_side.error_d_reg_prev_esr_RNISHIO_1Z0Z_11 ;
    wire \pid_side.error_d_reg_prev_esr_RNISKLO_0Z0Z_20 ;
    wire \pid_side.N_2398_i_cascade_ ;
    wire \pid_side.error_p_reg_esr_RNIL0VP1Z0Z_12 ;
    wire \pid_side.error_d_reg_prevZ0Z_11 ;
    wire \pid_side.N_2398_i ;
    wire \pid_side.un1_pid_prereg_79_cascade_ ;
    wire \pid_side.un1_pid_prereg_167_0_1_cascade_ ;
    wire \pid_side.un1_pid_prereg_167_0 ;
    wire \pid_side.g0_19_1_1 ;
    wire \pid_side.g0_19_1 ;
    wire \pid_side.un1_pid_prereg_135_0 ;
    wire \pid_side.N_3_i_1_1_cascade_ ;
    wire \pid_side.un1_pid_prereg_79 ;
    wire \pid_side.N_5_0 ;
    wire \pid_side.N_3_i_1_cascade_ ;
    wire \pid_side.error_i_reg_esr_RNIO6NRZ0Z_14 ;
    wire \pid_side.error_i_reg_esr_RNIM3MRZ0Z_13 ;
    wire \pid_side.error_d_reg_prev_esr_RNIQTGL4Z0Z_12_cascade_ ;
    wire \pid_side.error_d_reg_prev_esr_RNI6P1R3Z0Z_12 ;
    wire \pid_side.un1_pid_prereg_0_axb_14 ;
    wire \pid_side.error_d_reg_prev_fastZ0Z_12 ;
    wire \pid_side.g1_1_cascade_ ;
    wire \pid_side.g0_3_2 ;
    wire \pid_side.error_d_reg_fastZ0Z_12 ;
    wire \pid_side.N_5_1 ;
    wire \pid_side.error_d_reg_prevZ0Z_12 ;
    wire \pid_side.error_d_reg_fast_esr_RNIEIJH2Z0Z_12 ;
    wire \pid_side.error_d_reg_prev_esr_RNI41F23Z0Z_12 ;
    wire \pid_side.error_d_reg_prev_esr_RNI9BFR3Z0Z_1 ;
    wire \pid_side.error_p_reg_esr_RNIIQL11_0Z0Z_1_cascade_ ;
    wire \pid_side.error_d_reg_prev_esr_RNIBGIE2Z0Z_1 ;
    wire \pid_side.un1_error_i_acumm_prereg_cry_1_c_RNI0LLN ;
    wire \pid_side.error_d_reg_prev_esr_RNIBGIE2Z0Z_1_cascade_ ;
    wire \pid_side.error_d_reg_prev_esr_RNI905J4Z0Z_1 ;
    wire \pid_side.error_p_reg_esr_RNIIQL11Z0Z_1 ;
    wire \pid_side.error_d_reg_prev_esr_RNIIFEIZ0Z_1 ;
    wire \pid_side.error_d_reg_prevZ0Z_0 ;
    wire \pid_side.error_p_reg_esr_RNICBEQ_0Z0Z_2 ;
    wire \pid_side.O_0_2 ;
    wire \pid_side.error_d_regZ0Z_0 ;
    wire \pid_side.O_1_5 ;
    wire \pid_side.error_d_regZ0Z_3 ;
    wire \pid_side.O_2_5 ;
    wire \pid_side.error_d_reg_prevZ0Z_1 ;
    wire \pid_side.error_p_regZ0Z_1 ;
    wire \pid_side.un1_pid_prereg_9_0 ;
    wire \pid_side.error_d_regZ0Z_2 ;
    wire \pid_side.error_p_regZ0Z_2 ;
    wire \pid_side.error_d_reg_prevZ0Z_2 ;
    wire \pid_side.error_p_reg_esr_RNICBEQZ0Z_2 ;
    wire \pid_side.state_RNINK4UZ0Z_0 ;
    wire \pid_side.O_2_14 ;
    wire \pid_side.error_p_regZ0Z_11 ;
    wire \pid_side.O_1_17 ;
    wire \pid_side.error_d_regZ0Z_15 ;
    wire \pid_side.O_1_13 ;
    wire \pid_side.error_d_regZ0Z_11 ;
    wire \pid_side.O_1_14 ;
    wire \pid_side.error_d_regZ0Z_12 ;
    wire \pid_front.O_16 ;
    wire \pid_front.error_d_regZ0Z_14 ;
    wire xy_kp_1;
    wire \Commands_frame_decoder.state_RNIG48SZ0Z_7 ;
    wire \pid_side.error_d_reg_prev_esr_RNIB1JOZ0Z_16 ;
    wire \pid_side.error_d_reg_prev_esr_RNIE4JO_0Z0Z_17 ;
    wire \pid_side.error_d_reg_prevZ0Z_17 ;
    wire \pid_side.error_d_reg_prev_esr_RNIE4JOZ0Z_17 ;
    wire \pid_side.error_d_reg_prev_esr_RNIH7JO_0Z0Z_18 ;
    wire \pid_side.N_838_0 ;
    wire \pid_side.state_RNIIIOOZ0Z_0 ;
    wire \pid_side.error_d_reg_prevZ0Z_18 ;
    wire \pid_side.error_d_reg_prev_esr_RNIH7JOZ0Z_18 ;
    wire \pid_side.O_1_3 ;
    wire \pid_side.error_d_regZ0Z_1 ;
    wire \pid_side.error_d_reg_prev_esr_RNI2OIO_4Z0Z_13 ;
    wire \pid_side.error_d_reg_prevZ0Z_20 ;
    wire \pid_side.error_d_reg_prev_esr_RNISKLOZ0Z_20 ;
    wire \pid_side.error_d_reg_prevZ0Z_16 ;
    wire \pid_side.error_d_reg_prev_esr_RNIB1JO_0Z0Z_16 ;
    wire \pid_side.error_d_reg_prevZ0Z_14 ;
    wire \pid_side.N_2405_0_cascade_ ;
    wire \pid_side.g0_2 ;
    wire uart_pc_data_1;
    wire xy_kd_1;
    wire uart_pc_data_3;
    wire xy_kd_3;
    wire uart_pc_data_0;
    wire xy_kd_0;
    wire \pid_front.O_22 ;
    wire \pid_front.error_d_regZ0Z_20 ;
    wire \pid_side.O_2_22 ;
    wire \pid_side.error_p_regZ0Z_19 ;
    wire \pid_side.O_2_24 ;
    wire \pid_side.error_p_regZ0Z_21 ;
    wire \pid_side.O_2_21 ;
    wire \pid_side.error_p_regZ0Z_18 ;
    wire \pid_side.O_2_17 ;
    wire \pid_side.error_p_regZ0Z_14 ;
    wire \pid_side.O_2_10 ;
    wire \pid_side.error_p_regZ0Z_7 ;
    wire \pid_side.O_2_11 ;
    wire \pid_side.error_p_regZ0Z_8 ;
    wire \pid_side.O_2_16 ;
    wire \pid_side.O_2_20 ;
    wire \pid_side.error_p_regZ0Z_17 ;
    wire \pid_side.O_2_18 ;
    wire \pid_side.error_p_regZ0Z_15 ;
    wire \pid_side.O_2_19 ;
    wire \pid_side.error_p_regZ0Z_16 ;
    wire \pid_side.O_2_23 ;
    wire \pid_side.error_p_regZ0Z_20 ;
    wire \pid_side.O_2_15 ;
    wire \pid_side.error_p_regZ0Z_12 ;
    wire \pid_side.O_1_19 ;
    wire \pid_side.error_d_regZ0Z_17 ;
    wire \pid_side.O_1_20 ;
    wire \pid_side.error_d_regZ0Z_18 ;
    wire \pid_side.O_1_21 ;
    wire \pid_side.error_d_regZ0Z_19 ;
    wire \pid_side.O_1_23 ;
    wire \pid_side.error_d_regZ0Z_21 ;
    wire \pid_side.O_1_24 ;
    wire \pid_side.error_d_regZ0Z_22 ;
    wire \pid_side.O_1_22 ;
    wire \pid_side.error_d_regZ0Z_20 ;
    wire \pid_side.O_2_3 ;
    wire \pid_side.error_p_regZ0Z_0 ;
    wire \pid_side.O_1_15 ;
    wire \pid_side.O_1_16 ;
    wire \pid_side.error_d_regZ0Z_14 ;
    wire \pid_side.O_1_18 ;
    wire \pid_side.error_d_regZ0Z_16 ;
    wire \pid_side.N_873_0 ;
    wire \pid_side.N_5 ;
    wire \pid_side.error_d_regZ0Z_13 ;
    wire \pid_side.error_d_reg_prevZ0Z_13 ;
    wire \pid_side.error_p_regZ0Z_13 ;
    wire \pid_side.error_d_reg_prev_esr_RNI2OIO_1Z0Z_13 ;
    wire \pid_front.O_4 ;
    wire \pid_front.error_d_regZ0Z_2 ;
    wire uart_pc_data_7;
    wire xy_kd_7;
    wire uart_pc_data_5;
    wire xy_kd_5;
    wire uart_pc_data_4;
    wire xy_kd_4;
    wire \Commands_frame_decoder.state_RNITUI31Z0Z_13 ;
    wire \pid_front.O_19 ;
    wire \pid_front.error_d_regZ0Z_17 ;
    wire \pid_front.O_20 ;
    wire \pid_front.error_d_regZ0Z_18 ;
    wire \pid_front.O_21 ;
    wire \pid_front.error_d_regZ0Z_19 ;
    wire \pid_front.O_23 ;
    wire \pid_front.error_d_regZ0Z_21 ;
    wire \pid_front.O_24 ;
    wire \pid_front.error_d_regZ0Z_22 ;
    wire \pid_front.O_17 ;
    wire \pid_front.error_d_regZ0Z_15 ;
    wire \pid_front.O_18 ;
    wire \pid_front.error_d_regZ0Z_16 ;
    wire _gnd_net_;
    wire clk_system_pll_g;
    wire \pid_front.N_789_0 ;
    wire N_940_g;

    defparam \Pc2drone_pll_inst.Pc2drone_pll_inst_pll .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \Pc2drone_pll_inst.Pc2drone_pll_inst_pll .TEST_MODE=1'b0;
    defparam \Pc2drone_pll_inst.Pc2drone_pll_inst_pll .SHIFTREG_DIV_MODE=2'b00;
    defparam \Pc2drone_pll_inst.Pc2drone_pll_inst_pll .PLLOUT_SELECT="GENCLK";
    defparam \Pc2drone_pll_inst.Pc2drone_pll_inst_pll .FILTER_RANGE=3'b001;
    defparam \Pc2drone_pll_inst.Pc2drone_pll_inst_pll .FEEDBACK_PATH="SIMPLE";
    defparam \Pc2drone_pll_inst.Pc2drone_pll_inst_pll .FDA_RELATIVE=4'b0000;
    defparam \Pc2drone_pll_inst.Pc2drone_pll_inst_pll .FDA_FEEDBACK=4'b0000;
    defparam \Pc2drone_pll_inst.Pc2drone_pll_inst_pll .ENABLE_ICEGATE=1'b0;
    defparam \Pc2drone_pll_inst.Pc2drone_pll_inst_pll .DIVR=4'b0000;
    defparam \Pc2drone_pll_inst.Pc2drone_pll_inst_pll .DIVQ=3'b110;
    defparam \Pc2drone_pll_inst.Pc2drone_pll_inst_pll .DIVF=7'b0111111;
    defparam \Pc2drone_pll_inst.Pc2drone_pll_inst_pll .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    PLL40 \Pc2drone_pll_inst.Pc2drone_pll_inst_pll  (
            .PLLOUTGLOBAL(),
            .SDI(GNDG0),
            .BYPASS(GNDG0),
            .RESETB(N__56546),
            .PLLOUTCORE(\Pc2drone_pll_inst.clk_system_pll ),
            .LOCK(),
            .SDO(),
            .SCLK(GNDG0),
            .LATCHINPUTVALUE(GNDG0),
            .EXTFEEDBACK(GNDG0),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLIN(N__87702));
    defparam \pid_alt.un2_error_mulonly_0_24_0 .A_REG=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .NEG_TRIGGER=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .MODE_8x8=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .D_REG=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .C_REG=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .B_SIGNED=1'b1;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .B_REG=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .A_SIGNED=1'b1;
    SB_MAC16 \pid_alt.un2_error_mulonly_0_24_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__56630),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__56638),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_0,dangling_wire_1,dangling_wire_2,dangling_wire_3,dangling_wire_4,dangling_wire_5,dangling_wire_6,dangling_wire_7,dangling_wire_8,dangling_wire_9,dangling_wire_10,dangling_wire_11,dangling_wire_12,dangling_wire_13,dangling_wire_14,dangling_wire_15}),
            .ADDSUBBOT(),
            .A({N__36913,N__36952,N__37009,N__37057,N__37096,N__36409,N__36454,N__36496,N__36535,N__36608,N__36674,N__36736,N__36802,N__36250,N__36300,N__38911}),
            .C({dangling_wire_16,dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21,dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27,dangling_wire_28,dangling_wire_29,dangling_wire_30,dangling_wire_31}),
            .B({dangling_wire_32,dangling_wire_33,dangling_wire_34,dangling_wire_35,dangling_wire_36,dangling_wire_37,dangling_wire_38,dangling_wire_39,N__39180,N__39198,N__38931,N__38184,N__38949,N__38964,N__38976,N__38994}),
            .OHOLDTOP(),
            .O({dangling_wire_40,dangling_wire_41,dangling_wire_42,dangling_wire_43,dangling_wire_44,dangling_wire_45,dangling_wire_46,\pid_alt.O_5_24 ,\pid_alt.O_5_23 ,\pid_alt.O_5_22 ,\pid_alt.O_5_21 ,\pid_alt.O_5_20 ,\pid_alt.O_5_19 ,\pid_alt.O_5_18 ,\pid_alt.O_5_17 ,\pid_alt.O_5_16 ,\pid_alt.O_5_15 ,\pid_alt.O_5_14 ,\pid_alt.O_5_13 ,\pid_alt.O_5_12 ,\pid_alt.O_5_11 ,\pid_alt.O_5_10 ,\pid_alt.O_5_9 ,\pid_alt.O_5_8 ,\pid_alt.O_5_7 ,\pid_alt.O_5_6 ,\pid_alt.O_5_5 ,\pid_alt.O_5_4 ,dangling_wire_47,dangling_wire_48,dangling_wire_49,dangling_wire_50}));
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .A_REG=1'b0;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .NEG_TRIGGER=1'b0;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .MODE_8x8=1'b0;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .D_REG=1'b0;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .C_REG=1'b0;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .B_SIGNED=1'b1;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .B_REG=1'b0;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .A_SIGNED=1'b1;
    SB_MAC16 \pid_alt.un2_error_2_mulonly_0_24_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__56539),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__56580),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_51,dangling_wire_52,dangling_wire_53,dangling_wire_54,dangling_wire_55,dangling_wire_56,dangling_wire_57,dangling_wire_58,dangling_wire_59,dangling_wire_60,dangling_wire_61,dangling_wire_62,dangling_wire_63,dangling_wire_64,dangling_wire_65,dangling_wire_66}),
            .ADDSUBBOT(),
            .A({N__36921,N__36966,N__37014,N__37062,N__37104,N__36417,N__36462,N__36498,N__36543,N__36612,N__36678,N__36741,N__36807,N__36255,N__36299,N__38916}),
            .C({dangling_wire_67,dangling_wire_68,dangling_wire_69,dangling_wire_70,dangling_wire_71,dangling_wire_72,dangling_wire_73,dangling_wire_74,dangling_wire_75,dangling_wire_76,dangling_wire_77,dangling_wire_78,dangling_wire_79,dangling_wire_80,dangling_wire_81,dangling_wire_82}),
            .B({dangling_wire_83,dangling_wire_84,dangling_wire_85,dangling_wire_86,dangling_wire_87,dangling_wire_88,dangling_wire_89,dangling_wire_90,N__32082,N__32106,N__32121,N__32145,N__32133,N__32094,N__32157,N__33417}),
            .OHOLDTOP(),
            .O({dangling_wire_91,dangling_wire_92,dangling_wire_93,dangling_wire_94,dangling_wire_95,dangling_wire_96,dangling_wire_97,\pid_alt.O_3_24 ,\pid_alt.O_3_23 ,\pid_alt.O_3_22 ,\pid_alt.O_3_21 ,\pid_alt.O_3_20 ,\pid_alt.O_3_19 ,\pid_alt.O_3_18 ,\pid_alt.O_3_17 ,\pid_alt.O_3_16 ,\pid_alt.O_3_15 ,\pid_alt.O_3_14 ,\pid_alt.O_3_13 ,\pid_alt.O_3_12 ,\pid_alt.O_3_11 ,\pid_alt.O_3_10 ,\pid_alt.O_3_9 ,\pid_alt.O_3_8 ,\pid_alt.O_3_7 ,\pid_alt.O_3_6 ,\pid_alt.O_3_5 ,\pid_alt.O_3_4 ,dangling_wire_98,dangling_wire_99,dangling_wire_100,dangling_wire_101}));
    defparam \pid_side.un2_error_1_mulonly_0_24_0 .A_REG=1'b0;
    defparam \pid_side.un2_error_1_mulonly_0_24_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pid_side.un2_error_1_mulonly_0_24_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pid_side.un2_error_1_mulonly_0_24_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pid_side.un2_error_1_mulonly_0_24_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pid_side.un2_error_1_mulonly_0_24_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pid_side.un2_error_1_mulonly_0_24_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pid_side.un2_error_1_mulonly_0_24_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pid_side.un2_error_1_mulonly_0_24_0 .NEG_TRIGGER=1'b0;
    defparam \pid_side.un2_error_1_mulonly_0_24_0 .MODE_8x8=1'b0;
    defparam \pid_side.un2_error_1_mulonly_0_24_0 .D_REG=1'b0;
    defparam \pid_side.un2_error_1_mulonly_0_24_0 .C_REG=1'b0;
    defparam \pid_side.un2_error_1_mulonly_0_24_0 .B_SIGNED=1'b1;
    defparam \pid_side.un2_error_1_mulonly_0_24_0 .B_REG=1'b0;
    defparam \pid_side.un2_error_1_mulonly_0_24_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pid_side.un2_error_1_mulonly_0_24_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pid_side.un2_error_1_mulonly_0_24_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pid_side.un2_error_1_mulonly_0_24_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pid_side.un2_error_1_mulonly_0_24_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pid_side.un2_error_1_mulonly_0_24_0 .A_SIGNED=1'b1;
    SB_MAC16 \pid_side.un2_error_1_mulonly_0_24_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__56653),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__56652),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_102,dangling_wire_103,dangling_wire_104,dangling_wire_105,dangling_wire_106,dangling_wire_107,dangling_wire_108,dangling_wire_109,dangling_wire_110,dangling_wire_111,dangling_wire_112,dangling_wire_113,dangling_wire_114,dangling_wire_115,dangling_wire_116,dangling_wire_117}),
            .ADDSUBBOT(),
            .A({N__74930,N__74418,N__74509,N__74071,N__74189,N__74590,N__74657,N__74768,N__75824,N__75892,N__75073,N__75016,N__75197,N__75134,N__73873,N__81060}),
            .C({dangling_wire_118,dangling_wire_119,dangling_wire_120,dangling_wire_121,dangling_wire_122,dangling_wire_123,dangling_wire_124,dangling_wire_125,dangling_wire_126,dangling_wire_127,dangling_wire_128,dangling_wire_129,dangling_wire_130,dangling_wire_131,dangling_wire_132,dangling_wire_133}),
            .B({dangling_wire_134,dangling_wire_135,dangling_wire_136,dangling_wire_137,dangling_wire_138,dangling_wire_139,dangling_wire_140,dangling_wire_141,N__85232,N__54347,N__85061,N__84893,N__83870,N__54377,N__84053,N__83682}),
            .OHOLDTOP(),
            .O({dangling_wire_142,dangling_wire_143,dangling_wire_144,dangling_wire_145,dangling_wire_146,dangling_wire_147,dangling_wire_148,\pid_side.O_1_24 ,\pid_side.O_1_23 ,\pid_side.O_1_22 ,\pid_side.O_1_21 ,\pid_side.O_1_20 ,\pid_side.O_1_19 ,\pid_side.O_1_18 ,\pid_side.O_1_17 ,\pid_side.O_1_16 ,\pid_side.O_1_15 ,\pid_side.O_1_14 ,\pid_side.O_1_13 ,\pid_side.O_1_12 ,\pid_side.O_1_11 ,\pid_side.O_1_10 ,\pid_side.O_1_9 ,\pid_side.O_1_8 ,\pid_side.O_1_7 ,\pid_side.O_1_6 ,\pid_side.O_1_5 ,\pid_side.O_1_4 ,\pid_side.O_1_3 ,\pid_side.O_0_2 ,dangling_wire_149,dangling_wire_150}));
    defparam \pid_side.un2_error_mulonly_0_24_0 .A_REG=1'b0;
    defparam \pid_side.un2_error_mulonly_0_24_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pid_side.un2_error_mulonly_0_24_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pid_side.un2_error_mulonly_0_24_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pid_side.un2_error_mulonly_0_24_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pid_side.un2_error_mulonly_0_24_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pid_side.un2_error_mulonly_0_24_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pid_side.un2_error_mulonly_0_24_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pid_side.un2_error_mulonly_0_24_0 .NEG_TRIGGER=1'b0;
    defparam \pid_side.un2_error_mulonly_0_24_0 .MODE_8x8=1'b0;
    defparam \pid_side.un2_error_mulonly_0_24_0 .D_REG=1'b0;
    defparam \pid_side.un2_error_mulonly_0_24_0 .C_REG=1'b0;
    defparam \pid_side.un2_error_mulonly_0_24_0 .B_SIGNED=1'b1;
    defparam \pid_side.un2_error_mulonly_0_24_0 .B_REG=1'b0;
    defparam \pid_side.un2_error_mulonly_0_24_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pid_side.un2_error_mulonly_0_24_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pid_side.un2_error_mulonly_0_24_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pid_side.un2_error_mulonly_0_24_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pid_side.un2_error_mulonly_0_24_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pid_side.un2_error_mulonly_0_24_0 .A_SIGNED=1'b1;
    SB_MAC16 \pid_side.un2_error_mulonly_0_24_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__56640),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__56639),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_151,dangling_wire_152,dangling_wire_153,dangling_wire_154,dangling_wire_155,dangling_wire_156,dangling_wire_157,dangling_wire_158,dangling_wire_159,dangling_wire_160,dangling_wire_161,dangling_wire_162,dangling_wire_163,dangling_wire_164,dangling_wire_165,dangling_wire_166}),
            .ADDSUBBOT(),
            .A({N__74931,N__74408,N__74513,N__74073,N__74193,N__74592,N__74658,N__74772,N__75831,N__75909,N__75081,N__75027,N__75201,N__75138,N__73881,N__81075}),
            .C({dangling_wire_167,dangling_wire_168,dangling_wire_169,dangling_wire_170,dangling_wire_171,dangling_wire_172,dangling_wire_173,dangling_wire_174,dangling_wire_175,dangling_wire_176,dangling_wire_177,dangling_wire_178,dangling_wire_179,dangling_wire_180,dangling_wire_181,dangling_wire_182}),
            .B({dangling_wire_183,dangling_wire_184,dangling_wire_185,dangling_wire_186,dangling_wire_187,dangling_wire_188,dangling_wire_189,dangling_wire_190,N__51213,N__50675,N__50702,N__32388,N__51249,N__51288,N__82712,N__51318}),
            .OHOLDTOP(),
            .O({dangling_wire_191,dangling_wire_192,dangling_wire_193,dangling_wire_194,dangling_wire_195,dangling_wire_196,dangling_wire_197,\pid_side.O_2_24 ,\pid_side.O_2_23 ,\pid_side.O_2_22 ,\pid_side.O_2_21 ,\pid_side.O_2_20 ,\pid_side.O_2_19 ,\pid_side.O_2_18 ,\pid_side.O_2_17 ,\pid_side.O_2_16 ,\pid_side.O_2_15 ,\pid_side.O_2_14 ,\pid_side.O_2_13 ,\pid_side.O_2_12 ,\pid_side.O_2_11 ,\pid_side.O_2_10 ,\pid_side.O_2_9 ,\pid_side.O_2_8 ,\pid_side.O_2_7 ,\pid_side.O_2_6 ,\pid_side.O_2_5 ,\pid_side.O_2_4 ,\pid_side.O_2_3 ,dangling_wire_198,dangling_wire_199,dangling_wire_200}));
    defparam \pid_front.un2_error_1_mulonly_0_24_0 .A_REG=1'b0;
    defparam \pid_front.un2_error_1_mulonly_0_24_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pid_front.un2_error_1_mulonly_0_24_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pid_front.un2_error_1_mulonly_0_24_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pid_front.un2_error_1_mulonly_0_24_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pid_front.un2_error_1_mulonly_0_24_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pid_front.un2_error_1_mulonly_0_24_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pid_front.un2_error_1_mulonly_0_24_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pid_front.un2_error_1_mulonly_0_24_0 .NEG_TRIGGER=1'b0;
    defparam \pid_front.un2_error_1_mulonly_0_24_0 .MODE_8x8=1'b0;
    defparam \pid_front.un2_error_1_mulonly_0_24_0 .D_REG=1'b0;
    defparam \pid_front.un2_error_1_mulonly_0_24_0 .C_REG=1'b0;
    defparam \pid_front.un2_error_1_mulonly_0_24_0 .B_SIGNED=1'b1;
    defparam \pid_front.un2_error_1_mulonly_0_24_0 .B_REG=1'b0;
    defparam \pid_front.un2_error_1_mulonly_0_24_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pid_front.un2_error_1_mulonly_0_24_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pid_front.un2_error_1_mulonly_0_24_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pid_front.un2_error_1_mulonly_0_24_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pid_front.un2_error_1_mulonly_0_24_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pid_front.un2_error_1_mulonly_0_24_0 .A_SIGNED=1'b1;
    SB_MAC16 \pid_front.un2_error_1_mulonly_0_24_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__56667),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__56666),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_201,dangling_wire_202,dangling_wire_203,dangling_wire_204,dangling_wire_205,dangling_wire_206,dangling_wire_207,dangling_wire_208,dangling_wire_209,dangling_wire_210,dangling_wire_211,dangling_wire_212,dangling_wire_213,dangling_wire_214,dangling_wire_215,dangling_wire_216}),
            .ADDSUBBOT(),
            .A({N__71199,N__72152,N__67253,N__67184,N__67415,N__67334,N__59462,N__62996,N__67682,N__67754,N__67806,N__67850,N__77090,N__77138,N__77204,N__77279}),
            .C({dangling_wire_217,dangling_wire_218,dangling_wire_219,dangling_wire_220,dangling_wire_221,dangling_wire_222,dangling_wire_223,dangling_wire_224,dangling_wire_225,dangling_wire_226,dangling_wire_227,dangling_wire_228,dangling_wire_229,dangling_wire_230,dangling_wire_231,dangling_wire_232}),
            .B({dangling_wire_233,dangling_wire_234,dangling_wire_235,dangling_wire_236,dangling_wire_237,dangling_wire_238,dangling_wire_239,dangling_wire_240,N__85236,N__54348,N__85062,N__84894,N__83874,N__54378,N__84054,N__83681}),
            .OHOLDTOP(),
            .O({dangling_wire_241,dangling_wire_242,dangling_wire_243,dangling_wire_244,dangling_wire_245,dangling_wire_246,dangling_wire_247,\pid_front.O_24 ,\pid_front.O_23 ,\pid_front.O_22 ,\pid_front.O_21 ,\pid_front.O_20 ,\pid_front.O_19 ,\pid_front.O_18 ,\pid_front.O_17 ,\pid_front.O_16 ,\pid_front.O_15 ,\pid_front.O_14 ,\pid_front.O_13 ,\pid_front.O_12 ,\pid_front.O_11 ,\pid_front.O_10 ,\pid_front.O_9 ,\pid_front.O_8 ,\pid_front.O_7 ,\pid_front.O_6 ,\pid_front.O_5 ,\pid_front.O_4 ,\pid_front.O_3 ,\pid_front.O_2 ,dangling_wire_248,dangling_wire_249}));
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .A_REG=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .NEG_TRIGGER=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .MODE_8x8=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .D_REG=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .C_REG=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .B_SIGNED=1'b1;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .B_REG=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .A_SIGNED=1'b1;
    SB_MAC16 \pid_alt.un2_error_1_mulonly_0_24_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__56535),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__56528),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_250,dangling_wire_251,dangling_wire_252,dangling_wire_253,dangling_wire_254,dangling_wire_255,dangling_wire_256,dangling_wire_257,dangling_wire_258,dangling_wire_259,dangling_wire_260,dangling_wire_261,dangling_wire_262,dangling_wire_263,dangling_wire_264,dangling_wire_265}),
            .ADDSUBBOT(),
            .A({N__36914,N__36959,N__37010,N__37058,N__37097,N__36410,N__36455,N__36497,N__36536,N__36604,N__36670,N__36737,N__36803,N__36251,N__36295,N__38915}),
            .C({dangling_wire_266,dangling_wire_267,dangling_wire_268,dangling_wire_269,dangling_wire_270,dangling_wire_271,dangling_wire_272,dangling_wire_273,dangling_wire_274,dangling_wire_275,dangling_wire_276,dangling_wire_277,dangling_wire_278,dangling_wire_279,dangling_wire_280,dangling_wire_281}),
            .B({dangling_wire_282,dangling_wire_283,dangling_wire_284,dangling_wire_285,dangling_wire_286,dangling_wire_287,dangling_wire_288,dangling_wire_289,N__32283,N__32295,N__32307,N__32319,N__32328,N__32337,N__32235,N__32244}),
            .OHOLDTOP(),
            .O({dangling_wire_290,dangling_wire_291,dangling_wire_292,dangling_wire_293,dangling_wire_294,dangling_wire_295,dangling_wire_296,\pid_alt.O_4_24 ,\pid_alt.O_4_23 ,\pid_alt.O_4_22 ,\pid_alt.O_4_21 ,\pid_alt.O_4_20 ,\pid_alt.O_4_19 ,\pid_alt.O_4_18 ,\pid_alt.O_4_17 ,\pid_alt.O_4_16 ,\pid_alt.O_4_15 ,\pid_alt.O_4_14 ,\pid_alt.O_4_13 ,\pid_alt.O_4_12 ,\pid_alt.O_4_11 ,\pid_alt.O_4_10 ,\pid_alt.O_4_9 ,\pid_alt.O_4_8 ,\pid_alt.O_4_7 ,\pid_alt.O_4_6 ,\pid_alt.O_4_5 ,\pid_alt.O_4_4 ,dangling_wire_297,dangling_wire_298,dangling_wire_299,dangling_wire_300}));
    defparam \pid_front.un2_error_mulonly_0_24_0 .A_REG=1'b0;
    defparam \pid_front.un2_error_mulonly_0_24_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pid_front.un2_error_mulonly_0_24_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pid_front.un2_error_mulonly_0_24_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pid_front.un2_error_mulonly_0_24_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pid_front.un2_error_mulonly_0_24_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pid_front.un2_error_mulonly_0_24_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pid_front.un2_error_mulonly_0_24_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pid_front.un2_error_mulonly_0_24_0 .NEG_TRIGGER=1'b0;
    defparam \pid_front.un2_error_mulonly_0_24_0 .MODE_8x8=1'b0;
    defparam \pid_front.un2_error_mulonly_0_24_0 .D_REG=1'b0;
    defparam \pid_front.un2_error_mulonly_0_24_0 .C_REG=1'b0;
    defparam \pid_front.un2_error_mulonly_0_24_0 .B_SIGNED=1'b1;
    defparam \pid_front.un2_error_mulonly_0_24_0 .B_REG=1'b0;
    defparam \pid_front.un2_error_mulonly_0_24_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pid_front.un2_error_mulonly_0_24_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pid_front.un2_error_mulonly_0_24_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pid_front.un2_error_mulonly_0_24_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pid_front.un2_error_mulonly_0_24_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pid_front.un2_error_mulonly_0_24_0 .A_SIGNED=1'b1;
    SB_MAC16 \pid_front.un2_error_mulonly_0_24_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__56506),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__56576),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_301,dangling_wire_302,dangling_wire_303,dangling_wire_304,dangling_wire_305,dangling_wire_306,dangling_wire_307,dangling_wire_308,dangling_wire_309,dangling_wire_310,dangling_wire_311,dangling_wire_312,dangling_wire_313,dangling_wire_314,dangling_wire_315,dangling_wire_316}),
            .ADDSUBBOT(),
            .A({N__71198,N__72153,N__67257,N__67191,N__67416,N__67338,N__59472,N__62997,N__67683,N__67755,N__67805,N__67857,N__77091,N__77145,N__77205,N__77280}),
            .C({dangling_wire_317,dangling_wire_318,dangling_wire_319,dangling_wire_320,dangling_wire_321,dangling_wire_322,dangling_wire_323,dangling_wire_324,dangling_wire_325,dangling_wire_326,dangling_wire_327,dangling_wire_328,dangling_wire_329,dangling_wire_330,dangling_wire_331,dangling_wire_332}),
            .B({dangling_wire_333,dangling_wire_334,dangling_wire_335,dangling_wire_336,dangling_wire_337,dangling_wire_338,dangling_wire_339,dangling_wire_340,N__51209,N__50679,N__50703,N__32378,N__51242,N__51284,N__82716,N__51314}),
            .OHOLDTOP(),
            .O({dangling_wire_341,dangling_wire_342,dangling_wire_343,dangling_wire_344,dangling_wire_345,dangling_wire_346,dangling_wire_347,\pid_front.O_0_24 ,\pid_front.O_0_23 ,\pid_front.O_0_22 ,\pid_front.O_0_21 ,\pid_front.O_0_20 ,\pid_front.O_0_19 ,\pid_front.O_0_18 ,\pid_front.O_0_17 ,\pid_front.O_0_16 ,\pid_front.O_0_15 ,\pid_front.O_0_14 ,\pid_front.O_0_13 ,\pid_front.O_0_12 ,\pid_front.O_0_11 ,\pid_front.O_0_10 ,\pid_front.O_0_9 ,\pid_front.O_0_8 ,\pid_front.O_0_7 ,\pid_front.O_0_6 ,\pid_front.O_0_5 ,\pid_front.O_0_4 ,\pid_front.O_0_3 ,dangling_wire_348,dangling_wire_349,dangling_wire_350}));
    IO_PAD \Pc2drone_pll_inst.Pc2drone_pll_inst_iopad  (
            .OE(VCCG0),
            .DIN(),
            .DOUT(N__87702),
            .PACKAGEPIN(clk_system));
    defparam uart_input_pc_ibuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD uart_input_pc_ibuf_iopad (
            .OE(N__87688),
            .DIN(N__87687),
            .DOUT(N__87686),
            .PACKAGEPIN(uart_input_pc));
    defparam uart_input_pc_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam uart_input_pc_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO uart_input_pc_ibuf_preio (
            .PADOEN(N__87688),
            .PADOUT(N__87687),
            .PADIN(N__87686),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(uart_input_pc_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam debug_CH2_18A_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD debug_CH2_18A_obuf_iopad (
            .OE(N__87679),
            .DIN(N__87678),
            .DOUT(N__87677),
            .PACKAGEPIN(debug_CH2_18A));
    defparam debug_CH2_18A_obuf_preio.NEG_TRIGGER=1'b0;
    defparam debug_CH2_18A_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_CH2_18A_obuf_preio (
            .PADOEN(N__87679),
            .PADOUT(N__87678),
            .PADIN(N__87677),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__40254),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam debug_CH5_31B_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD debug_CH5_31B_obuf_iopad (
            .OE(N__87670),
            .DIN(N__87669),
            .DOUT(N__87668),
            .PACKAGEPIN(debug_CH5_31B));
    defparam debug_CH5_31B_obuf_preio.NEG_TRIGGER=1'b0;
    defparam debug_CH5_31B_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_CH5_31B_obuf_preio (
            .PADOEN(N__87670),
            .PADOUT(N__87669),
            .PADIN(N__87668),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam debug_CH4_2A_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD debug_CH4_2A_obuf_iopad (
            .OE(N__87661),
            .DIN(N__87660),
            .DOUT(N__87659),
            .PACKAGEPIN(debug_CH4_2A));
    defparam debug_CH4_2A_obuf_preio.NEG_TRIGGER=1'b0;
    defparam debug_CH4_2A_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_CH4_2A_obuf_preio (
            .PADOEN(N__87661),
            .PADOUT(N__87660),
            .PADIN(N__87659),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ppm_output_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD ppm_output_obuf_iopad (
            .OE(N__87652),
            .DIN(N__87651),
            .DOUT(N__87650),
            .PACKAGEPIN(ppm_output));
    defparam ppm_output_obuf_preio.NEG_TRIGGER=1'b0;
    defparam ppm_output_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO ppm_output_obuf_preio (
            .PADOEN(N__87652),
            .PADOUT(N__87651),
            .PADIN(N__87650),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__44391),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam debug_CH3_20A_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD debug_CH3_20A_obuf_iopad (
            .OE(N__87643),
            .DIN(N__87642),
            .DOUT(N__87641),
            .PACKAGEPIN(debug_CH3_20A));
    defparam debug_CH3_20A_obuf_preio.NEG_TRIGGER=1'b0;
    defparam debug_CH3_20A_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_CH3_20A_obuf_preio (
            .PADOEN(N__87643),
            .PADOUT(N__87642),
            .PADIN(N__87641),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__41373),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam debug_CH6_5B_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD debug_CH6_5B_obuf_iopad (
            .OE(N__87634),
            .DIN(N__87633),
            .DOUT(N__87632),
            .PACKAGEPIN(debug_CH6_5B));
    defparam debug_CH6_5B_obuf_preio.NEG_TRIGGER=1'b0;
    defparam debug_CH6_5B_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_CH6_5B_obuf_preio (
            .PADOEN(N__87634),
            .PADOUT(N__87633),
            .PADIN(N__87632),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam uart_input_drone_ibuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD uart_input_drone_ibuf_iopad (
            .OE(N__87625),
            .DIN(N__87624),
            .DOUT(N__87623),
            .PACKAGEPIN(uart_input_drone));
    defparam uart_input_drone_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam uart_input_drone_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO uart_input_drone_ibuf_preio (
            .PADOEN(N__87625),
            .PADOUT(N__87624),
            .PADIN(N__87623),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(uart_input_drone_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam debug_CH0_16A_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD debug_CH0_16A_obuf_iopad (
            .OE(N__87616),
            .DIN(N__87615),
            .DOUT(N__87614),
            .PACKAGEPIN(debug_CH0_16A));
    defparam debug_CH0_16A_obuf_preio.NEG_TRIGGER=1'b0;
    defparam debug_CH0_16A_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_CH0_16A_obuf_preio (
            .PADOEN(N__87616),
            .PADOUT(N__87615),
            .PADIN(N__87614),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__47997),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam debug_CH1_0A_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD debug_CH1_0A_obuf_iopad (
            .OE(N__87607),
            .DIN(N__87606),
            .DOUT(N__87605),
            .PACKAGEPIN(debug_CH1_0A));
    defparam debug_CH1_0A_obuf_preio.NEG_TRIGGER=1'b0;
    defparam debug_CH1_0A_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_CH1_0A_obuf_preio (
            .PADOEN(N__87607),
            .PADOUT(N__87606),
            .PADIN(N__87605),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__59964),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__21317 (
            .O(N__87588),
            .I(N__87585));
    LocalMux I__21316 (
            .O(N__87585),
            .I(N__87582));
    Odrv4 I__21315 (
            .O(N__87582),
            .I(\pid_front.O_19 ));
    InMux I__21314 (
            .O(N__87579),
            .I(N__87570));
    InMux I__21313 (
            .O(N__87578),
            .I(N__87570));
    InMux I__21312 (
            .O(N__87577),
            .I(N__87570));
    LocalMux I__21311 (
            .O(N__87570),
            .I(N__87567));
    Span4Mux_h I__21310 (
            .O(N__87567),
            .I(N__87564));
    Span4Mux_h I__21309 (
            .O(N__87564),
            .I(N__87561));
    Span4Mux_h I__21308 (
            .O(N__87561),
            .I(N__87558));
    Odrv4 I__21307 (
            .O(N__87558),
            .I(\pid_front.error_d_regZ0Z_17 ));
    InMux I__21306 (
            .O(N__87555),
            .I(N__87552));
    LocalMux I__21305 (
            .O(N__87552),
            .I(N__87549));
    Odrv4 I__21304 (
            .O(N__87549),
            .I(\pid_front.O_20 ));
    InMux I__21303 (
            .O(N__87546),
            .I(N__87540));
    InMux I__21302 (
            .O(N__87545),
            .I(N__87540));
    LocalMux I__21301 (
            .O(N__87540),
            .I(N__87536));
    InMux I__21300 (
            .O(N__87539),
            .I(N__87533));
    Span4Mux_h I__21299 (
            .O(N__87536),
            .I(N__87530));
    LocalMux I__21298 (
            .O(N__87533),
            .I(N__87527));
    Span4Mux_h I__21297 (
            .O(N__87530),
            .I(N__87524));
    Span12Mux_h I__21296 (
            .O(N__87527),
            .I(N__87521));
    Odrv4 I__21295 (
            .O(N__87524),
            .I(\pid_front.error_d_regZ0Z_18 ));
    Odrv12 I__21294 (
            .O(N__87521),
            .I(\pid_front.error_d_regZ0Z_18 ));
    InMux I__21293 (
            .O(N__87516),
            .I(N__87513));
    LocalMux I__21292 (
            .O(N__87513),
            .I(N__87510));
    Odrv4 I__21291 (
            .O(N__87510),
            .I(\pid_front.O_21 ));
    InMux I__21290 (
            .O(N__87507),
            .I(N__87504));
    LocalMux I__21289 (
            .O(N__87504),
            .I(N__87499));
    InMux I__21288 (
            .O(N__87503),
            .I(N__87494));
    InMux I__21287 (
            .O(N__87502),
            .I(N__87494));
    Sp12to4 I__21286 (
            .O(N__87499),
            .I(N__87491));
    LocalMux I__21285 (
            .O(N__87494),
            .I(N__87488));
    Span12Mux_h I__21284 (
            .O(N__87491),
            .I(N__87485));
    Span12Mux_h I__21283 (
            .O(N__87488),
            .I(N__87482));
    Odrv12 I__21282 (
            .O(N__87485),
            .I(\pid_front.error_d_regZ0Z_19 ));
    Odrv12 I__21281 (
            .O(N__87482),
            .I(\pid_front.error_d_regZ0Z_19 ));
    InMux I__21280 (
            .O(N__87477),
            .I(N__87474));
    LocalMux I__21279 (
            .O(N__87474),
            .I(N__87471));
    Span4Mux_h I__21278 (
            .O(N__87471),
            .I(N__87468));
    Odrv4 I__21277 (
            .O(N__87468),
            .I(\pid_front.O_23 ));
    InMux I__21276 (
            .O(N__87465),
            .I(N__87460));
    InMux I__21275 (
            .O(N__87464),
            .I(N__87455));
    InMux I__21274 (
            .O(N__87463),
            .I(N__87455));
    LocalMux I__21273 (
            .O(N__87460),
            .I(N__87450));
    LocalMux I__21272 (
            .O(N__87455),
            .I(N__87450));
    Span12Mux_v I__21271 (
            .O(N__87450),
            .I(N__87447));
    Span12Mux_h I__21270 (
            .O(N__87447),
            .I(N__87444));
    Odrv12 I__21269 (
            .O(N__87444),
            .I(\pid_front.error_d_regZ0Z_21 ));
    InMux I__21268 (
            .O(N__87441),
            .I(N__87438));
    LocalMux I__21267 (
            .O(N__87438),
            .I(N__87435));
    Span4Mux_h I__21266 (
            .O(N__87435),
            .I(N__87432));
    Odrv4 I__21265 (
            .O(N__87432),
            .I(\pid_front.O_24 ));
    CascadeMux I__21264 (
            .O(N__87429),
            .I(N__87426));
    InMux I__21263 (
            .O(N__87426),
            .I(N__87409));
    InMux I__21262 (
            .O(N__87425),
            .I(N__87409));
    InMux I__21261 (
            .O(N__87424),
            .I(N__87404));
    InMux I__21260 (
            .O(N__87423),
            .I(N__87404));
    InMux I__21259 (
            .O(N__87422),
            .I(N__87398));
    InMux I__21258 (
            .O(N__87421),
            .I(N__87398));
    InMux I__21257 (
            .O(N__87420),
            .I(N__87389));
    InMux I__21256 (
            .O(N__87419),
            .I(N__87389));
    InMux I__21255 (
            .O(N__87418),
            .I(N__87389));
    InMux I__21254 (
            .O(N__87417),
            .I(N__87389));
    InMux I__21253 (
            .O(N__87416),
            .I(N__87382));
    InMux I__21252 (
            .O(N__87415),
            .I(N__87382));
    InMux I__21251 (
            .O(N__87414),
            .I(N__87382));
    LocalMux I__21250 (
            .O(N__87409),
            .I(N__87379));
    LocalMux I__21249 (
            .O(N__87404),
            .I(N__87376));
    InMux I__21248 (
            .O(N__87403),
            .I(N__87373));
    LocalMux I__21247 (
            .O(N__87398),
            .I(N__87366));
    LocalMux I__21246 (
            .O(N__87389),
            .I(N__87366));
    LocalMux I__21245 (
            .O(N__87382),
            .I(N__87366));
    Span4Mux_h I__21244 (
            .O(N__87379),
            .I(N__87363));
    Span4Mux_v I__21243 (
            .O(N__87376),
            .I(N__87360));
    LocalMux I__21242 (
            .O(N__87373),
            .I(N__87355));
    Span4Mux_v I__21241 (
            .O(N__87366),
            .I(N__87355));
    Span4Mux_h I__21240 (
            .O(N__87363),
            .I(N__87352));
    Span4Mux_h I__21239 (
            .O(N__87360),
            .I(N__87347));
    Span4Mux_h I__21238 (
            .O(N__87355),
            .I(N__87347));
    Span4Mux_h I__21237 (
            .O(N__87352),
            .I(N__87344));
    Sp12to4 I__21236 (
            .O(N__87347),
            .I(N__87341));
    Span4Mux_h I__21235 (
            .O(N__87344),
            .I(N__87338));
    Odrv12 I__21234 (
            .O(N__87341),
            .I(\pid_front.error_d_regZ0Z_22 ));
    Odrv4 I__21233 (
            .O(N__87338),
            .I(\pid_front.error_d_regZ0Z_22 ));
    InMux I__21232 (
            .O(N__87333),
            .I(N__87330));
    LocalMux I__21231 (
            .O(N__87330),
            .I(N__87327));
    Odrv4 I__21230 (
            .O(N__87327),
            .I(\pid_front.O_17 ));
    InMux I__21229 (
            .O(N__87324),
            .I(N__87315));
    InMux I__21228 (
            .O(N__87323),
            .I(N__87315));
    InMux I__21227 (
            .O(N__87322),
            .I(N__87315));
    LocalMux I__21226 (
            .O(N__87315),
            .I(N__87312));
    Span12Mux_h I__21225 (
            .O(N__87312),
            .I(N__87309));
    Span12Mux_h I__21224 (
            .O(N__87309),
            .I(N__87306));
    Odrv12 I__21223 (
            .O(N__87306),
            .I(\pid_front.error_d_regZ0Z_15 ));
    InMux I__21222 (
            .O(N__87303),
            .I(N__87300));
    LocalMux I__21221 (
            .O(N__87300),
            .I(\pid_front.O_18 ));
    InMux I__21220 (
            .O(N__87297),
            .I(N__87288));
    InMux I__21219 (
            .O(N__87296),
            .I(N__87288));
    InMux I__21218 (
            .O(N__87295),
            .I(N__87288));
    LocalMux I__21217 (
            .O(N__87288),
            .I(N__87285));
    Span12Mux_h I__21216 (
            .O(N__87285),
            .I(N__87282));
    Odrv12 I__21215 (
            .O(N__87282),
            .I(\pid_front.error_d_regZ0Z_16 ));
    ClkMux I__21214 (
            .O(N__87279),
            .I(N__86346));
    ClkMux I__21213 (
            .O(N__87278),
            .I(N__86346));
    ClkMux I__21212 (
            .O(N__87277),
            .I(N__86346));
    ClkMux I__21211 (
            .O(N__87276),
            .I(N__86346));
    ClkMux I__21210 (
            .O(N__87275),
            .I(N__86346));
    ClkMux I__21209 (
            .O(N__87274),
            .I(N__86346));
    ClkMux I__21208 (
            .O(N__87273),
            .I(N__86346));
    ClkMux I__21207 (
            .O(N__87272),
            .I(N__86346));
    ClkMux I__21206 (
            .O(N__87271),
            .I(N__86346));
    ClkMux I__21205 (
            .O(N__87270),
            .I(N__86346));
    ClkMux I__21204 (
            .O(N__87269),
            .I(N__86346));
    ClkMux I__21203 (
            .O(N__87268),
            .I(N__86346));
    ClkMux I__21202 (
            .O(N__87267),
            .I(N__86346));
    ClkMux I__21201 (
            .O(N__87266),
            .I(N__86346));
    ClkMux I__21200 (
            .O(N__87265),
            .I(N__86346));
    ClkMux I__21199 (
            .O(N__87264),
            .I(N__86346));
    ClkMux I__21198 (
            .O(N__87263),
            .I(N__86346));
    ClkMux I__21197 (
            .O(N__87262),
            .I(N__86346));
    ClkMux I__21196 (
            .O(N__87261),
            .I(N__86346));
    ClkMux I__21195 (
            .O(N__87260),
            .I(N__86346));
    ClkMux I__21194 (
            .O(N__87259),
            .I(N__86346));
    ClkMux I__21193 (
            .O(N__87258),
            .I(N__86346));
    ClkMux I__21192 (
            .O(N__87257),
            .I(N__86346));
    ClkMux I__21191 (
            .O(N__87256),
            .I(N__86346));
    ClkMux I__21190 (
            .O(N__87255),
            .I(N__86346));
    ClkMux I__21189 (
            .O(N__87254),
            .I(N__86346));
    ClkMux I__21188 (
            .O(N__87253),
            .I(N__86346));
    ClkMux I__21187 (
            .O(N__87252),
            .I(N__86346));
    ClkMux I__21186 (
            .O(N__87251),
            .I(N__86346));
    ClkMux I__21185 (
            .O(N__87250),
            .I(N__86346));
    ClkMux I__21184 (
            .O(N__87249),
            .I(N__86346));
    ClkMux I__21183 (
            .O(N__87248),
            .I(N__86346));
    ClkMux I__21182 (
            .O(N__87247),
            .I(N__86346));
    ClkMux I__21181 (
            .O(N__87246),
            .I(N__86346));
    ClkMux I__21180 (
            .O(N__87245),
            .I(N__86346));
    ClkMux I__21179 (
            .O(N__87244),
            .I(N__86346));
    ClkMux I__21178 (
            .O(N__87243),
            .I(N__86346));
    ClkMux I__21177 (
            .O(N__87242),
            .I(N__86346));
    ClkMux I__21176 (
            .O(N__87241),
            .I(N__86346));
    ClkMux I__21175 (
            .O(N__87240),
            .I(N__86346));
    ClkMux I__21174 (
            .O(N__87239),
            .I(N__86346));
    ClkMux I__21173 (
            .O(N__87238),
            .I(N__86346));
    ClkMux I__21172 (
            .O(N__87237),
            .I(N__86346));
    ClkMux I__21171 (
            .O(N__87236),
            .I(N__86346));
    ClkMux I__21170 (
            .O(N__87235),
            .I(N__86346));
    ClkMux I__21169 (
            .O(N__87234),
            .I(N__86346));
    ClkMux I__21168 (
            .O(N__87233),
            .I(N__86346));
    ClkMux I__21167 (
            .O(N__87232),
            .I(N__86346));
    ClkMux I__21166 (
            .O(N__87231),
            .I(N__86346));
    ClkMux I__21165 (
            .O(N__87230),
            .I(N__86346));
    ClkMux I__21164 (
            .O(N__87229),
            .I(N__86346));
    ClkMux I__21163 (
            .O(N__87228),
            .I(N__86346));
    ClkMux I__21162 (
            .O(N__87227),
            .I(N__86346));
    ClkMux I__21161 (
            .O(N__87226),
            .I(N__86346));
    ClkMux I__21160 (
            .O(N__87225),
            .I(N__86346));
    ClkMux I__21159 (
            .O(N__87224),
            .I(N__86346));
    ClkMux I__21158 (
            .O(N__87223),
            .I(N__86346));
    ClkMux I__21157 (
            .O(N__87222),
            .I(N__86346));
    ClkMux I__21156 (
            .O(N__87221),
            .I(N__86346));
    ClkMux I__21155 (
            .O(N__87220),
            .I(N__86346));
    ClkMux I__21154 (
            .O(N__87219),
            .I(N__86346));
    ClkMux I__21153 (
            .O(N__87218),
            .I(N__86346));
    ClkMux I__21152 (
            .O(N__87217),
            .I(N__86346));
    ClkMux I__21151 (
            .O(N__87216),
            .I(N__86346));
    ClkMux I__21150 (
            .O(N__87215),
            .I(N__86346));
    ClkMux I__21149 (
            .O(N__87214),
            .I(N__86346));
    ClkMux I__21148 (
            .O(N__87213),
            .I(N__86346));
    ClkMux I__21147 (
            .O(N__87212),
            .I(N__86346));
    ClkMux I__21146 (
            .O(N__87211),
            .I(N__86346));
    ClkMux I__21145 (
            .O(N__87210),
            .I(N__86346));
    ClkMux I__21144 (
            .O(N__87209),
            .I(N__86346));
    ClkMux I__21143 (
            .O(N__87208),
            .I(N__86346));
    ClkMux I__21142 (
            .O(N__87207),
            .I(N__86346));
    ClkMux I__21141 (
            .O(N__87206),
            .I(N__86346));
    ClkMux I__21140 (
            .O(N__87205),
            .I(N__86346));
    ClkMux I__21139 (
            .O(N__87204),
            .I(N__86346));
    ClkMux I__21138 (
            .O(N__87203),
            .I(N__86346));
    ClkMux I__21137 (
            .O(N__87202),
            .I(N__86346));
    ClkMux I__21136 (
            .O(N__87201),
            .I(N__86346));
    ClkMux I__21135 (
            .O(N__87200),
            .I(N__86346));
    ClkMux I__21134 (
            .O(N__87199),
            .I(N__86346));
    ClkMux I__21133 (
            .O(N__87198),
            .I(N__86346));
    ClkMux I__21132 (
            .O(N__87197),
            .I(N__86346));
    ClkMux I__21131 (
            .O(N__87196),
            .I(N__86346));
    ClkMux I__21130 (
            .O(N__87195),
            .I(N__86346));
    ClkMux I__21129 (
            .O(N__87194),
            .I(N__86346));
    ClkMux I__21128 (
            .O(N__87193),
            .I(N__86346));
    ClkMux I__21127 (
            .O(N__87192),
            .I(N__86346));
    ClkMux I__21126 (
            .O(N__87191),
            .I(N__86346));
    ClkMux I__21125 (
            .O(N__87190),
            .I(N__86346));
    ClkMux I__21124 (
            .O(N__87189),
            .I(N__86346));
    ClkMux I__21123 (
            .O(N__87188),
            .I(N__86346));
    ClkMux I__21122 (
            .O(N__87187),
            .I(N__86346));
    ClkMux I__21121 (
            .O(N__87186),
            .I(N__86346));
    ClkMux I__21120 (
            .O(N__87185),
            .I(N__86346));
    ClkMux I__21119 (
            .O(N__87184),
            .I(N__86346));
    ClkMux I__21118 (
            .O(N__87183),
            .I(N__86346));
    ClkMux I__21117 (
            .O(N__87182),
            .I(N__86346));
    ClkMux I__21116 (
            .O(N__87181),
            .I(N__86346));
    ClkMux I__21115 (
            .O(N__87180),
            .I(N__86346));
    ClkMux I__21114 (
            .O(N__87179),
            .I(N__86346));
    ClkMux I__21113 (
            .O(N__87178),
            .I(N__86346));
    ClkMux I__21112 (
            .O(N__87177),
            .I(N__86346));
    ClkMux I__21111 (
            .O(N__87176),
            .I(N__86346));
    ClkMux I__21110 (
            .O(N__87175),
            .I(N__86346));
    ClkMux I__21109 (
            .O(N__87174),
            .I(N__86346));
    ClkMux I__21108 (
            .O(N__87173),
            .I(N__86346));
    ClkMux I__21107 (
            .O(N__87172),
            .I(N__86346));
    ClkMux I__21106 (
            .O(N__87171),
            .I(N__86346));
    ClkMux I__21105 (
            .O(N__87170),
            .I(N__86346));
    ClkMux I__21104 (
            .O(N__87169),
            .I(N__86346));
    ClkMux I__21103 (
            .O(N__87168),
            .I(N__86346));
    ClkMux I__21102 (
            .O(N__87167),
            .I(N__86346));
    ClkMux I__21101 (
            .O(N__87166),
            .I(N__86346));
    ClkMux I__21100 (
            .O(N__87165),
            .I(N__86346));
    ClkMux I__21099 (
            .O(N__87164),
            .I(N__86346));
    ClkMux I__21098 (
            .O(N__87163),
            .I(N__86346));
    ClkMux I__21097 (
            .O(N__87162),
            .I(N__86346));
    ClkMux I__21096 (
            .O(N__87161),
            .I(N__86346));
    ClkMux I__21095 (
            .O(N__87160),
            .I(N__86346));
    ClkMux I__21094 (
            .O(N__87159),
            .I(N__86346));
    ClkMux I__21093 (
            .O(N__87158),
            .I(N__86346));
    ClkMux I__21092 (
            .O(N__87157),
            .I(N__86346));
    ClkMux I__21091 (
            .O(N__87156),
            .I(N__86346));
    ClkMux I__21090 (
            .O(N__87155),
            .I(N__86346));
    ClkMux I__21089 (
            .O(N__87154),
            .I(N__86346));
    ClkMux I__21088 (
            .O(N__87153),
            .I(N__86346));
    ClkMux I__21087 (
            .O(N__87152),
            .I(N__86346));
    ClkMux I__21086 (
            .O(N__87151),
            .I(N__86346));
    ClkMux I__21085 (
            .O(N__87150),
            .I(N__86346));
    ClkMux I__21084 (
            .O(N__87149),
            .I(N__86346));
    ClkMux I__21083 (
            .O(N__87148),
            .I(N__86346));
    ClkMux I__21082 (
            .O(N__87147),
            .I(N__86346));
    ClkMux I__21081 (
            .O(N__87146),
            .I(N__86346));
    ClkMux I__21080 (
            .O(N__87145),
            .I(N__86346));
    ClkMux I__21079 (
            .O(N__87144),
            .I(N__86346));
    ClkMux I__21078 (
            .O(N__87143),
            .I(N__86346));
    ClkMux I__21077 (
            .O(N__87142),
            .I(N__86346));
    ClkMux I__21076 (
            .O(N__87141),
            .I(N__86346));
    ClkMux I__21075 (
            .O(N__87140),
            .I(N__86346));
    ClkMux I__21074 (
            .O(N__87139),
            .I(N__86346));
    ClkMux I__21073 (
            .O(N__87138),
            .I(N__86346));
    ClkMux I__21072 (
            .O(N__87137),
            .I(N__86346));
    ClkMux I__21071 (
            .O(N__87136),
            .I(N__86346));
    ClkMux I__21070 (
            .O(N__87135),
            .I(N__86346));
    ClkMux I__21069 (
            .O(N__87134),
            .I(N__86346));
    ClkMux I__21068 (
            .O(N__87133),
            .I(N__86346));
    ClkMux I__21067 (
            .O(N__87132),
            .I(N__86346));
    ClkMux I__21066 (
            .O(N__87131),
            .I(N__86346));
    ClkMux I__21065 (
            .O(N__87130),
            .I(N__86346));
    ClkMux I__21064 (
            .O(N__87129),
            .I(N__86346));
    ClkMux I__21063 (
            .O(N__87128),
            .I(N__86346));
    ClkMux I__21062 (
            .O(N__87127),
            .I(N__86346));
    ClkMux I__21061 (
            .O(N__87126),
            .I(N__86346));
    ClkMux I__21060 (
            .O(N__87125),
            .I(N__86346));
    ClkMux I__21059 (
            .O(N__87124),
            .I(N__86346));
    ClkMux I__21058 (
            .O(N__87123),
            .I(N__86346));
    ClkMux I__21057 (
            .O(N__87122),
            .I(N__86346));
    ClkMux I__21056 (
            .O(N__87121),
            .I(N__86346));
    ClkMux I__21055 (
            .O(N__87120),
            .I(N__86346));
    ClkMux I__21054 (
            .O(N__87119),
            .I(N__86346));
    ClkMux I__21053 (
            .O(N__87118),
            .I(N__86346));
    ClkMux I__21052 (
            .O(N__87117),
            .I(N__86346));
    ClkMux I__21051 (
            .O(N__87116),
            .I(N__86346));
    ClkMux I__21050 (
            .O(N__87115),
            .I(N__86346));
    ClkMux I__21049 (
            .O(N__87114),
            .I(N__86346));
    ClkMux I__21048 (
            .O(N__87113),
            .I(N__86346));
    ClkMux I__21047 (
            .O(N__87112),
            .I(N__86346));
    ClkMux I__21046 (
            .O(N__87111),
            .I(N__86346));
    ClkMux I__21045 (
            .O(N__87110),
            .I(N__86346));
    ClkMux I__21044 (
            .O(N__87109),
            .I(N__86346));
    ClkMux I__21043 (
            .O(N__87108),
            .I(N__86346));
    ClkMux I__21042 (
            .O(N__87107),
            .I(N__86346));
    ClkMux I__21041 (
            .O(N__87106),
            .I(N__86346));
    ClkMux I__21040 (
            .O(N__87105),
            .I(N__86346));
    ClkMux I__21039 (
            .O(N__87104),
            .I(N__86346));
    ClkMux I__21038 (
            .O(N__87103),
            .I(N__86346));
    ClkMux I__21037 (
            .O(N__87102),
            .I(N__86346));
    ClkMux I__21036 (
            .O(N__87101),
            .I(N__86346));
    ClkMux I__21035 (
            .O(N__87100),
            .I(N__86346));
    ClkMux I__21034 (
            .O(N__87099),
            .I(N__86346));
    ClkMux I__21033 (
            .O(N__87098),
            .I(N__86346));
    ClkMux I__21032 (
            .O(N__87097),
            .I(N__86346));
    ClkMux I__21031 (
            .O(N__87096),
            .I(N__86346));
    ClkMux I__21030 (
            .O(N__87095),
            .I(N__86346));
    ClkMux I__21029 (
            .O(N__87094),
            .I(N__86346));
    ClkMux I__21028 (
            .O(N__87093),
            .I(N__86346));
    ClkMux I__21027 (
            .O(N__87092),
            .I(N__86346));
    ClkMux I__21026 (
            .O(N__87091),
            .I(N__86346));
    ClkMux I__21025 (
            .O(N__87090),
            .I(N__86346));
    ClkMux I__21024 (
            .O(N__87089),
            .I(N__86346));
    ClkMux I__21023 (
            .O(N__87088),
            .I(N__86346));
    ClkMux I__21022 (
            .O(N__87087),
            .I(N__86346));
    ClkMux I__21021 (
            .O(N__87086),
            .I(N__86346));
    ClkMux I__21020 (
            .O(N__87085),
            .I(N__86346));
    ClkMux I__21019 (
            .O(N__87084),
            .I(N__86346));
    ClkMux I__21018 (
            .O(N__87083),
            .I(N__86346));
    ClkMux I__21017 (
            .O(N__87082),
            .I(N__86346));
    ClkMux I__21016 (
            .O(N__87081),
            .I(N__86346));
    ClkMux I__21015 (
            .O(N__87080),
            .I(N__86346));
    ClkMux I__21014 (
            .O(N__87079),
            .I(N__86346));
    ClkMux I__21013 (
            .O(N__87078),
            .I(N__86346));
    ClkMux I__21012 (
            .O(N__87077),
            .I(N__86346));
    ClkMux I__21011 (
            .O(N__87076),
            .I(N__86346));
    ClkMux I__21010 (
            .O(N__87075),
            .I(N__86346));
    ClkMux I__21009 (
            .O(N__87074),
            .I(N__86346));
    ClkMux I__21008 (
            .O(N__87073),
            .I(N__86346));
    ClkMux I__21007 (
            .O(N__87072),
            .I(N__86346));
    ClkMux I__21006 (
            .O(N__87071),
            .I(N__86346));
    ClkMux I__21005 (
            .O(N__87070),
            .I(N__86346));
    ClkMux I__21004 (
            .O(N__87069),
            .I(N__86346));
    ClkMux I__21003 (
            .O(N__87068),
            .I(N__86346));
    ClkMux I__21002 (
            .O(N__87067),
            .I(N__86346));
    ClkMux I__21001 (
            .O(N__87066),
            .I(N__86346));
    ClkMux I__21000 (
            .O(N__87065),
            .I(N__86346));
    ClkMux I__20999 (
            .O(N__87064),
            .I(N__86346));
    ClkMux I__20998 (
            .O(N__87063),
            .I(N__86346));
    ClkMux I__20997 (
            .O(N__87062),
            .I(N__86346));
    ClkMux I__20996 (
            .O(N__87061),
            .I(N__86346));
    ClkMux I__20995 (
            .O(N__87060),
            .I(N__86346));
    ClkMux I__20994 (
            .O(N__87059),
            .I(N__86346));
    ClkMux I__20993 (
            .O(N__87058),
            .I(N__86346));
    ClkMux I__20992 (
            .O(N__87057),
            .I(N__86346));
    ClkMux I__20991 (
            .O(N__87056),
            .I(N__86346));
    ClkMux I__20990 (
            .O(N__87055),
            .I(N__86346));
    ClkMux I__20989 (
            .O(N__87054),
            .I(N__86346));
    ClkMux I__20988 (
            .O(N__87053),
            .I(N__86346));
    ClkMux I__20987 (
            .O(N__87052),
            .I(N__86346));
    ClkMux I__20986 (
            .O(N__87051),
            .I(N__86346));
    ClkMux I__20985 (
            .O(N__87050),
            .I(N__86346));
    ClkMux I__20984 (
            .O(N__87049),
            .I(N__86346));
    ClkMux I__20983 (
            .O(N__87048),
            .I(N__86346));
    ClkMux I__20982 (
            .O(N__87047),
            .I(N__86346));
    ClkMux I__20981 (
            .O(N__87046),
            .I(N__86346));
    ClkMux I__20980 (
            .O(N__87045),
            .I(N__86346));
    ClkMux I__20979 (
            .O(N__87044),
            .I(N__86346));
    ClkMux I__20978 (
            .O(N__87043),
            .I(N__86346));
    ClkMux I__20977 (
            .O(N__87042),
            .I(N__86346));
    ClkMux I__20976 (
            .O(N__87041),
            .I(N__86346));
    ClkMux I__20975 (
            .O(N__87040),
            .I(N__86346));
    ClkMux I__20974 (
            .O(N__87039),
            .I(N__86346));
    ClkMux I__20973 (
            .O(N__87038),
            .I(N__86346));
    ClkMux I__20972 (
            .O(N__87037),
            .I(N__86346));
    ClkMux I__20971 (
            .O(N__87036),
            .I(N__86346));
    ClkMux I__20970 (
            .O(N__87035),
            .I(N__86346));
    ClkMux I__20969 (
            .O(N__87034),
            .I(N__86346));
    ClkMux I__20968 (
            .O(N__87033),
            .I(N__86346));
    ClkMux I__20967 (
            .O(N__87032),
            .I(N__86346));
    ClkMux I__20966 (
            .O(N__87031),
            .I(N__86346));
    ClkMux I__20965 (
            .O(N__87030),
            .I(N__86346));
    ClkMux I__20964 (
            .O(N__87029),
            .I(N__86346));
    ClkMux I__20963 (
            .O(N__87028),
            .I(N__86346));
    ClkMux I__20962 (
            .O(N__87027),
            .I(N__86346));
    ClkMux I__20961 (
            .O(N__87026),
            .I(N__86346));
    ClkMux I__20960 (
            .O(N__87025),
            .I(N__86346));
    ClkMux I__20959 (
            .O(N__87024),
            .I(N__86346));
    ClkMux I__20958 (
            .O(N__87023),
            .I(N__86346));
    ClkMux I__20957 (
            .O(N__87022),
            .I(N__86346));
    ClkMux I__20956 (
            .O(N__87021),
            .I(N__86346));
    ClkMux I__20955 (
            .O(N__87020),
            .I(N__86346));
    ClkMux I__20954 (
            .O(N__87019),
            .I(N__86346));
    ClkMux I__20953 (
            .O(N__87018),
            .I(N__86346));
    ClkMux I__20952 (
            .O(N__87017),
            .I(N__86346));
    ClkMux I__20951 (
            .O(N__87016),
            .I(N__86346));
    ClkMux I__20950 (
            .O(N__87015),
            .I(N__86346));
    ClkMux I__20949 (
            .O(N__87014),
            .I(N__86346));
    ClkMux I__20948 (
            .O(N__87013),
            .I(N__86346));
    ClkMux I__20947 (
            .O(N__87012),
            .I(N__86346));
    ClkMux I__20946 (
            .O(N__87011),
            .I(N__86346));
    ClkMux I__20945 (
            .O(N__87010),
            .I(N__86346));
    ClkMux I__20944 (
            .O(N__87009),
            .I(N__86346));
    ClkMux I__20943 (
            .O(N__87008),
            .I(N__86346));
    ClkMux I__20942 (
            .O(N__87007),
            .I(N__86346));
    ClkMux I__20941 (
            .O(N__87006),
            .I(N__86346));
    ClkMux I__20940 (
            .O(N__87005),
            .I(N__86346));
    ClkMux I__20939 (
            .O(N__87004),
            .I(N__86346));
    ClkMux I__20938 (
            .O(N__87003),
            .I(N__86346));
    ClkMux I__20937 (
            .O(N__87002),
            .I(N__86346));
    ClkMux I__20936 (
            .O(N__87001),
            .I(N__86346));
    ClkMux I__20935 (
            .O(N__87000),
            .I(N__86346));
    ClkMux I__20934 (
            .O(N__86999),
            .I(N__86346));
    ClkMux I__20933 (
            .O(N__86998),
            .I(N__86346));
    ClkMux I__20932 (
            .O(N__86997),
            .I(N__86346));
    ClkMux I__20931 (
            .O(N__86996),
            .I(N__86346));
    ClkMux I__20930 (
            .O(N__86995),
            .I(N__86346));
    ClkMux I__20929 (
            .O(N__86994),
            .I(N__86346));
    ClkMux I__20928 (
            .O(N__86993),
            .I(N__86346));
    ClkMux I__20927 (
            .O(N__86992),
            .I(N__86346));
    ClkMux I__20926 (
            .O(N__86991),
            .I(N__86346));
    ClkMux I__20925 (
            .O(N__86990),
            .I(N__86346));
    ClkMux I__20924 (
            .O(N__86989),
            .I(N__86346));
    ClkMux I__20923 (
            .O(N__86988),
            .I(N__86346));
    ClkMux I__20922 (
            .O(N__86987),
            .I(N__86346));
    ClkMux I__20921 (
            .O(N__86986),
            .I(N__86346));
    ClkMux I__20920 (
            .O(N__86985),
            .I(N__86346));
    ClkMux I__20919 (
            .O(N__86984),
            .I(N__86346));
    ClkMux I__20918 (
            .O(N__86983),
            .I(N__86346));
    ClkMux I__20917 (
            .O(N__86982),
            .I(N__86346));
    ClkMux I__20916 (
            .O(N__86981),
            .I(N__86346));
    ClkMux I__20915 (
            .O(N__86980),
            .I(N__86346));
    ClkMux I__20914 (
            .O(N__86979),
            .I(N__86346));
    ClkMux I__20913 (
            .O(N__86978),
            .I(N__86346));
    ClkMux I__20912 (
            .O(N__86977),
            .I(N__86346));
    ClkMux I__20911 (
            .O(N__86976),
            .I(N__86346));
    ClkMux I__20910 (
            .O(N__86975),
            .I(N__86346));
    ClkMux I__20909 (
            .O(N__86974),
            .I(N__86346));
    ClkMux I__20908 (
            .O(N__86973),
            .I(N__86346));
    ClkMux I__20907 (
            .O(N__86972),
            .I(N__86346));
    ClkMux I__20906 (
            .O(N__86971),
            .I(N__86346));
    ClkMux I__20905 (
            .O(N__86970),
            .I(N__86346));
    ClkMux I__20904 (
            .O(N__86969),
            .I(N__86346));
    GlobalMux I__20903 (
            .O(N__86346),
            .I(N__86343));
    gio2CtrlBuf I__20902 (
            .O(N__86343),
            .I(clk_system_pll_g));
    CEMux I__20901 (
            .O(N__86340),
            .I(N__86333));
    CEMux I__20900 (
            .O(N__86339),
            .I(N__86330));
    CEMux I__20899 (
            .O(N__86338),
            .I(N__86326));
    CEMux I__20898 (
            .O(N__86337),
            .I(N__86323));
    CEMux I__20897 (
            .O(N__86336),
            .I(N__86320));
    LocalMux I__20896 (
            .O(N__86333),
            .I(N__86314));
    LocalMux I__20895 (
            .O(N__86330),
            .I(N__86311));
    CEMux I__20894 (
            .O(N__86329),
            .I(N__86308));
    LocalMux I__20893 (
            .O(N__86326),
            .I(N__86304));
    LocalMux I__20892 (
            .O(N__86323),
            .I(N__86299));
    LocalMux I__20891 (
            .O(N__86320),
            .I(N__86299));
    CEMux I__20890 (
            .O(N__86319),
            .I(N__86296));
    CEMux I__20889 (
            .O(N__86318),
            .I(N__86293));
    CEMux I__20888 (
            .O(N__86317),
            .I(N__86289));
    Span4Mux_h I__20887 (
            .O(N__86314),
            .I(N__86283));
    Span4Mux_h I__20886 (
            .O(N__86311),
            .I(N__86283));
    LocalMux I__20885 (
            .O(N__86308),
            .I(N__86280));
    CEMux I__20884 (
            .O(N__86307),
            .I(N__86277));
    Span4Mux_v I__20883 (
            .O(N__86304),
            .I(N__86269));
    Span4Mux_v I__20882 (
            .O(N__86299),
            .I(N__86269));
    LocalMux I__20881 (
            .O(N__86296),
            .I(N__86269));
    LocalMux I__20880 (
            .O(N__86293),
            .I(N__86266));
    CEMux I__20879 (
            .O(N__86292),
            .I(N__86263));
    LocalMux I__20878 (
            .O(N__86289),
            .I(N__86260));
    CEMux I__20877 (
            .O(N__86288),
            .I(N__86257));
    Span4Mux_h I__20876 (
            .O(N__86283),
            .I(N__86252));
    Span4Mux_h I__20875 (
            .O(N__86280),
            .I(N__86252));
    LocalMux I__20874 (
            .O(N__86277),
            .I(N__86249));
    CEMux I__20873 (
            .O(N__86276),
            .I(N__86246));
    Span4Mux_v I__20872 (
            .O(N__86269),
            .I(N__86243));
    Span4Mux_h I__20871 (
            .O(N__86266),
            .I(N__86240));
    LocalMux I__20870 (
            .O(N__86263),
            .I(N__86237));
    Span4Mux_h I__20869 (
            .O(N__86260),
            .I(N__86232));
    LocalMux I__20868 (
            .O(N__86257),
            .I(N__86232));
    Span4Mux_h I__20867 (
            .O(N__86252),
            .I(N__86225));
    Span4Mux_h I__20866 (
            .O(N__86249),
            .I(N__86225));
    LocalMux I__20865 (
            .O(N__86246),
            .I(N__86225));
    Span4Mux_h I__20864 (
            .O(N__86243),
            .I(N__86222));
    Span4Mux_h I__20863 (
            .O(N__86240),
            .I(N__86219));
    Span4Mux_v I__20862 (
            .O(N__86237),
            .I(N__86216));
    Span4Mux_h I__20861 (
            .O(N__86232),
            .I(N__86213));
    Span4Mux_v I__20860 (
            .O(N__86225),
            .I(N__86210));
    Span4Mux_h I__20859 (
            .O(N__86222),
            .I(N__86207));
    Span4Mux_h I__20858 (
            .O(N__86219),
            .I(N__86204));
    Span4Mux_v I__20857 (
            .O(N__86216),
            .I(N__86197));
    Span4Mux_h I__20856 (
            .O(N__86213),
            .I(N__86197));
    Span4Mux_h I__20855 (
            .O(N__86210),
            .I(N__86197));
    Odrv4 I__20854 (
            .O(N__86207),
            .I(\pid_front.N_789_0 ));
    Odrv4 I__20853 (
            .O(N__86204),
            .I(\pid_front.N_789_0 ));
    Odrv4 I__20852 (
            .O(N__86197),
            .I(\pid_front.N_789_0 ));
    InMux I__20851 (
            .O(N__86190),
            .I(N__86137));
    InMux I__20850 (
            .O(N__86189),
            .I(N__86137));
    InMux I__20849 (
            .O(N__86188),
            .I(N__86137));
    InMux I__20848 (
            .O(N__86187),
            .I(N__86137));
    InMux I__20847 (
            .O(N__86186),
            .I(N__86137));
    InMux I__20846 (
            .O(N__86185),
            .I(N__86134));
    InMux I__20845 (
            .O(N__86184),
            .I(N__86129));
    InMux I__20844 (
            .O(N__86183),
            .I(N__86129));
    InMux I__20843 (
            .O(N__86182),
            .I(N__86112));
    InMux I__20842 (
            .O(N__86181),
            .I(N__86112));
    InMux I__20841 (
            .O(N__86180),
            .I(N__86112));
    InMux I__20840 (
            .O(N__86179),
            .I(N__86112));
    InMux I__20839 (
            .O(N__86178),
            .I(N__86112));
    InMux I__20838 (
            .O(N__86177),
            .I(N__86112));
    InMux I__20837 (
            .O(N__86176),
            .I(N__86112));
    InMux I__20836 (
            .O(N__86175),
            .I(N__86112));
    InMux I__20835 (
            .O(N__86174),
            .I(N__86107));
    InMux I__20834 (
            .O(N__86173),
            .I(N__86107));
    InMux I__20833 (
            .O(N__86172),
            .I(N__86092));
    InMux I__20832 (
            .O(N__86171),
            .I(N__86092));
    InMux I__20831 (
            .O(N__86170),
            .I(N__86092));
    InMux I__20830 (
            .O(N__86169),
            .I(N__86092));
    InMux I__20829 (
            .O(N__86168),
            .I(N__86092));
    InMux I__20828 (
            .O(N__86167),
            .I(N__86092));
    InMux I__20827 (
            .O(N__86166),
            .I(N__86092));
    InMux I__20826 (
            .O(N__86165),
            .I(N__86089));
    InMux I__20825 (
            .O(N__86164),
            .I(N__86080));
    InMux I__20824 (
            .O(N__86163),
            .I(N__86080));
    InMux I__20823 (
            .O(N__86162),
            .I(N__86080));
    InMux I__20822 (
            .O(N__86161),
            .I(N__86080));
    InMux I__20821 (
            .O(N__86160),
            .I(N__86077));
    InMux I__20820 (
            .O(N__86159),
            .I(N__86072));
    InMux I__20819 (
            .O(N__86158),
            .I(N__86072));
    InMux I__20818 (
            .O(N__86157),
            .I(N__86069));
    InMux I__20817 (
            .O(N__86156),
            .I(N__86064));
    InMux I__20816 (
            .O(N__86155),
            .I(N__86064));
    InMux I__20815 (
            .O(N__86154),
            .I(N__86061));
    InMux I__20814 (
            .O(N__86153),
            .I(N__86058));
    InMux I__20813 (
            .O(N__86152),
            .I(N__86055));
    InMux I__20812 (
            .O(N__86151),
            .I(N__86052));
    InMux I__20811 (
            .O(N__86150),
            .I(N__86045));
    InMux I__20810 (
            .O(N__86149),
            .I(N__86045));
    InMux I__20809 (
            .O(N__86148),
            .I(N__86045));
    LocalMux I__20808 (
            .O(N__86137),
            .I(N__85999));
    LocalMux I__20807 (
            .O(N__86134),
            .I(N__85996));
    LocalMux I__20806 (
            .O(N__86129),
            .I(N__85993));
    LocalMux I__20805 (
            .O(N__86112),
            .I(N__85990));
    LocalMux I__20804 (
            .O(N__86107),
            .I(N__85987));
    LocalMux I__20803 (
            .O(N__86092),
            .I(N__85984));
    LocalMux I__20802 (
            .O(N__86089),
            .I(N__85981));
    LocalMux I__20801 (
            .O(N__86080),
            .I(N__85978));
    LocalMux I__20800 (
            .O(N__86077),
            .I(N__85975));
    LocalMux I__20799 (
            .O(N__86072),
            .I(N__85972));
    LocalMux I__20798 (
            .O(N__86069),
            .I(N__85969));
    LocalMux I__20797 (
            .O(N__86064),
            .I(N__85966));
    LocalMux I__20796 (
            .O(N__86061),
            .I(N__85963));
    LocalMux I__20795 (
            .O(N__86058),
            .I(N__85960));
    LocalMux I__20794 (
            .O(N__86055),
            .I(N__85957));
    LocalMux I__20793 (
            .O(N__86052),
            .I(N__85954));
    LocalMux I__20792 (
            .O(N__86045),
            .I(N__85951));
    SRMux I__20791 (
            .O(N__86044),
            .I(N__85830));
    SRMux I__20790 (
            .O(N__86043),
            .I(N__85830));
    SRMux I__20789 (
            .O(N__86042),
            .I(N__85830));
    SRMux I__20788 (
            .O(N__86041),
            .I(N__85830));
    SRMux I__20787 (
            .O(N__86040),
            .I(N__85830));
    SRMux I__20786 (
            .O(N__86039),
            .I(N__85830));
    SRMux I__20785 (
            .O(N__86038),
            .I(N__85830));
    SRMux I__20784 (
            .O(N__86037),
            .I(N__85830));
    SRMux I__20783 (
            .O(N__86036),
            .I(N__85830));
    SRMux I__20782 (
            .O(N__86035),
            .I(N__85830));
    SRMux I__20781 (
            .O(N__86034),
            .I(N__85830));
    SRMux I__20780 (
            .O(N__86033),
            .I(N__85830));
    SRMux I__20779 (
            .O(N__86032),
            .I(N__85830));
    SRMux I__20778 (
            .O(N__86031),
            .I(N__85830));
    SRMux I__20777 (
            .O(N__86030),
            .I(N__85830));
    SRMux I__20776 (
            .O(N__86029),
            .I(N__85830));
    SRMux I__20775 (
            .O(N__86028),
            .I(N__85830));
    SRMux I__20774 (
            .O(N__86027),
            .I(N__85830));
    SRMux I__20773 (
            .O(N__86026),
            .I(N__85830));
    SRMux I__20772 (
            .O(N__86025),
            .I(N__85830));
    SRMux I__20771 (
            .O(N__86024),
            .I(N__85830));
    SRMux I__20770 (
            .O(N__86023),
            .I(N__85830));
    SRMux I__20769 (
            .O(N__86022),
            .I(N__85830));
    SRMux I__20768 (
            .O(N__86021),
            .I(N__85830));
    SRMux I__20767 (
            .O(N__86020),
            .I(N__85830));
    SRMux I__20766 (
            .O(N__86019),
            .I(N__85830));
    SRMux I__20765 (
            .O(N__86018),
            .I(N__85830));
    SRMux I__20764 (
            .O(N__86017),
            .I(N__85830));
    SRMux I__20763 (
            .O(N__86016),
            .I(N__85830));
    SRMux I__20762 (
            .O(N__86015),
            .I(N__85830));
    SRMux I__20761 (
            .O(N__86014),
            .I(N__85830));
    SRMux I__20760 (
            .O(N__86013),
            .I(N__85830));
    SRMux I__20759 (
            .O(N__86012),
            .I(N__85830));
    SRMux I__20758 (
            .O(N__86011),
            .I(N__85830));
    SRMux I__20757 (
            .O(N__86010),
            .I(N__85830));
    SRMux I__20756 (
            .O(N__86009),
            .I(N__85830));
    SRMux I__20755 (
            .O(N__86008),
            .I(N__85830));
    SRMux I__20754 (
            .O(N__86007),
            .I(N__85830));
    SRMux I__20753 (
            .O(N__86006),
            .I(N__85830));
    SRMux I__20752 (
            .O(N__86005),
            .I(N__85830));
    SRMux I__20751 (
            .O(N__86004),
            .I(N__85830));
    SRMux I__20750 (
            .O(N__86003),
            .I(N__85830));
    SRMux I__20749 (
            .O(N__86002),
            .I(N__85830));
    Glb2LocalMux I__20748 (
            .O(N__85999),
            .I(N__85830));
    Glb2LocalMux I__20747 (
            .O(N__85996),
            .I(N__85830));
    Glb2LocalMux I__20746 (
            .O(N__85993),
            .I(N__85830));
    Glb2LocalMux I__20745 (
            .O(N__85990),
            .I(N__85830));
    Glb2LocalMux I__20744 (
            .O(N__85987),
            .I(N__85830));
    Glb2LocalMux I__20743 (
            .O(N__85984),
            .I(N__85830));
    Glb2LocalMux I__20742 (
            .O(N__85981),
            .I(N__85830));
    Glb2LocalMux I__20741 (
            .O(N__85978),
            .I(N__85830));
    Glb2LocalMux I__20740 (
            .O(N__85975),
            .I(N__85830));
    Glb2LocalMux I__20739 (
            .O(N__85972),
            .I(N__85830));
    Glb2LocalMux I__20738 (
            .O(N__85969),
            .I(N__85830));
    Glb2LocalMux I__20737 (
            .O(N__85966),
            .I(N__85830));
    Glb2LocalMux I__20736 (
            .O(N__85963),
            .I(N__85830));
    Glb2LocalMux I__20735 (
            .O(N__85960),
            .I(N__85830));
    Glb2LocalMux I__20734 (
            .O(N__85957),
            .I(N__85830));
    Glb2LocalMux I__20733 (
            .O(N__85954),
            .I(N__85830));
    Glb2LocalMux I__20732 (
            .O(N__85951),
            .I(N__85830));
    GlobalMux I__20731 (
            .O(N__85830),
            .I(N__85827));
    gio2CtrlBuf I__20730 (
            .O(N__85827),
            .I(N_940_g));
    InMux I__20729 (
            .O(N__85824),
            .I(N__85821));
    LocalMux I__20728 (
            .O(N__85821),
            .I(N__85818));
    Odrv4 I__20727 (
            .O(N__85818),
            .I(\pid_side.O_1_16 ));
    InMux I__20726 (
            .O(N__85815),
            .I(N__85812));
    LocalMux I__20725 (
            .O(N__85812),
            .I(N__85806));
    InMux I__20724 (
            .O(N__85811),
            .I(N__85799));
    InMux I__20723 (
            .O(N__85810),
            .I(N__85799));
    InMux I__20722 (
            .O(N__85809),
            .I(N__85799));
    Span4Mux_h I__20721 (
            .O(N__85806),
            .I(N__85795));
    LocalMux I__20720 (
            .O(N__85799),
            .I(N__85792));
    InMux I__20719 (
            .O(N__85798),
            .I(N__85789));
    Odrv4 I__20718 (
            .O(N__85795),
            .I(\pid_side.error_d_regZ0Z_14 ));
    Odrv12 I__20717 (
            .O(N__85792),
            .I(\pid_side.error_d_regZ0Z_14 ));
    LocalMux I__20716 (
            .O(N__85789),
            .I(\pid_side.error_d_regZ0Z_14 ));
    InMux I__20715 (
            .O(N__85782),
            .I(N__85779));
    LocalMux I__20714 (
            .O(N__85779),
            .I(N__85776));
    Odrv4 I__20713 (
            .O(N__85776),
            .I(\pid_side.O_1_18 ));
    InMux I__20712 (
            .O(N__85773),
            .I(N__85767));
    InMux I__20711 (
            .O(N__85772),
            .I(N__85767));
    LocalMux I__20710 (
            .O(N__85767),
            .I(N__85763));
    InMux I__20709 (
            .O(N__85766),
            .I(N__85760));
    Odrv4 I__20708 (
            .O(N__85763),
            .I(\pid_side.error_d_regZ0Z_16 ));
    LocalMux I__20707 (
            .O(N__85760),
            .I(\pid_side.error_d_regZ0Z_16 ));
    CEMux I__20706 (
            .O(N__85755),
            .I(N__85748));
    CEMux I__20705 (
            .O(N__85754),
            .I(N__85742));
    CEMux I__20704 (
            .O(N__85753),
            .I(N__85738));
    CEMux I__20703 (
            .O(N__85752),
            .I(N__85735));
    CEMux I__20702 (
            .O(N__85751),
            .I(N__85732));
    LocalMux I__20701 (
            .O(N__85748),
            .I(N__85729));
    CEMux I__20700 (
            .O(N__85747),
            .I(N__85725));
    CEMux I__20699 (
            .O(N__85746),
            .I(N__85720));
    CEMux I__20698 (
            .O(N__85745),
            .I(N__85717));
    LocalMux I__20697 (
            .O(N__85742),
            .I(N__85714));
    CEMux I__20696 (
            .O(N__85741),
            .I(N__85711));
    LocalMux I__20695 (
            .O(N__85738),
            .I(N__85705));
    LocalMux I__20694 (
            .O(N__85735),
            .I(N__85702));
    LocalMux I__20693 (
            .O(N__85732),
            .I(N__85699));
    Span4Mux_s2_h I__20692 (
            .O(N__85729),
            .I(N__85696));
    CEMux I__20691 (
            .O(N__85728),
            .I(N__85693));
    LocalMux I__20690 (
            .O(N__85725),
            .I(N__85690));
    CEMux I__20689 (
            .O(N__85724),
            .I(N__85687));
    CEMux I__20688 (
            .O(N__85723),
            .I(N__85684));
    LocalMux I__20687 (
            .O(N__85720),
            .I(N__85681));
    LocalMux I__20686 (
            .O(N__85717),
            .I(N__85676));
    Span4Mux_h I__20685 (
            .O(N__85714),
            .I(N__85676));
    LocalMux I__20684 (
            .O(N__85711),
            .I(N__85673));
    CEMux I__20683 (
            .O(N__85710),
            .I(N__85670));
    CEMux I__20682 (
            .O(N__85709),
            .I(N__85667));
    CEMux I__20681 (
            .O(N__85708),
            .I(N__85664));
    Span4Mux_v I__20680 (
            .O(N__85705),
            .I(N__85657));
    Span4Mux_v I__20679 (
            .O(N__85702),
            .I(N__85657));
    Span4Mux_v I__20678 (
            .O(N__85699),
            .I(N__85657));
    Span4Mux_h I__20677 (
            .O(N__85696),
            .I(N__85652));
    LocalMux I__20676 (
            .O(N__85693),
            .I(N__85652));
    Sp12to4 I__20675 (
            .O(N__85690),
            .I(N__85647));
    LocalMux I__20674 (
            .O(N__85687),
            .I(N__85647));
    LocalMux I__20673 (
            .O(N__85684),
            .I(N__85644));
    Span4Mux_h I__20672 (
            .O(N__85681),
            .I(N__85631));
    Span4Mux_s3_h I__20671 (
            .O(N__85676),
            .I(N__85631));
    Span4Mux_s3_h I__20670 (
            .O(N__85673),
            .I(N__85631));
    LocalMux I__20669 (
            .O(N__85670),
            .I(N__85631));
    LocalMux I__20668 (
            .O(N__85667),
            .I(N__85631));
    LocalMux I__20667 (
            .O(N__85664),
            .I(N__85631));
    Odrv4 I__20666 (
            .O(N__85657),
            .I(\pid_side.N_873_0 ));
    Odrv4 I__20665 (
            .O(N__85652),
            .I(\pid_side.N_873_0 ));
    Odrv12 I__20664 (
            .O(N__85647),
            .I(\pid_side.N_873_0 ));
    Odrv12 I__20663 (
            .O(N__85644),
            .I(\pid_side.N_873_0 ));
    Odrv4 I__20662 (
            .O(N__85631),
            .I(\pid_side.N_873_0 ));
    InMux I__20661 (
            .O(N__85620),
            .I(N__85617));
    LocalMux I__20660 (
            .O(N__85617),
            .I(N__85614));
    Odrv4 I__20659 (
            .O(N__85614),
            .I(\pid_side.N_5 ));
    InMux I__20658 (
            .O(N__85611),
            .I(N__85605));
    InMux I__20657 (
            .O(N__85610),
            .I(N__85602));
    InMux I__20656 (
            .O(N__85609),
            .I(N__85597));
    InMux I__20655 (
            .O(N__85608),
            .I(N__85597));
    LocalMux I__20654 (
            .O(N__85605),
            .I(N__85594));
    LocalMux I__20653 (
            .O(N__85602),
            .I(N__85587));
    LocalMux I__20652 (
            .O(N__85597),
            .I(N__85587));
    Span4Mux_v I__20651 (
            .O(N__85594),
            .I(N__85582));
    InMux I__20650 (
            .O(N__85593),
            .I(N__85577));
    InMux I__20649 (
            .O(N__85592),
            .I(N__85577));
    Span4Mux_h I__20648 (
            .O(N__85587),
            .I(N__85574));
    InMux I__20647 (
            .O(N__85586),
            .I(N__85571));
    InMux I__20646 (
            .O(N__85585),
            .I(N__85568));
    Odrv4 I__20645 (
            .O(N__85582),
            .I(\pid_side.error_d_regZ0Z_13 ));
    LocalMux I__20644 (
            .O(N__85577),
            .I(\pid_side.error_d_regZ0Z_13 ));
    Odrv4 I__20643 (
            .O(N__85574),
            .I(\pid_side.error_d_regZ0Z_13 ));
    LocalMux I__20642 (
            .O(N__85571),
            .I(\pid_side.error_d_regZ0Z_13 ));
    LocalMux I__20641 (
            .O(N__85568),
            .I(\pid_side.error_d_regZ0Z_13 ));
    CascadeMux I__20640 (
            .O(N__85557),
            .I(N__85553));
    CascadeMux I__20639 (
            .O(N__85556),
            .I(N__85549));
    InMux I__20638 (
            .O(N__85553),
            .I(N__85543));
    InMux I__20637 (
            .O(N__85552),
            .I(N__85543));
    InMux I__20636 (
            .O(N__85549),
            .I(N__85538));
    InMux I__20635 (
            .O(N__85548),
            .I(N__85538));
    LocalMux I__20634 (
            .O(N__85543),
            .I(N__85534));
    LocalMux I__20633 (
            .O(N__85538),
            .I(N__85531));
    InMux I__20632 (
            .O(N__85537),
            .I(N__85526));
    Span4Mux_s1_h I__20631 (
            .O(N__85534),
            .I(N__85521));
    Span4Mux_v I__20630 (
            .O(N__85531),
            .I(N__85521));
    InMux I__20629 (
            .O(N__85530),
            .I(N__85518));
    InMux I__20628 (
            .O(N__85529),
            .I(N__85515));
    LocalMux I__20627 (
            .O(N__85526),
            .I(\pid_side.error_d_reg_prevZ0Z_13 ));
    Odrv4 I__20626 (
            .O(N__85521),
            .I(\pid_side.error_d_reg_prevZ0Z_13 ));
    LocalMux I__20625 (
            .O(N__85518),
            .I(\pid_side.error_d_reg_prevZ0Z_13 ));
    LocalMux I__20624 (
            .O(N__85515),
            .I(\pid_side.error_d_reg_prevZ0Z_13 ));
    InMux I__20623 (
            .O(N__85506),
            .I(N__85500));
    InMux I__20622 (
            .O(N__85505),
            .I(N__85495));
    InMux I__20621 (
            .O(N__85504),
            .I(N__85495));
    CascadeMux I__20620 (
            .O(N__85503),
            .I(N__85492));
    LocalMux I__20619 (
            .O(N__85500),
            .I(N__85486));
    LocalMux I__20618 (
            .O(N__85495),
            .I(N__85483));
    InMux I__20617 (
            .O(N__85492),
            .I(N__85480));
    InMux I__20616 (
            .O(N__85491),
            .I(N__85475));
    InMux I__20615 (
            .O(N__85490),
            .I(N__85475));
    InMux I__20614 (
            .O(N__85489),
            .I(N__85472));
    Span4Mux_v I__20613 (
            .O(N__85486),
            .I(N__85469));
    Span4Mux_v I__20612 (
            .O(N__85483),
            .I(N__85466));
    LocalMux I__20611 (
            .O(N__85480),
            .I(N__85463));
    LocalMux I__20610 (
            .O(N__85475),
            .I(N__85458));
    LocalMux I__20609 (
            .O(N__85472),
            .I(N__85458));
    Span4Mux_h I__20608 (
            .O(N__85469),
            .I(N__85455));
    Span4Mux_h I__20607 (
            .O(N__85466),
            .I(N__85448));
    Span4Mux_v I__20606 (
            .O(N__85463),
            .I(N__85448));
    Span4Mux_v I__20605 (
            .O(N__85458),
            .I(N__85448));
    Odrv4 I__20604 (
            .O(N__85455),
            .I(\pid_side.error_p_regZ0Z_13 ));
    Odrv4 I__20603 (
            .O(N__85448),
            .I(\pid_side.error_p_regZ0Z_13 ));
    InMux I__20602 (
            .O(N__85443),
            .I(N__85440));
    LocalMux I__20601 (
            .O(N__85440),
            .I(N__85437));
    Odrv12 I__20600 (
            .O(N__85437),
            .I(\pid_side.error_d_reg_prev_esr_RNI2OIO_1Z0Z_13 ));
    InMux I__20599 (
            .O(N__85434),
            .I(N__85431));
    LocalMux I__20598 (
            .O(N__85431),
            .I(N__85428));
    Span4Mux_v I__20597 (
            .O(N__85428),
            .I(N__85425));
    Odrv4 I__20596 (
            .O(N__85425),
            .I(\pid_front.O_4 ));
    InMux I__20595 (
            .O(N__85422),
            .I(N__85413));
    InMux I__20594 (
            .O(N__85421),
            .I(N__85413));
    InMux I__20593 (
            .O(N__85420),
            .I(N__85413));
    LocalMux I__20592 (
            .O(N__85413),
            .I(N__85410));
    Span12Mux_h I__20591 (
            .O(N__85410),
            .I(N__85407));
    Odrv12 I__20590 (
            .O(N__85407),
            .I(\pid_front.error_d_regZ0Z_2 ));
    InMux I__20589 (
            .O(N__85404),
            .I(N__85401));
    LocalMux I__20588 (
            .O(N__85401),
            .I(N__85397));
    InMux I__20587 (
            .O(N__85400),
            .I(N__85393));
    Span4Mux_v I__20586 (
            .O(N__85397),
            .I(N__85390));
    InMux I__20585 (
            .O(N__85396),
            .I(N__85387));
    LocalMux I__20584 (
            .O(N__85393),
            .I(N__85384));
    Span4Mux_h I__20583 (
            .O(N__85390),
            .I(N__85381));
    LocalMux I__20582 (
            .O(N__85387),
            .I(N__85375));
    Span4Mux_v I__20581 (
            .O(N__85384),
            .I(N__85371));
    Span4Mux_h I__20580 (
            .O(N__85381),
            .I(N__85368));
    InMux I__20579 (
            .O(N__85380),
            .I(N__85365));
    InMux I__20578 (
            .O(N__85379),
            .I(N__85358));
    CascadeMux I__20577 (
            .O(N__85378),
            .I(N__85353));
    Span4Mux_v I__20576 (
            .O(N__85375),
            .I(N__85350));
    InMux I__20575 (
            .O(N__85374),
            .I(N__85347));
    Span4Mux_v I__20574 (
            .O(N__85371),
            .I(N__85340));
    Span4Mux_h I__20573 (
            .O(N__85368),
            .I(N__85340));
    LocalMux I__20572 (
            .O(N__85365),
            .I(N__85340));
    InMux I__20571 (
            .O(N__85364),
            .I(N__85337));
    InMux I__20570 (
            .O(N__85363),
            .I(N__85334));
    InMux I__20569 (
            .O(N__85362),
            .I(N__85331));
    InMux I__20568 (
            .O(N__85361),
            .I(N__85328));
    LocalMux I__20567 (
            .O(N__85358),
            .I(N__85325));
    InMux I__20566 (
            .O(N__85357),
            .I(N__85322));
    InMux I__20565 (
            .O(N__85356),
            .I(N__85318));
    InMux I__20564 (
            .O(N__85353),
            .I(N__85315));
    Span4Mux_h I__20563 (
            .O(N__85350),
            .I(N__85312));
    LocalMux I__20562 (
            .O(N__85347),
            .I(N__85309));
    Span4Mux_h I__20561 (
            .O(N__85340),
            .I(N__85305));
    LocalMux I__20560 (
            .O(N__85337),
            .I(N__85302));
    LocalMux I__20559 (
            .O(N__85334),
            .I(N__85295));
    LocalMux I__20558 (
            .O(N__85331),
            .I(N__85295));
    LocalMux I__20557 (
            .O(N__85328),
            .I(N__85295));
    Span4Mux_h I__20556 (
            .O(N__85325),
            .I(N__85292));
    LocalMux I__20555 (
            .O(N__85322),
            .I(N__85289));
    CascadeMux I__20554 (
            .O(N__85321),
            .I(N__85285));
    LocalMux I__20553 (
            .O(N__85318),
            .I(N__85280));
    LocalMux I__20552 (
            .O(N__85315),
            .I(N__85280));
    Sp12to4 I__20551 (
            .O(N__85312),
            .I(N__85277));
    Span12Mux_h I__20550 (
            .O(N__85309),
            .I(N__85274));
    InMux I__20549 (
            .O(N__85308),
            .I(N__85271));
    Span4Mux_h I__20548 (
            .O(N__85305),
            .I(N__85268));
    Span4Mux_h I__20547 (
            .O(N__85302),
            .I(N__85259));
    Span4Mux_v I__20546 (
            .O(N__85295),
            .I(N__85259));
    Span4Mux_v I__20545 (
            .O(N__85292),
            .I(N__85259));
    Span4Mux_h I__20544 (
            .O(N__85289),
            .I(N__85259));
    InMux I__20543 (
            .O(N__85288),
            .I(N__85254));
    InMux I__20542 (
            .O(N__85285),
            .I(N__85254));
    Span4Mux_h I__20541 (
            .O(N__85280),
            .I(N__85251));
    Odrv12 I__20540 (
            .O(N__85277),
            .I(uart_pc_data_7));
    Odrv12 I__20539 (
            .O(N__85274),
            .I(uart_pc_data_7));
    LocalMux I__20538 (
            .O(N__85271),
            .I(uart_pc_data_7));
    Odrv4 I__20537 (
            .O(N__85268),
            .I(uart_pc_data_7));
    Odrv4 I__20536 (
            .O(N__85259),
            .I(uart_pc_data_7));
    LocalMux I__20535 (
            .O(N__85254),
            .I(uart_pc_data_7));
    Odrv4 I__20534 (
            .O(N__85251),
            .I(uart_pc_data_7));
    InMux I__20533 (
            .O(N__85236),
            .I(N__85233));
    LocalMux I__20532 (
            .O(N__85233),
            .I(N__85229));
    InMux I__20531 (
            .O(N__85232),
            .I(N__85226));
    Span4Mux_v I__20530 (
            .O(N__85229),
            .I(N__85223));
    LocalMux I__20529 (
            .O(N__85226),
            .I(N__85220));
    Odrv4 I__20528 (
            .O(N__85223),
            .I(xy_kd_7));
    Odrv4 I__20527 (
            .O(N__85220),
            .I(xy_kd_7));
    InMux I__20526 (
            .O(N__85215),
            .I(N__85211));
    InMux I__20525 (
            .O(N__85214),
            .I(N__85206));
    LocalMux I__20524 (
            .O(N__85211),
            .I(N__85203));
    InMux I__20523 (
            .O(N__85210),
            .I(N__85200));
    InMux I__20522 (
            .O(N__85209),
            .I(N__85195));
    LocalMux I__20521 (
            .O(N__85206),
            .I(N__85192));
    Span4Mux_v I__20520 (
            .O(N__85203),
            .I(N__85189));
    LocalMux I__20519 (
            .O(N__85200),
            .I(N__85184));
    InMux I__20518 (
            .O(N__85199),
            .I(N__85181));
    InMux I__20517 (
            .O(N__85198),
            .I(N__85178));
    LocalMux I__20516 (
            .O(N__85195),
            .I(N__85174));
    Span4Mux_h I__20515 (
            .O(N__85192),
            .I(N__85169));
    Span4Mux_h I__20514 (
            .O(N__85189),
            .I(N__85169));
    InMux I__20513 (
            .O(N__85188),
            .I(N__85165));
    InMux I__20512 (
            .O(N__85187),
            .I(N__85162));
    Span4Mux_h I__20511 (
            .O(N__85184),
            .I(N__85159));
    LocalMux I__20510 (
            .O(N__85181),
            .I(N__85155));
    LocalMux I__20509 (
            .O(N__85178),
            .I(N__85152));
    InMux I__20508 (
            .O(N__85177),
            .I(N__85149));
    Span4Mux_v I__20507 (
            .O(N__85174),
            .I(N__85146));
    Span4Mux_v I__20506 (
            .O(N__85169),
            .I(N__85143));
    InMux I__20505 (
            .O(N__85168),
            .I(N__85140));
    LocalMux I__20504 (
            .O(N__85165),
            .I(N__85133));
    LocalMux I__20503 (
            .O(N__85162),
            .I(N__85133));
    Span4Mux_h I__20502 (
            .O(N__85159),
            .I(N__85133));
    InMux I__20501 (
            .O(N__85158),
            .I(N__85127));
    Span4Mux_v I__20500 (
            .O(N__85155),
            .I(N__85122));
    Span4Mux_v I__20499 (
            .O(N__85152),
            .I(N__85122));
    LocalMux I__20498 (
            .O(N__85149),
            .I(N__85119));
    Span4Mux_v I__20497 (
            .O(N__85146),
            .I(N__85116));
    Sp12to4 I__20496 (
            .O(N__85143),
            .I(N__85113));
    LocalMux I__20495 (
            .O(N__85140),
            .I(N__85110));
    Span4Mux_v I__20494 (
            .O(N__85133),
            .I(N__85107));
    InMux I__20493 (
            .O(N__85132),
            .I(N__85104));
    InMux I__20492 (
            .O(N__85131),
            .I(N__85099));
    InMux I__20491 (
            .O(N__85130),
            .I(N__85099));
    LocalMux I__20490 (
            .O(N__85127),
            .I(N__85086));
    Sp12to4 I__20489 (
            .O(N__85122),
            .I(N__85086));
    Span12Mux_s11_v I__20488 (
            .O(N__85119),
            .I(N__85086));
    Sp12to4 I__20487 (
            .O(N__85116),
            .I(N__85086));
    Span12Mux_s11_h I__20486 (
            .O(N__85113),
            .I(N__85086));
    Span4Mux_v I__20485 (
            .O(N__85110),
            .I(N__85079));
    Span4Mux_v I__20484 (
            .O(N__85107),
            .I(N__85079));
    LocalMux I__20483 (
            .O(N__85104),
            .I(N__85079));
    LocalMux I__20482 (
            .O(N__85099),
            .I(N__85076));
    InMux I__20481 (
            .O(N__85098),
            .I(N__85071));
    InMux I__20480 (
            .O(N__85097),
            .I(N__85071));
    Odrv12 I__20479 (
            .O(N__85086),
            .I(uart_pc_data_5));
    Odrv4 I__20478 (
            .O(N__85079),
            .I(uart_pc_data_5));
    Odrv4 I__20477 (
            .O(N__85076),
            .I(uart_pc_data_5));
    LocalMux I__20476 (
            .O(N__85071),
            .I(uart_pc_data_5));
    InMux I__20475 (
            .O(N__85062),
            .I(N__85058));
    InMux I__20474 (
            .O(N__85061),
            .I(N__85055));
    LocalMux I__20473 (
            .O(N__85058),
            .I(N__85052));
    LocalMux I__20472 (
            .O(N__85055),
            .I(N__85049));
    Span4Mux_v I__20471 (
            .O(N__85052),
            .I(N__85044));
    Span4Mux_s0_h I__20470 (
            .O(N__85049),
            .I(N__85044));
    Odrv4 I__20469 (
            .O(N__85044),
            .I(xy_kd_5));
    InMux I__20468 (
            .O(N__85041),
            .I(N__85036));
    InMux I__20467 (
            .O(N__85040),
            .I(N__85033));
    InMux I__20466 (
            .O(N__85039),
            .I(N__85030));
    LocalMux I__20465 (
            .O(N__85036),
            .I(N__85023));
    LocalMux I__20464 (
            .O(N__85033),
            .I(N__85020));
    LocalMux I__20463 (
            .O(N__85030),
            .I(N__85016));
    CascadeMux I__20462 (
            .O(N__85029),
            .I(N__85013));
    InMux I__20461 (
            .O(N__85028),
            .I(N__85010));
    InMux I__20460 (
            .O(N__85027),
            .I(N__85006));
    InMux I__20459 (
            .O(N__85026),
            .I(N__85003));
    Span4Mux_v I__20458 (
            .O(N__85023),
            .I(N__85000));
    Span4Mux_v I__20457 (
            .O(N__85020),
            .I(N__84997));
    InMux I__20456 (
            .O(N__85019),
            .I(N__84994));
    Span4Mux_v I__20455 (
            .O(N__85016),
            .I(N__84991));
    InMux I__20454 (
            .O(N__85013),
            .I(N__84988));
    LocalMux I__20453 (
            .O(N__85010),
            .I(N__84984));
    InMux I__20452 (
            .O(N__85009),
            .I(N__84980));
    LocalMux I__20451 (
            .O(N__85006),
            .I(N__84974));
    LocalMux I__20450 (
            .O(N__85003),
            .I(N__84974));
    Span4Mux_v I__20449 (
            .O(N__85000),
            .I(N__84971));
    Span4Mux_v I__20448 (
            .O(N__84997),
            .I(N__84968));
    LocalMux I__20447 (
            .O(N__84994),
            .I(N__84961));
    Span4Mux_v I__20446 (
            .O(N__84991),
            .I(N__84961));
    LocalMux I__20445 (
            .O(N__84988),
            .I(N__84961));
    InMux I__20444 (
            .O(N__84987),
            .I(N__84957));
    Span12Mux_v I__20443 (
            .O(N__84984),
            .I(N__84954));
    InMux I__20442 (
            .O(N__84983),
            .I(N__84951));
    LocalMux I__20441 (
            .O(N__84980),
            .I(N__84948));
    InMux I__20440 (
            .O(N__84979),
            .I(N__84945));
    Span4Mux_v I__20439 (
            .O(N__84974),
            .I(N__84940));
    Span4Mux_v I__20438 (
            .O(N__84971),
            .I(N__84940));
    Sp12to4 I__20437 (
            .O(N__84968),
            .I(N__84937));
    Span4Mux_v I__20436 (
            .O(N__84961),
            .I(N__84933));
    InMux I__20435 (
            .O(N__84960),
            .I(N__84930));
    LocalMux I__20434 (
            .O(N__84957),
            .I(N__84927));
    Span12Mux_h I__20433 (
            .O(N__84954),
            .I(N__84924));
    LocalMux I__20432 (
            .O(N__84951),
            .I(N__84913));
    Span12Mux_s10_v I__20431 (
            .O(N__84948),
            .I(N__84913));
    LocalMux I__20430 (
            .O(N__84945),
            .I(N__84913));
    Sp12to4 I__20429 (
            .O(N__84940),
            .I(N__84913));
    Span12Mux_s11_h I__20428 (
            .O(N__84937),
            .I(N__84913));
    InMux I__20427 (
            .O(N__84936),
            .I(N__84910));
    Span4Mux_v I__20426 (
            .O(N__84933),
            .I(N__84907));
    LocalMux I__20425 (
            .O(N__84930),
            .I(uart_pc_data_4));
    Odrv4 I__20424 (
            .O(N__84927),
            .I(uart_pc_data_4));
    Odrv12 I__20423 (
            .O(N__84924),
            .I(uart_pc_data_4));
    Odrv12 I__20422 (
            .O(N__84913),
            .I(uart_pc_data_4));
    LocalMux I__20421 (
            .O(N__84910),
            .I(uart_pc_data_4));
    Odrv4 I__20420 (
            .O(N__84907),
            .I(uart_pc_data_4));
    InMux I__20419 (
            .O(N__84894),
            .I(N__84890));
    InMux I__20418 (
            .O(N__84893),
            .I(N__84887));
    LocalMux I__20417 (
            .O(N__84890),
            .I(N__84884));
    LocalMux I__20416 (
            .O(N__84887),
            .I(N__84881));
    Span4Mux_v I__20415 (
            .O(N__84884),
            .I(N__84876));
    Span4Mux_s0_h I__20414 (
            .O(N__84881),
            .I(N__84876));
    Odrv4 I__20413 (
            .O(N__84876),
            .I(xy_kd_4));
    CEMux I__20412 (
            .O(N__84873),
            .I(N__84870));
    LocalMux I__20411 (
            .O(N__84870),
            .I(N__84863));
    CEMux I__20410 (
            .O(N__84869),
            .I(N__84860));
    CEMux I__20409 (
            .O(N__84868),
            .I(N__84857));
    CEMux I__20408 (
            .O(N__84867),
            .I(N__84854));
    CEMux I__20407 (
            .O(N__84866),
            .I(N__84851));
    Span4Mux_v I__20406 (
            .O(N__84863),
            .I(N__84846));
    LocalMux I__20405 (
            .O(N__84860),
            .I(N__84846));
    LocalMux I__20404 (
            .O(N__84857),
            .I(N__84839));
    LocalMux I__20403 (
            .O(N__84854),
            .I(N__84839));
    LocalMux I__20402 (
            .O(N__84851),
            .I(N__84839));
    Span4Mux_v I__20401 (
            .O(N__84846),
            .I(N__84834));
    Span4Mux_v I__20400 (
            .O(N__84839),
            .I(N__84834));
    Span4Mux_v I__20399 (
            .O(N__84834),
            .I(N__84831));
    Sp12to4 I__20398 (
            .O(N__84831),
            .I(N__84827));
    CEMux I__20397 (
            .O(N__84830),
            .I(N__84824));
    Span12Mux_h I__20396 (
            .O(N__84827),
            .I(N__84819));
    LocalMux I__20395 (
            .O(N__84824),
            .I(N__84819));
    Span12Mux_v I__20394 (
            .O(N__84819),
            .I(N__84816));
    Odrv12 I__20393 (
            .O(N__84816),
            .I(\Commands_frame_decoder.state_RNITUI31Z0Z_13 ));
    InMux I__20392 (
            .O(N__84813),
            .I(N__84810));
    LocalMux I__20391 (
            .O(N__84810),
            .I(\pid_side.O_2_15 ));
    CascadeMux I__20390 (
            .O(N__84807),
            .I(N__84801));
    InMux I__20389 (
            .O(N__84806),
            .I(N__84793));
    InMux I__20388 (
            .O(N__84805),
            .I(N__84793));
    InMux I__20387 (
            .O(N__84804),
            .I(N__84788));
    InMux I__20386 (
            .O(N__84801),
            .I(N__84788));
    InMux I__20385 (
            .O(N__84800),
            .I(N__84785));
    InMux I__20384 (
            .O(N__84799),
            .I(N__84780));
    InMux I__20383 (
            .O(N__84798),
            .I(N__84780));
    LocalMux I__20382 (
            .O(N__84793),
            .I(N__84775));
    LocalMux I__20381 (
            .O(N__84788),
            .I(N__84775));
    LocalMux I__20380 (
            .O(N__84785),
            .I(N__84772));
    LocalMux I__20379 (
            .O(N__84780),
            .I(N__84769));
    Span4Mux_h I__20378 (
            .O(N__84775),
            .I(N__84766));
    Span12Mux_v I__20377 (
            .O(N__84772),
            .I(N__84763));
    Span4Mux_v I__20376 (
            .O(N__84769),
            .I(N__84760));
    Span4Mux_v I__20375 (
            .O(N__84766),
            .I(N__84757));
    Odrv12 I__20374 (
            .O(N__84763),
            .I(\pid_side.error_p_regZ0Z_12 ));
    Odrv4 I__20373 (
            .O(N__84760),
            .I(\pid_side.error_p_regZ0Z_12 ));
    Odrv4 I__20372 (
            .O(N__84757),
            .I(\pid_side.error_p_regZ0Z_12 ));
    InMux I__20371 (
            .O(N__84750),
            .I(N__84747));
    LocalMux I__20370 (
            .O(N__84747),
            .I(N__84744));
    Span4Mux_h I__20369 (
            .O(N__84744),
            .I(N__84741));
    Odrv4 I__20368 (
            .O(N__84741),
            .I(\pid_side.O_1_19 ));
    InMux I__20367 (
            .O(N__84738),
            .I(N__84729));
    InMux I__20366 (
            .O(N__84737),
            .I(N__84729));
    InMux I__20365 (
            .O(N__84736),
            .I(N__84729));
    LocalMux I__20364 (
            .O(N__84729),
            .I(\pid_side.error_d_regZ0Z_17 ));
    InMux I__20363 (
            .O(N__84726),
            .I(N__84723));
    LocalMux I__20362 (
            .O(N__84723),
            .I(N__84720));
    Odrv4 I__20361 (
            .O(N__84720),
            .I(\pid_side.O_1_20 ));
    InMux I__20360 (
            .O(N__84717),
            .I(N__84708));
    InMux I__20359 (
            .O(N__84716),
            .I(N__84708));
    InMux I__20358 (
            .O(N__84715),
            .I(N__84708));
    LocalMux I__20357 (
            .O(N__84708),
            .I(\pid_side.error_d_regZ0Z_18 ));
    InMux I__20356 (
            .O(N__84705),
            .I(N__84702));
    LocalMux I__20355 (
            .O(N__84702),
            .I(N__84699));
    Span4Mux_v I__20354 (
            .O(N__84699),
            .I(N__84696));
    Odrv4 I__20353 (
            .O(N__84696),
            .I(\pid_side.O_1_21 ));
    InMux I__20352 (
            .O(N__84693),
            .I(N__84684));
    InMux I__20351 (
            .O(N__84692),
            .I(N__84684));
    InMux I__20350 (
            .O(N__84691),
            .I(N__84684));
    LocalMux I__20349 (
            .O(N__84684),
            .I(N__84681));
    Odrv4 I__20348 (
            .O(N__84681),
            .I(\pid_side.error_d_regZ0Z_19 ));
    InMux I__20347 (
            .O(N__84678),
            .I(N__84675));
    LocalMux I__20346 (
            .O(N__84675),
            .I(N__84672));
    Span4Mux_v I__20345 (
            .O(N__84672),
            .I(N__84669));
    Odrv4 I__20344 (
            .O(N__84669),
            .I(\pid_side.O_1_23 ));
    InMux I__20343 (
            .O(N__84666),
            .I(N__84657));
    InMux I__20342 (
            .O(N__84665),
            .I(N__84657));
    InMux I__20341 (
            .O(N__84664),
            .I(N__84657));
    LocalMux I__20340 (
            .O(N__84657),
            .I(N__84654));
    Span4Mux_h I__20339 (
            .O(N__84654),
            .I(N__84651));
    Span4Mux_h I__20338 (
            .O(N__84651),
            .I(N__84648));
    Odrv4 I__20337 (
            .O(N__84648),
            .I(\pid_side.error_d_regZ0Z_21 ));
    InMux I__20336 (
            .O(N__84645),
            .I(N__84642));
    LocalMux I__20335 (
            .O(N__84642),
            .I(N__84639));
    Span4Mux_v I__20334 (
            .O(N__84639),
            .I(N__84636));
    Odrv4 I__20333 (
            .O(N__84636),
            .I(\pid_side.O_1_24 ));
    CascadeMux I__20332 (
            .O(N__84633),
            .I(N__84626));
    InMux I__20331 (
            .O(N__84632),
            .I(N__84614));
    InMux I__20330 (
            .O(N__84631),
            .I(N__84614));
    InMux I__20329 (
            .O(N__84630),
            .I(N__84614));
    InMux I__20328 (
            .O(N__84629),
            .I(N__84605));
    InMux I__20327 (
            .O(N__84626),
            .I(N__84605));
    InMux I__20326 (
            .O(N__84625),
            .I(N__84605));
    InMux I__20325 (
            .O(N__84624),
            .I(N__84605));
    InMux I__20324 (
            .O(N__84623),
            .I(N__84598));
    InMux I__20323 (
            .O(N__84622),
            .I(N__84598));
    InMux I__20322 (
            .O(N__84621),
            .I(N__84598));
    LocalMux I__20321 (
            .O(N__84614),
            .I(N__84595));
    LocalMux I__20320 (
            .O(N__84605),
            .I(N__84588));
    LocalMux I__20319 (
            .O(N__84598),
            .I(N__84585));
    Span4Mux_h I__20318 (
            .O(N__84595),
            .I(N__84582));
    InMux I__20317 (
            .O(N__84594),
            .I(N__84573));
    InMux I__20316 (
            .O(N__84593),
            .I(N__84573));
    InMux I__20315 (
            .O(N__84592),
            .I(N__84573));
    InMux I__20314 (
            .O(N__84591),
            .I(N__84573));
    Span4Mux_h I__20313 (
            .O(N__84588),
            .I(N__84570));
    Span4Mux_h I__20312 (
            .O(N__84585),
            .I(N__84567));
    Span4Mux_h I__20311 (
            .O(N__84582),
            .I(N__84564));
    LocalMux I__20310 (
            .O(N__84573),
            .I(N__84561));
    Span4Mux_h I__20309 (
            .O(N__84570),
            .I(N__84558));
    Span4Mux_h I__20308 (
            .O(N__84567),
            .I(N__84555));
    Odrv4 I__20307 (
            .O(N__84564),
            .I(\pid_side.error_d_regZ0Z_22 ));
    Odrv12 I__20306 (
            .O(N__84561),
            .I(\pid_side.error_d_regZ0Z_22 ));
    Odrv4 I__20305 (
            .O(N__84558),
            .I(\pid_side.error_d_regZ0Z_22 ));
    Odrv4 I__20304 (
            .O(N__84555),
            .I(\pid_side.error_d_regZ0Z_22 ));
    InMux I__20303 (
            .O(N__84546),
            .I(N__84543));
    LocalMux I__20302 (
            .O(N__84543),
            .I(N__84540));
    Odrv4 I__20301 (
            .O(N__84540),
            .I(\pid_side.O_1_22 ));
    InMux I__20300 (
            .O(N__84537),
            .I(N__84530));
    InMux I__20299 (
            .O(N__84536),
            .I(N__84530));
    InMux I__20298 (
            .O(N__84535),
            .I(N__84527));
    LocalMux I__20297 (
            .O(N__84530),
            .I(N__84524));
    LocalMux I__20296 (
            .O(N__84527),
            .I(N__84519));
    Span4Mux_v I__20295 (
            .O(N__84524),
            .I(N__84519));
    Odrv4 I__20294 (
            .O(N__84519),
            .I(\pid_side.error_d_regZ0Z_20 ));
    InMux I__20293 (
            .O(N__84516),
            .I(N__84513));
    LocalMux I__20292 (
            .O(N__84513),
            .I(N__84510));
    Span4Mux_v I__20291 (
            .O(N__84510),
            .I(N__84507));
    Odrv4 I__20290 (
            .O(N__84507),
            .I(\pid_side.O_2_3 ));
    CascadeMux I__20289 (
            .O(N__84504),
            .I(N__84501));
    InMux I__20288 (
            .O(N__84501),
            .I(N__84497));
    InMux I__20287 (
            .O(N__84500),
            .I(N__84494));
    LocalMux I__20286 (
            .O(N__84497),
            .I(N__84489));
    LocalMux I__20285 (
            .O(N__84494),
            .I(N__84489));
    Span4Mux_h I__20284 (
            .O(N__84489),
            .I(N__84486));
    Span4Mux_h I__20283 (
            .O(N__84486),
            .I(N__84483));
    Span4Mux_s0_h I__20282 (
            .O(N__84483),
            .I(N__84480));
    Odrv4 I__20281 (
            .O(N__84480),
            .I(\pid_side.error_p_regZ0Z_0 ));
    InMux I__20280 (
            .O(N__84477),
            .I(N__84474));
    LocalMux I__20279 (
            .O(N__84474),
            .I(\pid_side.O_1_15 ));
    InMux I__20278 (
            .O(N__84471),
            .I(N__84468));
    LocalMux I__20277 (
            .O(N__84468),
            .I(N__84465));
    Odrv4 I__20276 (
            .O(N__84465),
            .I(\pid_side.O_2_17 ));
    InMux I__20275 (
            .O(N__84462),
            .I(N__84459));
    LocalMux I__20274 (
            .O(N__84459),
            .I(N__84453));
    InMux I__20273 (
            .O(N__84458),
            .I(N__84450));
    InMux I__20272 (
            .O(N__84457),
            .I(N__84445));
    InMux I__20271 (
            .O(N__84456),
            .I(N__84445));
    Span4Mux_h I__20270 (
            .O(N__84453),
            .I(N__84442));
    LocalMux I__20269 (
            .O(N__84450),
            .I(N__84439));
    LocalMux I__20268 (
            .O(N__84445),
            .I(N__84436));
    Span4Mux_v I__20267 (
            .O(N__84442),
            .I(N__84431));
    Span4Mux_v I__20266 (
            .O(N__84439),
            .I(N__84431));
    Span12Mux_h I__20265 (
            .O(N__84436),
            .I(N__84428));
    Odrv4 I__20264 (
            .O(N__84431),
            .I(\pid_side.error_p_regZ0Z_14 ));
    Odrv12 I__20263 (
            .O(N__84428),
            .I(\pid_side.error_p_regZ0Z_14 ));
    InMux I__20262 (
            .O(N__84423),
            .I(N__84420));
    LocalMux I__20261 (
            .O(N__84420),
            .I(\pid_side.O_2_10 ));
    CascadeMux I__20260 (
            .O(N__84417),
            .I(N__84413));
    CascadeMux I__20259 (
            .O(N__84416),
            .I(N__84410));
    InMux I__20258 (
            .O(N__84413),
            .I(N__84405));
    InMux I__20257 (
            .O(N__84410),
            .I(N__84405));
    LocalMux I__20256 (
            .O(N__84405),
            .I(N__84402));
    Span4Mux_v I__20255 (
            .O(N__84402),
            .I(N__84399));
    Span4Mux_h I__20254 (
            .O(N__84399),
            .I(N__84396));
    Span4Mux_h I__20253 (
            .O(N__84396),
            .I(N__84393));
    Odrv4 I__20252 (
            .O(N__84393),
            .I(\pid_side.error_p_regZ0Z_7 ));
    InMux I__20251 (
            .O(N__84390),
            .I(N__84387));
    LocalMux I__20250 (
            .O(N__84387),
            .I(\pid_side.O_2_11 ));
    InMux I__20249 (
            .O(N__84384),
            .I(N__84378));
    InMux I__20248 (
            .O(N__84383),
            .I(N__84378));
    LocalMux I__20247 (
            .O(N__84378),
            .I(N__84375));
    Span4Mux_h I__20246 (
            .O(N__84375),
            .I(N__84372));
    Span4Mux_h I__20245 (
            .O(N__84372),
            .I(N__84369));
    Span4Mux_h I__20244 (
            .O(N__84369),
            .I(N__84366));
    Odrv4 I__20243 (
            .O(N__84366),
            .I(\pid_side.error_p_regZ0Z_8 ));
    InMux I__20242 (
            .O(N__84363),
            .I(N__84360));
    LocalMux I__20241 (
            .O(N__84360),
            .I(\pid_side.O_2_16 ));
    InMux I__20240 (
            .O(N__84357),
            .I(N__84354));
    LocalMux I__20239 (
            .O(N__84354),
            .I(\pid_side.O_2_20 ));
    InMux I__20238 (
            .O(N__84351),
            .I(N__84345));
    InMux I__20237 (
            .O(N__84350),
            .I(N__84345));
    LocalMux I__20236 (
            .O(N__84345),
            .I(N__84342));
    Span4Mux_v I__20235 (
            .O(N__84342),
            .I(N__84339));
    Odrv4 I__20234 (
            .O(N__84339),
            .I(\pid_side.error_p_regZ0Z_17 ));
    InMux I__20233 (
            .O(N__84336),
            .I(N__84333));
    LocalMux I__20232 (
            .O(N__84333),
            .I(\pid_side.O_2_18 ));
    InMux I__20231 (
            .O(N__84330),
            .I(N__84324));
    InMux I__20230 (
            .O(N__84329),
            .I(N__84324));
    LocalMux I__20229 (
            .O(N__84324),
            .I(N__84321));
    Span12Mux_h I__20228 (
            .O(N__84321),
            .I(N__84318));
    Odrv12 I__20227 (
            .O(N__84318),
            .I(\pid_side.error_p_regZ0Z_15 ));
    InMux I__20226 (
            .O(N__84315),
            .I(N__84312));
    LocalMux I__20225 (
            .O(N__84312),
            .I(\pid_side.O_2_19 ));
    InMux I__20224 (
            .O(N__84309),
            .I(N__84305));
    InMux I__20223 (
            .O(N__84308),
            .I(N__84302));
    LocalMux I__20222 (
            .O(N__84305),
            .I(N__84297));
    LocalMux I__20221 (
            .O(N__84302),
            .I(N__84297));
    Span4Mux_v I__20220 (
            .O(N__84297),
            .I(N__84294));
    Odrv4 I__20219 (
            .O(N__84294),
            .I(\pid_side.error_p_regZ0Z_16 ));
    InMux I__20218 (
            .O(N__84291),
            .I(N__84288));
    LocalMux I__20217 (
            .O(N__84288),
            .I(\pid_side.O_2_23 ));
    InMux I__20216 (
            .O(N__84285),
            .I(N__84281));
    InMux I__20215 (
            .O(N__84284),
            .I(N__84278));
    LocalMux I__20214 (
            .O(N__84281),
            .I(N__84275));
    LocalMux I__20213 (
            .O(N__84278),
            .I(N__84272));
    Span4Mux_v I__20212 (
            .O(N__84275),
            .I(N__84267));
    Span4Mux_h I__20211 (
            .O(N__84272),
            .I(N__84267));
    Odrv4 I__20210 (
            .O(N__84267),
            .I(\pid_side.error_p_regZ0Z_20 ));
    InMux I__20209 (
            .O(N__84264),
            .I(N__84261));
    LocalMux I__20208 (
            .O(N__84261),
            .I(N__84257));
    InMux I__20207 (
            .O(N__84260),
            .I(N__84254));
    Span4Mux_v I__20206 (
            .O(N__84257),
            .I(N__84247));
    LocalMux I__20205 (
            .O(N__84254),
            .I(N__84247));
    InMux I__20204 (
            .O(N__84253),
            .I(N__84242));
    InMux I__20203 (
            .O(N__84252),
            .I(N__84242));
    Span4Mux_h I__20202 (
            .O(N__84247),
            .I(N__84239));
    LocalMux I__20201 (
            .O(N__84242),
            .I(\pid_side.error_d_reg_prevZ0Z_14 ));
    Odrv4 I__20200 (
            .O(N__84239),
            .I(\pid_side.error_d_reg_prevZ0Z_14 ));
    CascadeMux I__20199 (
            .O(N__84234),
            .I(\pid_side.N_2405_0_cascade_ ));
    InMux I__20198 (
            .O(N__84231),
            .I(N__84228));
    LocalMux I__20197 (
            .O(N__84228),
            .I(N__84225));
    Odrv12 I__20196 (
            .O(N__84225),
            .I(\pid_side.g0_2 ));
    InMux I__20195 (
            .O(N__84222),
            .I(N__84216));
    InMux I__20194 (
            .O(N__84221),
            .I(N__84216));
    LocalMux I__20193 (
            .O(N__84216),
            .I(N__84211));
    InMux I__20192 (
            .O(N__84215),
            .I(N__84205));
    InMux I__20191 (
            .O(N__84214),
            .I(N__84201));
    Span4Mux_v I__20190 (
            .O(N__84211),
            .I(N__84198));
    InMux I__20189 (
            .O(N__84210),
            .I(N__84195));
    InMux I__20188 (
            .O(N__84209),
            .I(N__84192));
    InMux I__20187 (
            .O(N__84208),
            .I(N__84189));
    LocalMux I__20186 (
            .O(N__84205),
            .I(N__84186));
    InMux I__20185 (
            .O(N__84204),
            .I(N__84183));
    LocalMux I__20184 (
            .O(N__84201),
            .I(N__84179));
    Span4Mux_h I__20183 (
            .O(N__84198),
            .I(N__84174));
    LocalMux I__20182 (
            .O(N__84195),
            .I(N__84174));
    LocalMux I__20181 (
            .O(N__84192),
            .I(N__84171));
    LocalMux I__20180 (
            .O(N__84189),
            .I(N__84168));
    Span4Mux_v I__20179 (
            .O(N__84186),
            .I(N__84165));
    LocalMux I__20178 (
            .O(N__84183),
            .I(N__84162));
    InMux I__20177 (
            .O(N__84182),
            .I(N__84157));
    Span4Mux_h I__20176 (
            .O(N__84179),
            .I(N__84151));
    Span4Mux_v I__20175 (
            .O(N__84174),
            .I(N__84151));
    Span4Mux_v I__20174 (
            .O(N__84171),
            .I(N__84148));
    Span4Mux_v I__20173 (
            .O(N__84168),
            .I(N__84144));
    Span4Mux_v I__20172 (
            .O(N__84165),
            .I(N__84139));
    Span4Mux_v I__20171 (
            .O(N__84162),
            .I(N__84139));
    InMux I__20170 (
            .O(N__84161),
            .I(N__84136));
    InMux I__20169 (
            .O(N__84160),
            .I(N__84133));
    LocalMux I__20168 (
            .O(N__84157),
            .I(N__84128));
    InMux I__20167 (
            .O(N__84156),
            .I(N__84125));
    Span4Mux_v I__20166 (
            .O(N__84151),
            .I(N__84120));
    Span4Mux_v I__20165 (
            .O(N__84148),
            .I(N__84117));
    InMux I__20164 (
            .O(N__84147),
            .I(N__84114));
    Sp12to4 I__20163 (
            .O(N__84144),
            .I(N__84109));
    Sp12to4 I__20162 (
            .O(N__84139),
            .I(N__84109));
    LocalMux I__20161 (
            .O(N__84136),
            .I(N__84106));
    LocalMux I__20160 (
            .O(N__84133),
            .I(N__84103));
    InMux I__20159 (
            .O(N__84132),
            .I(N__84098));
    InMux I__20158 (
            .O(N__84131),
            .I(N__84098));
    Span4Mux_v I__20157 (
            .O(N__84128),
            .I(N__84093));
    LocalMux I__20156 (
            .O(N__84125),
            .I(N__84093));
    InMux I__20155 (
            .O(N__84124),
            .I(N__84090));
    InMux I__20154 (
            .O(N__84123),
            .I(N__84087));
    Sp12to4 I__20153 (
            .O(N__84120),
            .I(N__84078));
    Sp12to4 I__20152 (
            .O(N__84117),
            .I(N__84078));
    LocalMux I__20151 (
            .O(N__84114),
            .I(N__84078));
    Span12Mux_h I__20150 (
            .O(N__84109),
            .I(N__84078));
    Span4Mux_h I__20149 (
            .O(N__84106),
            .I(N__84073));
    Span4Mux_v I__20148 (
            .O(N__84103),
            .I(N__84073));
    LocalMux I__20147 (
            .O(N__84098),
            .I(N__84070));
    Span4Mux_v I__20146 (
            .O(N__84093),
            .I(N__84065));
    LocalMux I__20145 (
            .O(N__84090),
            .I(N__84065));
    LocalMux I__20144 (
            .O(N__84087),
            .I(uart_pc_data_1));
    Odrv12 I__20143 (
            .O(N__84078),
            .I(uart_pc_data_1));
    Odrv4 I__20142 (
            .O(N__84073),
            .I(uart_pc_data_1));
    Odrv4 I__20141 (
            .O(N__84070),
            .I(uart_pc_data_1));
    Odrv4 I__20140 (
            .O(N__84065),
            .I(uart_pc_data_1));
    InMux I__20139 (
            .O(N__84054),
            .I(N__84050));
    InMux I__20138 (
            .O(N__84053),
            .I(N__84047));
    LocalMux I__20137 (
            .O(N__84050),
            .I(N__84044));
    LocalMux I__20136 (
            .O(N__84047),
            .I(N__84041));
    Span12Mux_s2_h I__20135 (
            .O(N__84044),
            .I(N__84038));
    Span4Mux_s1_h I__20134 (
            .O(N__84041),
            .I(N__84035));
    Odrv12 I__20133 (
            .O(N__84038),
            .I(xy_kd_1));
    Odrv4 I__20132 (
            .O(N__84035),
            .I(xy_kd_1));
    InMux I__20131 (
            .O(N__84030),
            .I(N__84025));
    InMux I__20130 (
            .O(N__84029),
            .I(N__84022));
    InMux I__20129 (
            .O(N__84028),
            .I(N__84016));
    LocalMux I__20128 (
            .O(N__84025),
            .I(N__84013));
    LocalMux I__20127 (
            .O(N__84022),
            .I(N__84010));
    InMux I__20126 (
            .O(N__84021),
            .I(N__84003));
    InMux I__20125 (
            .O(N__84020),
            .I(N__84003));
    InMux I__20124 (
            .O(N__84019),
            .I(N__84003));
    LocalMux I__20123 (
            .O(N__84016),
            .I(N__83997));
    Span4Mux_h I__20122 (
            .O(N__84013),
            .I(N__83994));
    Span4Mux_h I__20121 (
            .O(N__84010),
            .I(N__83989));
    LocalMux I__20120 (
            .O(N__84003),
            .I(N__83989));
    InMux I__20119 (
            .O(N__84002),
            .I(N__83985));
    InMux I__20118 (
            .O(N__84001),
            .I(N__83981));
    InMux I__20117 (
            .O(N__84000),
            .I(N__83977));
    Span4Mux_v I__20116 (
            .O(N__83997),
            .I(N__83974));
    Span4Mux_h I__20115 (
            .O(N__83994),
            .I(N__83969));
    Span4Mux_v I__20114 (
            .O(N__83989),
            .I(N__83969));
    InMux I__20113 (
            .O(N__83988),
            .I(N__83965));
    LocalMux I__20112 (
            .O(N__83985),
            .I(N__83962));
    InMux I__20111 (
            .O(N__83984),
            .I(N__83959));
    LocalMux I__20110 (
            .O(N__83981),
            .I(N__83956));
    InMux I__20109 (
            .O(N__83980),
            .I(N__83953));
    LocalMux I__20108 (
            .O(N__83977),
            .I(N__83948));
    Sp12to4 I__20107 (
            .O(N__83974),
            .I(N__83948));
    Span4Mux_v I__20106 (
            .O(N__83969),
            .I(N__83942));
    InMux I__20105 (
            .O(N__83968),
            .I(N__83939));
    LocalMux I__20104 (
            .O(N__83965),
            .I(N__83935));
    Span4Mux_h I__20103 (
            .O(N__83962),
            .I(N__83932));
    LocalMux I__20102 (
            .O(N__83959),
            .I(N__83929));
    Span4Mux_h I__20101 (
            .O(N__83956),
            .I(N__83926));
    LocalMux I__20100 (
            .O(N__83953),
            .I(N__83923));
    Span12Mux_s9_h I__20099 (
            .O(N__83948),
            .I(N__83920));
    InMux I__20098 (
            .O(N__83947),
            .I(N__83915));
    InMux I__20097 (
            .O(N__83946),
            .I(N__83915));
    InMux I__20096 (
            .O(N__83945),
            .I(N__83912));
    Sp12to4 I__20095 (
            .O(N__83942),
            .I(N__83907));
    LocalMux I__20094 (
            .O(N__83939),
            .I(N__83907));
    InMux I__20093 (
            .O(N__83938),
            .I(N__83904));
    Span4Mux_h I__20092 (
            .O(N__83935),
            .I(N__83893));
    Span4Mux_h I__20091 (
            .O(N__83932),
            .I(N__83893));
    Span4Mux_v I__20090 (
            .O(N__83929),
            .I(N__83893));
    Span4Mux_v I__20089 (
            .O(N__83926),
            .I(N__83893));
    Span4Mux_h I__20088 (
            .O(N__83923),
            .I(N__83893));
    Span12Mux_h I__20087 (
            .O(N__83920),
            .I(N__83888));
    LocalMux I__20086 (
            .O(N__83915),
            .I(N__83888));
    LocalMux I__20085 (
            .O(N__83912),
            .I(N__83885));
    Odrv12 I__20084 (
            .O(N__83907),
            .I(uart_pc_data_3));
    LocalMux I__20083 (
            .O(N__83904),
            .I(uart_pc_data_3));
    Odrv4 I__20082 (
            .O(N__83893),
            .I(uart_pc_data_3));
    Odrv12 I__20081 (
            .O(N__83888),
            .I(uart_pc_data_3));
    Odrv4 I__20080 (
            .O(N__83885),
            .I(uart_pc_data_3));
    InMux I__20079 (
            .O(N__83874),
            .I(N__83871));
    LocalMux I__20078 (
            .O(N__83871),
            .I(N__83867));
    InMux I__20077 (
            .O(N__83870),
            .I(N__83864));
    Span4Mux_v I__20076 (
            .O(N__83867),
            .I(N__83861));
    LocalMux I__20075 (
            .O(N__83864),
            .I(N__83858));
    Span4Mux_v I__20074 (
            .O(N__83861),
            .I(N__83853));
    Span4Mux_v I__20073 (
            .O(N__83858),
            .I(N__83853));
    Odrv4 I__20072 (
            .O(N__83853),
            .I(xy_kd_3));
    InMux I__20071 (
            .O(N__83850),
            .I(N__83841));
    InMux I__20070 (
            .O(N__83849),
            .I(N__83841));
    InMux I__20069 (
            .O(N__83848),
            .I(N__83841));
    LocalMux I__20068 (
            .O(N__83841),
            .I(N__83838));
    Span4Mux_v I__20067 (
            .O(N__83838),
            .I(N__83832));
    InMux I__20066 (
            .O(N__83837),
            .I(N__83829));
    InMux I__20065 (
            .O(N__83836),
            .I(N__83825));
    InMux I__20064 (
            .O(N__83835),
            .I(N__83822));
    Span4Mux_v I__20063 (
            .O(N__83832),
            .I(N__83817));
    LocalMux I__20062 (
            .O(N__83829),
            .I(N__83817));
    InMux I__20061 (
            .O(N__83828),
            .I(N__83814));
    LocalMux I__20060 (
            .O(N__83825),
            .I(N__83811));
    LocalMux I__20059 (
            .O(N__83822),
            .I(N__83808));
    Span4Mux_v I__20058 (
            .O(N__83817),
            .I(N__83804));
    LocalMux I__20057 (
            .O(N__83814),
            .I(N__83801));
    Span4Mux_v I__20056 (
            .O(N__83811),
            .I(N__83798));
    Span4Mux_v I__20055 (
            .O(N__83808),
            .I(N__83791));
    InMux I__20054 (
            .O(N__83807),
            .I(N__83788));
    Span4Mux_h I__20053 (
            .O(N__83804),
            .I(N__83782));
    Span4Mux_v I__20052 (
            .O(N__83801),
            .I(N__83782));
    Sp12to4 I__20051 (
            .O(N__83798),
            .I(N__83779));
    InMux I__20050 (
            .O(N__83797),
            .I(N__83776));
    InMux I__20049 (
            .O(N__83796),
            .I(N__83773));
    InMux I__20048 (
            .O(N__83795),
            .I(N__83770));
    InMux I__20047 (
            .O(N__83794),
            .I(N__83766));
    Span4Mux_v I__20046 (
            .O(N__83791),
            .I(N__83761));
    LocalMux I__20045 (
            .O(N__83788),
            .I(N__83761));
    InMux I__20044 (
            .O(N__83787),
            .I(N__83758));
    Sp12to4 I__20043 (
            .O(N__83782),
            .I(N__83750));
    Span12Mux_s9_h I__20042 (
            .O(N__83779),
            .I(N__83750));
    LocalMux I__20041 (
            .O(N__83776),
            .I(N__83747));
    LocalMux I__20040 (
            .O(N__83773),
            .I(N__83744));
    LocalMux I__20039 (
            .O(N__83770),
            .I(N__83741));
    InMux I__20038 (
            .O(N__83769),
            .I(N__83738));
    LocalMux I__20037 (
            .O(N__83766),
            .I(N__83735));
    Span4Mux_h I__20036 (
            .O(N__83761),
            .I(N__83732));
    LocalMux I__20035 (
            .O(N__83758),
            .I(N__83729));
    InMux I__20034 (
            .O(N__83757),
            .I(N__83724));
    InMux I__20033 (
            .O(N__83756),
            .I(N__83724));
    InMux I__20032 (
            .O(N__83755),
            .I(N__83720));
    Span12Mux_h I__20031 (
            .O(N__83750),
            .I(N__83717));
    Span4Mux_v I__20030 (
            .O(N__83747),
            .I(N__83714));
    Span4Mux_h I__20029 (
            .O(N__83744),
            .I(N__83707));
    Span4Mux_v I__20028 (
            .O(N__83741),
            .I(N__83707));
    LocalMux I__20027 (
            .O(N__83738),
            .I(N__83707));
    Span4Mux_h I__20026 (
            .O(N__83735),
            .I(N__83698));
    Span4Mux_h I__20025 (
            .O(N__83732),
            .I(N__83698));
    Span4Mux_v I__20024 (
            .O(N__83729),
            .I(N__83698));
    LocalMux I__20023 (
            .O(N__83724),
            .I(N__83698));
    InMux I__20022 (
            .O(N__83723),
            .I(N__83695));
    LocalMux I__20021 (
            .O(N__83720),
            .I(uart_pc_data_0));
    Odrv12 I__20020 (
            .O(N__83717),
            .I(uart_pc_data_0));
    Odrv4 I__20019 (
            .O(N__83714),
            .I(uart_pc_data_0));
    Odrv4 I__20018 (
            .O(N__83707),
            .I(uart_pc_data_0));
    Odrv4 I__20017 (
            .O(N__83698),
            .I(uart_pc_data_0));
    LocalMux I__20016 (
            .O(N__83695),
            .I(uart_pc_data_0));
    InMux I__20015 (
            .O(N__83682),
            .I(N__83678));
    InMux I__20014 (
            .O(N__83681),
            .I(N__83675));
    LocalMux I__20013 (
            .O(N__83678),
            .I(N__83672));
    LocalMux I__20012 (
            .O(N__83675),
            .I(N__83669));
    Span4Mux_v I__20011 (
            .O(N__83672),
            .I(N__83666));
    Span4Mux_v I__20010 (
            .O(N__83669),
            .I(N__83663));
    Span4Mux_v I__20009 (
            .O(N__83666),
            .I(N__83658));
    Span4Mux_s0_h I__20008 (
            .O(N__83663),
            .I(N__83658));
    Odrv4 I__20007 (
            .O(N__83658),
            .I(xy_kd_0));
    InMux I__20006 (
            .O(N__83655),
            .I(N__83652));
    LocalMux I__20005 (
            .O(N__83652),
            .I(N__83649));
    Span4Mux_h I__20004 (
            .O(N__83649),
            .I(N__83646));
    Odrv4 I__20003 (
            .O(N__83646),
            .I(\pid_front.O_22 ));
    InMux I__20002 (
            .O(N__83643),
            .I(N__83636));
    InMux I__20001 (
            .O(N__83642),
            .I(N__83636));
    InMux I__20000 (
            .O(N__83641),
            .I(N__83633));
    LocalMux I__19999 (
            .O(N__83636),
            .I(N__83630));
    LocalMux I__19998 (
            .O(N__83633),
            .I(N__83627));
    Span4Mux_h I__19997 (
            .O(N__83630),
            .I(N__83624));
    Span12Mux_v I__19996 (
            .O(N__83627),
            .I(N__83621));
    Span4Mux_h I__19995 (
            .O(N__83624),
            .I(N__83618));
    Span12Mux_h I__19994 (
            .O(N__83621),
            .I(N__83615));
    Span4Mux_h I__19993 (
            .O(N__83618),
            .I(N__83612));
    Odrv12 I__19992 (
            .O(N__83615),
            .I(\pid_front.error_d_regZ0Z_20 ));
    Odrv4 I__19991 (
            .O(N__83612),
            .I(\pid_front.error_d_regZ0Z_20 ));
    InMux I__19990 (
            .O(N__83607),
            .I(N__83604));
    LocalMux I__19989 (
            .O(N__83604),
            .I(N__83601));
    Odrv4 I__19988 (
            .O(N__83601),
            .I(\pid_side.O_2_22 ));
    InMux I__19987 (
            .O(N__83598),
            .I(N__83592));
    InMux I__19986 (
            .O(N__83597),
            .I(N__83592));
    LocalMux I__19985 (
            .O(N__83592),
            .I(N__83589));
    Span4Mux_v I__19984 (
            .O(N__83589),
            .I(N__83586));
    Odrv4 I__19983 (
            .O(N__83586),
            .I(\pid_side.error_p_regZ0Z_19 ));
    InMux I__19982 (
            .O(N__83583),
            .I(N__83580));
    LocalMux I__19981 (
            .O(N__83580),
            .I(N__83577));
    Odrv4 I__19980 (
            .O(N__83577),
            .I(\pid_side.O_2_24 ));
    CascadeMux I__19979 (
            .O(N__83574),
            .I(N__83570));
    CascadeMux I__19978 (
            .O(N__83573),
            .I(N__83563));
    InMux I__19977 (
            .O(N__83570),
            .I(N__83553));
    InMux I__19976 (
            .O(N__83569),
            .I(N__83553));
    InMux I__19975 (
            .O(N__83568),
            .I(N__83553));
    InMux I__19974 (
            .O(N__83567),
            .I(N__83553));
    InMux I__19973 (
            .O(N__83566),
            .I(N__83541));
    InMux I__19972 (
            .O(N__83563),
            .I(N__83541));
    InMux I__19971 (
            .O(N__83562),
            .I(N__83541));
    LocalMux I__19970 (
            .O(N__83553),
            .I(N__83538));
    CascadeMux I__19969 (
            .O(N__83552),
            .I(N__83534));
    InMux I__19968 (
            .O(N__83551),
            .I(N__83523));
    InMux I__19967 (
            .O(N__83550),
            .I(N__83523));
    InMux I__19966 (
            .O(N__83549),
            .I(N__83523));
    InMux I__19965 (
            .O(N__83548),
            .I(N__83523));
    LocalMux I__19964 (
            .O(N__83541),
            .I(N__83520));
    Span4Mux_h I__19963 (
            .O(N__83538),
            .I(N__83517));
    InMux I__19962 (
            .O(N__83537),
            .I(N__83508));
    InMux I__19961 (
            .O(N__83534),
            .I(N__83508));
    InMux I__19960 (
            .O(N__83533),
            .I(N__83508));
    InMux I__19959 (
            .O(N__83532),
            .I(N__83508));
    LocalMux I__19958 (
            .O(N__83523),
            .I(N__83505));
    Span4Mux_v I__19957 (
            .O(N__83520),
            .I(N__83502));
    Span4Mux_v I__19956 (
            .O(N__83517),
            .I(N__83499));
    LocalMux I__19955 (
            .O(N__83508),
            .I(N__83496));
    Span4Mux_h I__19954 (
            .O(N__83505),
            .I(N__83493));
    Span4Mux_h I__19953 (
            .O(N__83502),
            .I(N__83490));
    Sp12to4 I__19952 (
            .O(N__83499),
            .I(N__83485));
    Sp12to4 I__19951 (
            .O(N__83496),
            .I(N__83485));
    Span4Mux_h I__19950 (
            .O(N__83493),
            .I(N__83480));
    Span4Mux_h I__19949 (
            .O(N__83490),
            .I(N__83480));
    Odrv12 I__19948 (
            .O(N__83485),
            .I(\pid_side.error_p_regZ0Z_21 ));
    Odrv4 I__19947 (
            .O(N__83480),
            .I(\pid_side.error_p_regZ0Z_21 ));
    InMux I__19946 (
            .O(N__83475),
            .I(N__83472));
    LocalMux I__19945 (
            .O(N__83472),
            .I(N__83469));
    Odrv4 I__19944 (
            .O(N__83469),
            .I(\pid_side.O_2_21 ));
    InMux I__19943 (
            .O(N__83466),
            .I(N__83460));
    InMux I__19942 (
            .O(N__83465),
            .I(N__83460));
    LocalMux I__19941 (
            .O(N__83460),
            .I(N__83457));
    Span4Mux_h I__19940 (
            .O(N__83457),
            .I(N__83454));
    Odrv4 I__19939 (
            .O(N__83454),
            .I(\pid_side.error_p_regZ0Z_18 ));
    InMux I__19938 (
            .O(N__83451),
            .I(N__83445));
    InMux I__19937 (
            .O(N__83450),
            .I(N__83445));
    LocalMux I__19936 (
            .O(N__83445),
            .I(\pid_side.error_d_reg_prevZ0Z_17 ));
    InMux I__19935 (
            .O(N__83442),
            .I(N__83436));
    InMux I__19934 (
            .O(N__83441),
            .I(N__83436));
    LocalMux I__19933 (
            .O(N__83436),
            .I(N__83433));
    Span4Mux_h I__19932 (
            .O(N__83433),
            .I(N__83430));
    Span4Mux_h I__19931 (
            .O(N__83430),
            .I(N__83427));
    Odrv4 I__19930 (
            .O(N__83427),
            .I(\pid_side.error_d_reg_prev_esr_RNIE4JOZ0Z_17 ));
    InMux I__19929 (
            .O(N__83424),
            .I(N__83418));
    InMux I__19928 (
            .O(N__83423),
            .I(N__83418));
    LocalMux I__19927 (
            .O(N__83418),
            .I(N__83415));
    Span4Mux_v I__19926 (
            .O(N__83415),
            .I(N__83412));
    Span4Mux_h I__19925 (
            .O(N__83412),
            .I(N__83409));
    Odrv4 I__19924 (
            .O(N__83409),
            .I(\pid_side.error_d_reg_prev_esr_RNIH7JO_0Z0Z_18 ));
    CEMux I__19923 (
            .O(N__83406),
            .I(N__83394));
    CEMux I__19922 (
            .O(N__83405),
            .I(N__83389));
    CEMux I__19921 (
            .O(N__83404),
            .I(N__83386));
    CEMux I__19920 (
            .O(N__83403),
            .I(N__83382));
    CEMux I__19919 (
            .O(N__83402),
            .I(N__83379));
    CEMux I__19918 (
            .O(N__83401),
            .I(N__83376));
    CEMux I__19917 (
            .O(N__83400),
            .I(N__83373));
    CEMux I__19916 (
            .O(N__83399),
            .I(N__83370));
    CEMux I__19915 (
            .O(N__83398),
            .I(N__83367));
    CEMux I__19914 (
            .O(N__83397),
            .I(N__83364));
    LocalMux I__19913 (
            .O(N__83394),
            .I(N__83361));
    CEMux I__19912 (
            .O(N__83393),
            .I(N__83358));
    CEMux I__19911 (
            .O(N__83392),
            .I(N__83355));
    LocalMux I__19910 (
            .O(N__83389),
            .I(N__83350));
    LocalMux I__19909 (
            .O(N__83386),
            .I(N__83350));
    CEMux I__19908 (
            .O(N__83385),
            .I(N__83347));
    LocalMux I__19907 (
            .O(N__83382),
            .I(N__83342));
    LocalMux I__19906 (
            .O(N__83379),
            .I(N__83342));
    LocalMux I__19905 (
            .O(N__83376),
            .I(N__83339));
    LocalMux I__19904 (
            .O(N__83373),
            .I(N__83336));
    LocalMux I__19903 (
            .O(N__83370),
            .I(N__83333));
    LocalMux I__19902 (
            .O(N__83367),
            .I(N__83330));
    LocalMux I__19901 (
            .O(N__83364),
            .I(N__83326));
    Span4Mux_s3_h I__19900 (
            .O(N__83361),
            .I(N__83321));
    LocalMux I__19899 (
            .O(N__83358),
            .I(N__83321));
    LocalMux I__19898 (
            .O(N__83355),
            .I(N__83316));
    Span4Mux_v I__19897 (
            .O(N__83350),
            .I(N__83316));
    LocalMux I__19896 (
            .O(N__83347),
            .I(N__83313));
    Span4Mux_v I__19895 (
            .O(N__83342),
            .I(N__83308));
    Span4Mux_v I__19894 (
            .O(N__83339),
            .I(N__83308));
    Span4Mux_v I__19893 (
            .O(N__83336),
            .I(N__83303));
    Span4Mux_v I__19892 (
            .O(N__83333),
            .I(N__83303));
    Span4Mux_h I__19891 (
            .O(N__83330),
            .I(N__83300));
    CEMux I__19890 (
            .O(N__83329),
            .I(N__83297));
    Span4Mux_v I__19889 (
            .O(N__83326),
            .I(N__83290));
    Span4Mux_h I__19888 (
            .O(N__83321),
            .I(N__83290));
    Span4Mux_h I__19887 (
            .O(N__83316),
            .I(N__83290));
    Span4Mux_v I__19886 (
            .O(N__83313),
            .I(N__83285));
    Span4Mux_h I__19885 (
            .O(N__83308),
            .I(N__83285));
    Span4Mux_h I__19884 (
            .O(N__83303),
            .I(N__83282));
    Span4Mux_h I__19883 (
            .O(N__83300),
            .I(N__83279));
    LocalMux I__19882 (
            .O(N__83297),
            .I(N__83274));
    Span4Mux_h I__19881 (
            .O(N__83290),
            .I(N__83274));
    Span4Mux_h I__19880 (
            .O(N__83285),
            .I(N__83271));
    Odrv4 I__19879 (
            .O(N__83282),
            .I(\pid_side.N_838_0 ));
    Odrv4 I__19878 (
            .O(N__83279),
            .I(\pid_side.N_838_0 ));
    Odrv4 I__19877 (
            .O(N__83274),
            .I(\pid_side.N_838_0 ));
    Odrv4 I__19876 (
            .O(N__83271),
            .I(\pid_side.N_838_0 ));
    SRMux I__19875 (
            .O(N__83262),
            .I(N__83258));
    SRMux I__19874 (
            .O(N__83261),
            .I(N__83251));
    LocalMux I__19873 (
            .O(N__83258),
            .I(N__83248));
    SRMux I__19872 (
            .O(N__83257),
            .I(N__83245));
    SRMux I__19871 (
            .O(N__83256),
            .I(N__83241));
    SRMux I__19870 (
            .O(N__83255),
            .I(N__83237));
    SRMux I__19869 (
            .O(N__83254),
            .I(N__83233));
    LocalMux I__19868 (
            .O(N__83251),
            .I(N__83230));
    Span4Mux_h I__19867 (
            .O(N__83248),
            .I(N__83223));
    LocalMux I__19866 (
            .O(N__83245),
            .I(N__83223));
    SRMux I__19865 (
            .O(N__83244),
            .I(N__83220));
    LocalMux I__19864 (
            .O(N__83241),
            .I(N__83215));
    SRMux I__19863 (
            .O(N__83240),
            .I(N__83212));
    LocalMux I__19862 (
            .O(N__83237),
            .I(N__83209));
    SRMux I__19861 (
            .O(N__83236),
            .I(N__83206));
    LocalMux I__19860 (
            .O(N__83233),
            .I(N__83201));
    Span4Mux_v I__19859 (
            .O(N__83230),
            .I(N__83201));
    SRMux I__19858 (
            .O(N__83229),
            .I(N__83198));
    SRMux I__19857 (
            .O(N__83228),
            .I(N__83195));
    Span4Mux_v I__19856 (
            .O(N__83223),
            .I(N__83190));
    LocalMux I__19855 (
            .O(N__83220),
            .I(N__83190));
    SRMux I__19854 (
            .O(N__83219),
            .I(N__83187));
    SRMux I__19853 (
            .O(N__83218),
            .I(N__83184));
    Span4Mux_v I__19852 (
            .O(N__83215),
            .I(N__83178));
    LocalMux I__19851 (
            .O(N__83212),
            .I(N__83178));
    Span4Mux_v I__19850 (
            .O(N__83209),
            .I(N__83174));
    LocalMux I__19849 (
            .O(N__83206),
            .I(N__83171));
    Span4Mux_h I__19848 (
            .O(N__83201),
            .I(N__83166));
    LocalMux I__19847 (
            .O(N__83198),
            .I(N__83166));
    LocalMux I__19846 (
            .O(N__83195),
            .I(N__83159));
    Span4Mux_v I__19845 (
            .O(N__83190),
            .I(N__83159));
    LocalMux I__19844 (
            .O(N__83187),
            .I(N__83159));
    LocalMux I__19843 (
            .O(N__83184),
            .I(N__83156));
    SRMux I__19842 (
            .O(N__83183),
            .I(N__83153));
    Span4Mux_v I__19841 (
            .O(N__83178),
            .I(N__83150));
    InMux I__19840 (
            .O(N__83177),
            .I(N__83147));
    Span4Mux_h I__19839 (
            .O(N__83174),
            .I(N__83142));
    Span4Mux_h I__19838 (
            .O(N__83171),
            .I(N__83142));
    Span4Mux_h I__19837 (
            .O(N__83166),
            .I(N__83139));
    Span4Mux_h I__19836 (
            .O(N__83159),
            .I(N__83136));
    Span4Mux_v I__19835 (
            .O(N__83156),
            .I(N__83131));
    LocalMux I__19834 (
            .O(N__83153),
            .I(N__83131));
    Span4Mux_h I__19833 (
            .O(N__83150),
            .I(N__83128));
    LocalMux I__19832 (
            .O(N__83147),
            .I(N__83125));
    Span4Mux_h I__19831 (
            .O(N__83142),
            .I(N__83120));
    Span4Mux_v I__19830 (
            .O(N__83139),
            .I(N__83120));
    Span4Mux_h I__19829 (
            .O(N__83136),
            .I(N__83115));
    Span4Mux_v I__19828 (
            .O(N__83131),
            .I(N__83115));
    Span4Mux_h I__19827 (
            .O(N__83128),
            .I(N__83110));
    Span4Mux_v I__19826 (
            .O(N__83125),
            .I(N__83110));
    Odrv4 I__19825 (
            .O(N__83120),
            .I(\pid_side.state_RNIIIOOZ0Z_0 ));
    Odrv4 I__19824 (
            .O(N__83115),
            .I(\pid_side.state_RNIIIOOZ0Z_0 ));
    Odrv4 I__19823 (
            .O(N__83110),
            .I(\pid_side.state_RNIIIOOZ0Z_0 ));
    InMux I__19822 (
            .O(N__83103),
            .I(N__83097));
    InMux I__19821 (
            .O(N__83102),
            .I(N__83097));
    LocalMux I__19820 (
            .O(N__83097),
            .I(\pid_side.error_d_reg_prevZ0Z_18 ));
    InMux I__19819 (
            .O(N__83094),
            .I(N__83090));
    InMux I__19818 (
            .O(N__83093),
            .I(N__83087));
    LocalMux I__19817 (
            .O(N__83090),
            .I(N__83084));
    LocalMux I__19816 (
            .O(N__83087),
            .I(N__83081));
    Span4Mux_h I__19815 (
            .O(N__83084),
            .I(N__83078));
    Span4Mux_h I__19814 (
            .O(N__83081),
            .I(N__83075));
    Span4Mux_h I__19813 (
            .O(N__83078),
            .I(N__83072));
    Span4Mux_h I__19812 (
            .O(N__83075),
            .I(N__83069));
    Odrv4 I__19811 (
            .O(N__83072),
            .I(\pid_side.error_d_reg_prev_esr_RNIH7JOZ0Z_18 ));
    Odrv4 I__19810 (
            .O(N__83069),
            .I(\pid_side.error_d_reg_prev_esr_RNIH7JOZ0Z_18 ));
    InMux I__19809 (
            .O(N__83064),
            .I(N__83061));
    LocalMux I__19808 (
            .O(N__83061),
            .I(N__83058));
    Span4Mux_v I__19807 (
            .O(N__83058),
            .I(N__83055));
    Odrv4 I__19806 (
            .O(N__83055),
            .I(\pid_side.O_1_3 ));
    InMux I__19805 (
            .O(N__83052),
            .I(N__83049));
    LocalMux I__19804 (
            .O(N__83049),
            .I(N__83046));
    Span4Mux_v I__19803 (
            .O(N__83046),
            .I(N__83038));
    InMux I__19802 (
            .O(N__83045),
            .I(N__83029));
    InMux I__19801 (
            .O(N__83044),
            .I(N__83029));
    InMux I__19800 (
            .O(N__83043),
            .I(N__83029));
    InMux I__19799 (
            .O(N__83042),
            .I(N__83029));
    InMux I__19798 (
            .O(N__83041),
            .I(N__83026));
    Span4Mux_h I__19797 (
            .O(N__83038),
            .I(N__83021));
    LocalMux I__19796 (
            .O(N__83029),
            .I(N__83021));
    LocalMux I__19795 (
            .O(N__83026),
            .I(\pid_side.error_d_regZ0Z_1 ));
    Odrv4 I__19794 (
            .O(N__83021),
            .I(\pid_side.error_d_regZ0Z_1 ));
    InMux I__19793 (
            .O(N__83016),
            .I(N__83013));
    LocalMux I__19792 (
            .O(N__83013),
            .I(N__83008));
    InMux I__19791 (
            .O(N__83012),
            .I(N__83003));
    InMux I__19790 (
            .O(N__83011),
            .I(N__83003));
    Span4Mux_h I__19789 (
            .O(N__83008),
            .I(N__82999));
    LocalMux I__19788 (
            .O(N__83003),
            .I(N__82996));
    InMux I__19787 (
            .O(N__83002),
            .I(N__82993));
    Span4Mux_v I__19786 (
            .O(N__82999),
            .I(N__82986));
    Span4Mux_v I__19785 (
            .O(N__82996),
            .I(N__82986));
    LocalMux I__19784 (
            .O(N__82993),
            .I(N__82986));
    Odrv4 I__19783 (
            .O(N__82986),
            .I(\pid_side.error_d_reg_prev_esr_RNI2OIO_4Z0Z_13 ));
    InMux I__19782 (
            .O(N__82983),
            .I(N__82980));
    LocalMux I__19781 (
            .O(N__82980),
            .I(N__82977));
    Span4Mux_s3_h I__19780 (
            .O(N__82977),
            .I(N__82973));
    InMux I__19779 (
            .O(N__82976),
            .I(N__82970));
    Odrv4 I__19778 (
            .O(N__82973),
            .I(\pid_side.error_d_reg_prevZ0Z_20 ));
    LocalMux I__19777 (
            .O(N__82970),
            .I(\pid_side.error_d_reg_prevZ0Z_20 ));
    InMux I__19776 (
            .O(N__82965),
            .I(N__82962));
    LocalMux I__19775 (
            .O(N__82962),
            .I(N__82958));
    InMux I__19774 (
            .O(N__82961),
            .I(N__82955));
    Span4Mux_h I__19773 (
            .O(N__82958),
            .I(N__82952));
    LocalMux I__19772 (
            .O(N__82955),
            .I(N__82949));
    Span4Mux_h I__19771 (
            .O(N__82952),
            .I(N__82946));
    Span4Mux_h I__19770 (
            .O(N__82949),
            .I(N__82943));
    Odrv4 I__19769 (
            .O(N__82946),
            .I(\pid_side.error_d_reg_prev_esr_RNISKLOZ0Z_20 ));
    Odrv4 I__19768 (
            .O(N__82943),
            .I(\pid_side.error_d_reg_prev_esr_RNISKLOZ0Z_20 ));
    InMux I__19767 (
            .O(N__82938),
            .I(N__82934));
    InMux I__19766 (
            .O(N__82937),
            .I(N__82931));
    LocalMux I__19765 (
            .O(N__82934),
            .I(N__82928));
    LocalMux I__19764 (
            .O(N__82931),
            .I(\pid_side.error_d_reg_prevZ0Z_16 ));
    Odrv4 I__19763 (
            .O(N__82928),
            .I(\pid_side.error_d_reg_prevZ0Z_16 ));
    CascadeMux I__19762 (
            .O(N__82923),
            .I(N__82920));
    InMux I__19761 (
            .O(N__82920),
            .I(N__82914));
    InMux I__19760 (
            .O(N__82919),
            .I(N__82914));
    LocalMux I__19759 (
            .O(N__82914),
            .I(N__82911));
    Span4Mux_h I__19758 (
            .O(N__82911),
            .I(N__82908));
    Odrv4 I__19757 (
            .O(N__82908),
            .I(\pid_side.error_d_reg_prev_esr_RNIB1JO_0Z0Z_16 ));
    InMux I__19756 (
            .O(N__82905),
            .I(N__82902));
    LocalMux I__19755 (
            .O(N__82902),
            .I(N__82899));
    Span4Mux_h I__19754 (
            .O(N__82899),
            .I(N__82896));
    Odrv4 I__19753 (
            .O(N__82896),
            .I(\pid_side.O_1_13 ));
    InMux I__19752 (
            .O(N__82893),
            .I(N__82882));
    InMux I__19751 (
            .O(N__82892),
            .I(N__82882));
    InMux I__19750 (
            .O(N__82891),
            .I(N__82882));
    InMux I__19749 (
            .O(N__82890),
            .I(N__82877));
    InMux I__19748 (
            .O(N__82889),
            .I(N__82877));
    LocalMux I__19747 (
            .O(N__82882),
            .I(\pid_side.error_d_regZ0Z_11 ));
    LocalMux I__19746 (
            .O(N__82877),
            .I(\pid_side.error_d_regZ0Z_11 ));
    InMux I__19745 (
            .O(N__82872),
            .I(N__82869));
    LocalMux I__19744 (
            .O(N__82869),
            .I(N__82865));
    InMux I__19743 (
            .O(N__82868),
            .I(N__82862));
    Span4Mux_v I__19742 (
            .O(N__82865),
            .I(N__82857));
    LocalMux I__19741 (
            .O(N__82862),
            .I(N__82857));
    Span4Mux_h I__19740 (
            .O(N__82857),
            .I(N__82854));
    Odrv4 I__19739 (
            .O(N__82854),
            .I(\pid_side.O_1_14 ));
    InMux I__19738 (
            .O(N__82851),
            .I(N__82847));
    InMux I__19737 (
            .O(N__82850),
            .I(N__82844));
    LocalMux I__19736 (
            .O(N__82847),
            .I(N__82838));
    LocalMux I__19735 (
            .O(N__82844),
            .I(N__82835));
    CascadeMux I__19734 (
            .O(N__82843),
            .I(N__82828));
    InMux I__19733 (
            .O(N__82842),
            .I(N__82822));
    InMux I__19732 (
            .O(N__82841),
            .I(N__82822));
    Span4Mux_h I__19731 (
            .O(N__82838),
            .I(N__82819));
    Span4Mux_h I__19730 (
            .O(N__82835),
            .I(N__82816));
    InMux I__19729 (
            .O(N__82834),
            .I(N__82811));
    InMux I__19728 (
            .O(N__82833),
            .I(N__82811));
    InMux I__19727 (
            .O(N__82832),
            .I(N__82802));
    InMux I__19726 (
            .O(N__82831),
            .I(N__82802));
    InMux I__19725 (
            .O(N__82828),
            .I(N__82802));
    InMux I__19724 (
            .O(N__82827),
            .I(N__82802));
    LocalMux I__19723 (
            .O(N__82822),
            .I(N__82799));
    Odrv4 I__19722 (
            .O(N__82819),
            .I(\pid_side.error_d_regZ0Z_12 ));
    Odrv4 I__19721 (
            .O(N__82816),
            .I(\pid_side.error_d_regZ0Z_12 ));
    LocalMux I__19720 (
            .O(N__82811),
            .I(\pid_side.error_d_regZ0Z_12 ));
    LocalMux I__19719 (
            .O(N__82802),
            .I(\pid_side.error_d_regZ0Z_12 ));
    Odrv4 I__19718 (
            .O(N__82799),
            .I(\pid_side.error_d_regZ0Z_12 ));
    InMux I__19717 (
            .O(N__82788),
            .I(N__82785));
    LocalMux I__19716 (
            .O(N__82785),
            .I(N__82782));
    Span4Mux_v I__19715 (
            .O(N__82782),
            .I(N__82779));
    Odrv4 I__19714 (
            .O(N__82779),
            .I(\pid_front.O_16 ));
    InMux I__19713 (
            .O(N__82776),
            .I(N__82772));
    InMux I__19712 (
            .O(N__82775),
            .I(N__82766));
    LocalMux I__19711 (
            .O(N__82772),
            .I(N__82763));
    InMux I__19710 (
            .O(N__82771),
            .I(N__82760));
    InMux I__19709 (
            .O(N__82770),
            .I(N__82757));
    InMux I__19708 (
            .O(N__82769),
            .I(N__82754));
    LocalMux I__19707 (
            .O(N__82766),
            .I(N__82747));
    Span4Mux_v I__19706 (
            .O(N__82763),
            .I(N__82747));
    LocalMux I__19705 (
            .O(N__82760),
            .I(N__82747));
    LocalMux I__19704 (
            .O(N__82757),
            .I(N__82744));
    LocalMux I__19703 (
            .O(N__82754),
            .I(N__82741));
    Span4Mux_h I__19702 (
            .O(N__82747),
            .I(N__82738));
    Span4Mux_h I__19701 (
            .O(N__82744),
            .I(N__82733));
    Span4Mux_v I__19700 (
            .O(N__82741),
            .I(N__82733));
    Span4Mux_h I__19699 (
            .O(N__82738),
            .I(N__82730));
    Span4Mux_h I__19698 (
            .O(N__82733),
            .I(N__82727));
    Span4Mux_h I__19697 (
            .O(N__82730),
            .I(N__82724));
    Span4Mux_h I__19696 (
            .O(N__82727),
            .I(N__82721));
    Odrv4 I__19695 (
            .O(N__82724),
            .I(\pid_front.error_d_regZ0Z_14 ));
    Odrv4 I__19694 (
            .O(N__82721),
            .I(\pid_front.error_d_regZ0Z_14 ));
    InMux I__19693 (
            .O(N__82716),
            .I(N__82713));
    LocalMux I__19692 (
            .O(N__82713),
            .I(N__82709));
    InMux I__19691 (
            .O(N__82712),
            .I(N__82706));
    Span12Mux_v I__19690 (
            .O(N__82709),
            .I(N__82703));
    LocalMux I__19689 (
            .O(N__82706),
            .I(N__82700));
    Span12Mux_h I__19688 (
            .O(N__82703),
            .I(N__82697));
    Odrv4 I__19687 (
            .O(N__82700),
            .I(xy_kp_1));
    Odrv12 I__19686 (
            .O(N__82697),
            .I(xy_kp_1));
    CEMux I__19685 (
            .O(N__82692),
            .I(N__82689));
    LocalMux I__19684 (
            .O(N__82689),
            .I(N__82685));
    CEMux I__19683 (
            .O(N__82688),
            .I(N__82682));
    Span4Mux_h I__19682 (
            .O(N__82685),
            .I(N__82679));
    LocalMux I__19681 (
            .O(N__82682),
            .I(N__82676));
    Span4Mux_h I__19680 (
            .O(N__82679),
            .I(N__82672));
    Span4Mux_h I__19679 (
            .O(N__82676),
            .I(N__82669));
    CEMux I__19678 (
            .O(N__82675),
            .I(N__82666));
    Span4Mux_h I__19677 (
            .O(N__82672),
            .I(N__82659));
    Span4Mux_v I__19676 (
            .O(N__82669),
            .I(N__82659));
    LocalMux I__19675 (
            .O(N__82666),
            .I(N__82659));
    Span4Mux_h I__19674 (
            .O(N__82659),
            .I(N__82656));
    Span4Mux_h I__19673 (
            .O(N__82656),
            .I(N__82653));
    Odrv4 I__19672 (
            .O(N__82653),
            .I(\Commands_frame_decoder.state_RNIG48SZ0Z_7 ));
    InMux I__19671 (
            .O(N__82650),
            .I(N__82646));
    InMux I__19670 (
            .O(N__82649),
            .I(N__82643));
    LocalMux I__19669 (
            .O(N__82646),
            .I(N__82640));
    LocalMux I__19668 (
            .O(N__82643),
            .I(N__82637));
    Span4Mux_v I__19667 (
            .O(N__82640),
            .I(N__82632));
    Span4Mux_v I__19666 (
            .O(N__82637),
            .I(N__82632));
    Span4Mux_h I__19665 (
            .O(N__82632),
            .I(N__82629));
    Odrv4 I__19664 (
            .O(N__82629),
            .I(\pid_side.error_d_reg_prev_esr_RNIB1JOZ0Z_16 ));
    InMux I__19663 (
            .O(N__82626),
            .I(N__82622));
    InMux I__19662 (
            .O(N__82625),
            .I(N__82619));
    LocalMux I__19661 (
            .O(N__82622),
            .I(N__82614));
    LocalMux I__19660 (
            .O(N__82619),
            .I(N__82614));
    Span12Mux_v I__19659 (
            .O(N__82614),
            .I(N__82611));
    Odrv12 I__19658 (
            .O(N__82611),
            .I(\pid_side.error_d_reg_prev_esr_RNIE4JO_0Z0Z_17 ));
    InMux I__19657 (
            .O(N__82608),
            .I(N__82604));
    InMux I__19656 (
            .O(N__82607),
            .I(N__82601));
    LocalMux I__19655 (
            .O(N__82604),
            .I(\pid_side.error_p_reg_esr_RNICBEQ_0Z0Z_2 ));
    LocalMux I__19654 (
            .O(N__82601),
            .I(\pid_side.error_p_reg_esr_RNICBEQ_0Z0Z_2 ));
    InMux I__19653 (
            .O(N__82596),
            .I(N__82593));
    LocalMux I__19652 (
            .O(N__82593),
            .I(N__82590));
    Span4Mux_h I__19651 (
            .O(N__82590),
            .I(N__82587));
    Odrv4 I__19650 (
            .O(N__82587),
            .I(\pid_side.O_0_2 ));
    InMux I__19649 (
            .O(N__82584),
            .I(N__82580));
    InMux I__19648 (
            .O(N__82583),
            .I(N__82577));
    LocalMux I__19647 (
            .O(N__82580),
            .I(N__82574));
    LocalMux I__19646 (
            .O(N__82577),
            .I(N__82571));
    Span4Mux_v I__19645 (
            .O(N__82574),
            .I(N__82566));
    Span4Mux_v I__19644 (
            .O(N__82571),
            .I(N__82566));
    Span4Mux_h I__19643 (
            .O(N__82566),
            .I(N__82560));
    InMux I__19642 (
            .O(N__82565),
            .I(N__82553));
    InMux I__19641 (
            .O(N__82564),
            .I(N__82553));
    InMux I__19640 (
            .O(N__82563),
            .I(N__82553));
    Odrv4 I__19639 (
            .O(N__82560),
            .I(\pid_side.error_d_regZ0Z_0 ));
    LocalMux I__19638 (
            .O(N__82553),
            .I(\pid_side.error_d_regZ0Z_0 ));
    InMux I__19637 (
            .O(N__82548),
            .I(N__82545));
    LocalMux I__19636 (
            .O(N__82545),
            .I(N__82542));
    Span4Mux_v I__19635 (
            .O(N__82542),
            .I(N__82539));
    Odrv4 I__19634 (
            .O(N__82539),
            .I(\pid_side.O_1_5 ));
    InMux I__19633 (
            .O(N__82536),
            .I(N__82527));
    InMux I__19632 (
            .O(N__82535),
            .I(N__82527));
    InMux I__19631 (
            .O(N__82534),
            .I(N__82527));
    LocalMux I__19630 (
            .O(N__82527),
            .I(\pid_side.error_d_regZ0Z_3 ));
    InMux I__19629 (
            .O(N__82524),
            .I(N__82521));
    LocalMux I__19628 (
            .O(N__82521),
            .I(N__82518));
    Span4Mux_v I__19627 (
            .O(N__82518),
            .I(N__82515));
    Odrv4 I__19626 (
            .O(N__82515),
            .I(\pid_side.O_2_5 ));
    InMux I__19625 (
            .O(N__82512),
            .I(N__82508));
    CascadeMux I__19624 (
            .O(N__82511),
            .I(N__82505));
    LocalMux I__19623 (
            .O(N__82508),
            .I(N__82500));
    InMux I__19622 (
            .O(N__82505),
            .I(N__82493));
    InMux I__19621 (
            .O(N__82504),
            .I(N__82493));
    InMux I__19620 (
            .O(N__82503),
            .I(N__82493));
    Span4Mux_v I__19619 (
            .O(N__82500),
            .I(N__82488));
    LocalMux I__19618 (
            .O(N__82493),
            .I(N__82488));
    Span4Mux_h I__19617 (
            .O(N__82488),
            .I(N__82485));
    Odrv4 I__19616 (
            .O(N__82485),
            .I(\pid_side.error_d_reg_prevZ0Z_1 ));
    CascadeMux I__19615 (
            .O(N__82482),
            .I(N__82477));
    InMux I__19614 (
            .O(N__82481),
            .I(N__82474));
    InMux I__19613 (
            .O(N__82480),
            .I(N__82469));
    InMux I__19612 (
            .O(N__82477),
            .I(N__82469));
    LocalMux I__19611 (
            .O(N__82474),
            .I(\pid_side.error_p_regZ0Z_1 ));
    LocalMux I__19610 (
            .O(N__82469),
            .I(\pid_side.error_p_regZ0Z_1 ));
    InMux I__19609 (
            .O(N__82464),
            .I(N__82461));
    LocalMux I__19608 (
            .O(N__82461),
            .I(N__82458));
    Span4Mux_v I__19607 (
            .O(N__82458),
            .I(N__82455));
    Span4Mux_h I__19606 (
            .O(N__82455),
            .I(N__82452));
    Odrv4 I__19605 (
            .O(N__82452),
            .I(\pid_side.un1_pid_prereg_9_0 ));
    InMux I__19604 (
            .O(N__82449),
            .I(N__82446));
    LocalMux I__19603 (
            .O(N__82446),
            .I(N__82442));
    InMux I__19602 (
            .O(N__82445),
            .I(N__82439));
    Sp12to4 I__19601 (
            .O(N__82442),
            .I(N__82435));
    LocalMux I__19600 (
            .O(N__82439),
            .I(N__82432));
    InMux I__19599 (
            .O(N__82438),
            .I(N__82429));
    Odrv12 I__19598 (
            .O(N__82435),
            .I(\pid_side.error_d_regZ0Z_2 ));
    Odrv4 I__19597 (
            .O(N__82432),
            .I(\pid_side.error_d_regZ0Z_2 ));
    LocalMux I__19596 (
            .O(N__82429),
            .I(\pid_side.error_d_regZ0Z_2 ));
    InMux I__19595 (
            .O(N__82422),
            .I(N__82418));
    InMux I__19594 (
            .O(N__82421),
            .I(N__82415));
    LocalMux I__19593 (
            .O(N__82418),
            .I(\pid_side.error_p_regZ0Z_2 ));
    LocalMux I__19592 (
            .O(N__82415),
            .I(\pid_side.error_p_regZ0Z_2 ));
    InMux I__19591 (
            .O(N__82410),
            .I(N__82407));
    LocalMux I__19590 (
            .O(N__82407),
            .I(N__82403));
    InMux I__19589 (
            .O(N__82406),
            .I(N__82400));
    Span4Mux_h I__19588 (
            .O(N__82403),
            .I(N__82397));
    LocalMux I__19587 (
            .O(N__82400),
            .I(N__82394));
    Span4Mux_h I__19586 (
            .O(N__82397),
            .I(N__82391));
    Span4Mux_h I__19585 (
            .O(N__82394),
            .I(N__82388));
    Span4Mux_h I__19584 (
            .O(N__82391),
            .I(N__82385));
    Span4Mux_h I__19583 (
            .O(N__82388),
            .I(N__82382));
    Odrv4 I__19582 (
            .O(N__82385),
            .I(\pid_side.error_d_reg_prevZ0Z_2 ));
    Odrv4 I__19581 (
            .O(N__82382),
            .I(\pid_side.error_d_reg_prevZ0Z_2 ));
    InMux I__19580 (
            .O(N__82377),
            .I(N__82371));
    InMux I__19579 (
            .O(N__82376),
            .I(N__82371));
    LocalMux I__19578 (
            .O(N__82371),
            .I(\pid_side.error_p_reg_esr_RNICBEQZ0Z_2 ));
    InMux I__19577 (
            .O(N__82368),
            .I(N__82365));
    LocalMux I__19576 (
            .O(N__82365),
            .I(N__82362));
    Span4Mux_h I__19575 (
            .O(N__82362),
            .I(N__82359));
    Span4Mux_h I__19574 (
            .O(N__82359),
            .I(N__82356));
    Odrv4 I__19573 (
            .O(N__82356),
            .I(\pid_side.state_RNINK4UZ0Z_0 ));
    InMux I__19572 (
            .O(N__82353),
            .I(N__82350));
    LocalMux I__19571 (
            .O(N__82350),
            .I(N__82347));
    Span4Mux_h I__19570 (
            .O(N__82347),
            .I(N__82344));
    Odrv4 I__19569 (
            .O(N__82344),
            .I(\pid_side.O_2_14 ));
    CascadeMux I__19568 (
            .O(N__82341),
            .I(N__82336));
    CascadeMux I__19567 (
            .O(N__82340),
            .I(N__82333));
    CascadeMux I__19566 (
            .O(N__82339),
            .I(N__82329));
    InMux I__19565 (
            .O(N__82336),
            .I(N__82321));
    InMux I__19564 (
            .O(N__82333),
            .I(N__82321));
    InMux I__19563 (
            .O(N__82332),
            .I(N__82321));
    InMux I__19562 (
            .O(N__82329),
            .I(N__82316));
    InMux I__19561 (
            .O(N__82328),
            .I(N__82316));
    LocalMux I__19560 (
            .O(N__82321),
            .I(\pid_side.error_p_regZ0Z_11 ));
    LocalMux I__19559 (
            .O(N__82316),
            .I(\pid_side.error_p_regZ0Z_11 ));
    InMux I__19558 (
            .O(N__82311),
            .I(N__82308));
    LocalMux I__19557 (
            .O(N__82308),
            .I(N__82305));
    Span4Mux_h I__19556 (
            .O(N__82305),
            .I(N__82302));
    Odrv4 I__19555 (
            .O(N__82302),
            .I(\pid_side.O_1_17 ));
    InMux I__19554 (
            .O(N__82299),
            .I(N__82290));
    InMux I__19553 (
            .O(N__82298),
            .I(N__82290));
    InMux I__19552 (
            .O(N__82297),
            .I(N__82290));
    LocalMux I__19551 (
            .O(N__82290),
            .I(N__82287));
    Odrv4 I__19550 (
            .O(N__82287),
            .I(\pid_side.error_d_regZ0Z_15 ));
    InMux I__19549 (
            .O(N__82284),
            .I(N__82281));
    LocalMux I__19548 (
            .O(N__82281),
            .I(\pid_side.N_5_1 ));
    CascadeMux I__19547 (
            .O(N__82278),
            .I(N__82274));
    InMux I__19546 (
            .O(N__82277),
            .I(N__82266));
    InMux I__19545 (
            .O(N__82274),
            .I(N__82261));
    InMux I__19544 (
            .O(N__82273),
            .I(N__82261));
    CascadeMux I__19543 (
            .O(N__82272),
            .I(N__82258));
    InMux I__19542 (
            .O(N__82271),
            .I(N__82254));
    InMux I__19541 (
            .O(N__82270),
            .I(N__82251));
    InMux I__19540 (
            .O(N__82269),
            .I(N__82248));
    LocalMux I__19539 (
            .O(N__82266),
            .I(N__82243));
    LocalMux I__19538 (
            .O(N__82261),
            .I(N__82243));
    InMux I__19537 (
            .O(N__82258),
            .I(N__82238));
    InMux I__19536 (
            .O(N__82257),
            .I(N__82238));
    LocalMux I__19535 (
            .O(N__82254),
            .I(\pid_side.error_d_reg_prevZ0Z_12 ));
    LocalMux I__19534 (
            .O(N__82251),
            .I(\pid_side.error_d_reg_prevZ0Z_12 ));
    LocalMux I__19533 (
            .O(N__82248),
            .I(\pid_side.error_d_reg_prevZ0Z_12 ));
    Odrv4 I__19532 (
            .O(N__82243),
            .I(\pid_side.error_d_reg_prevZ0Z_12 ));
    LocalMux I__19531 (
            .O(N__82238),
            .I(\pid_side.error_d_reg_prevZ0Z_12 ));
    InMux I__19530 (
            .O(N__82227),
            .I(N__82223));
    InMux I__19529 (
            .O(N__82226),
            .I(N__82220));
    LocalMux I__19528 (
            .O(N__82223),
            .I(\pid_side.error_d_reg_fast_esr_RNIEIJH2Z0Z_12 ));
    LocalMux I__19527 (
            .O(N__82220),
            .I(\pid_side.error_d_reg_fast_esr_RNIEIJH2Z0Z_12 ));
    InMux I__19526 (
            .O(N__82215),
            .I(N__82212));
    LocalMux I__19525 (
            .O(N__82212),
            .I(N__82209));
    Span4Mux_h I__19524 (
            .O(N__82209),
            .I(N__82206));
    Span4Mux_v I__19523 (
            .O(N__82206),
            .I(N__82203));
    Odrv4 I__19522 (
            .O(N__82203),
            .I(\pid_side.error_d_reg_prev_esr_RNI41F23Z0Z_12 ));
    InMux I__19521 (
            .O(N__82200),
            .I(N__82196));
    InMux I__19520 (
            .O(N__82199),
            .I(N__82193));
    LocalMux I__19519 (
            .O(N__82196),
            .I(N__82190));
    LocalMux I__19518 (
            .O(N__82193),
            .I(N__82187));
    Span4Mux_v I__19517 (
            .O(N__82190),
            .I(N__82182));
    Span4Mux_h I__19516 (
            .O(N__82187),
            .I(N__82182));
    Odrv4 I__19515 (
            .O(N__82182),
            .I(\pid_side.error_d_reg_prev_esr_RNI9BFR3Z0Z_1 ));
    CascadeMux I__19514 (
            .O(N__82179),
            .I(\pid_side.error_p_reg_esr_RNIIQL11_0Z0Z_1_cascade_ ));
    InMux I__19513 (
            .O(N__82176),
            .I(N__82173));
    LocalMux I__19512 (
            .O(N__82173),
            .I(\pid_side.error_d_reg_prev_esr_RNIBGIE2Z0Z_1 ));
    InMux I__19511 (
            .O(N__82170),
            .I(N__82167));
    LocalMux I__19510 (
            .O(N__82167),
            .I(N__82163));
    CascadeMux I__19509 (
            .O(N__82166),
            .I(N__82159));
    Span4Mux_v I__19508 (
            .O(N__82163),
            .I(N__82156));
    InMux I__19507 (
            .O(N__82162),
            .I(N__82153));
    InMux I__19506 (
            .O(N__82159),
            .I(N__82150));
    Span4Mux_h I__19505 (
            .O(N__82156),
            .I(N__82147));
    LocalMux I__19504 (
            .O(N__82153),
            .I(N__82144));
    LocalMux I__19503 (
            .O(N__82150),
            .I(N__82141));
    Odrv4 I__19502 (
            .O(N__82147),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_1_c_RNI0LLN ));
    Odrv4 I__19501 (
            .O(N__82144),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_1_c_RNI0LLN ));
    Odrv4 I__19500 (
            .O(N__82141),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_1_c_RNI0LLN ));
    CascadeMux I__19499 (
            .O(N__82134),
            .I(\pid_side.error_d_reg_prev_esr_RNIBGIE2Z0Z_1_cascade_ ));
    InMux I__19498 (
            .O(N__82131),
            .I(N__82128));
    LocalMux I__19497 (
            .O(N__82128),
            .I(N__82125));
    Odrv12 I__19496 (
            .O(N__82125),
            .I(\pid_side.error_d_reg_prev_esr_RNI905J4Z0Z_1 ));
    InMux I__19495 (
            .O(N__82122),
            .I(N__82119));
    LocalMux I__19494 (
            .O(N__82119),
            .I(\pid_side.error_p_reg_esr_RNIIQL11Z0Z_1 ));
    InMux I__19493 (
            .O(N__82116),
            .I(N__82113));
    LocalMux I__19492 (
            .O(N__82113),
            .I(\pid_side.error_d_reg_prev_esr_RNIIFEIZ0Z_1 ));
    InMux I__19491 (
            .O(N__82110),
            .I(N__82106));
    InMux I__19490 (
            .O(N__82109),
            .I(N__82103));
    LocalMux I__19489 (
            .O(N__82106),
            .I(N__82099));
    LocalMux I__19488 (
            .O(N__82103),
            .I(N__82096));
    CascadeMux I__19487 (
            .O(N__82102),
            .I(N__82093));
    Span4Mux_h I__19486 (
            .O(N__82099),
            .I(N__82087));
    Span4Mux_v I__19485 (
            .O(N__82096),
            .I(N__82087));
    InMux I__19484 (
            .O(N__82093),
            .I(N__82082));
    InMux I__19483 (
            .O(N__82092),
            .I(N__82082));
    Odrv4 I__19482 (
            .O(N__82087),
            .I(\pid_side.error_d_reg_prevZ0Z_0 ));
    LocalMux I__19481 (
            .O(N__82082),
            .I(\pid_side.error_d_reg_prevZ0Z_0 ));
    InMux I__19480 (
            .O(N__82077),
            .I(N__82071));
    InMux I__19479 (
            .O(N__82076),
            .I(N__82066));
    InMux I__19478 (
            .O(N__82075),
            .I(N__82066));
    InMux I__19477 (
            .O(N__82074),
            .I(N__82063));
    LocalMux I__19476 (
            .O(N__82071),
            .I(\pid_side.un1_pid_prereg_135_0 ));
    LocalMux I__19475 (
            .O(N__82066),
            .I(\pid_side.un1_pid_prereg_135_0 ));
    LocalMux I__19474 (
            .O(N__82063),
            .I(\pid_side.un1_pid_prereg_135_0 ));
    CascadeMux I__19473 (
            .O(N__82056),
            .I(\pid_side.N_3_i_1_1_cascade_ ));
    InMux I__19472 (
            .O(N__82053),
            .I(N__82048));
    InMux I__19471 (
            .O(N__82052),
            .I(N__82045));
    InMux I__19470 (
            .O(N__82051),
            .I(N__82042));
    LocalMux I__19469 (
            .O(N__82048),
            .I(\pid_side.un1_pid_prereg_79 ));
    LocalMux I__19468 (
            .O(N__82045),
            .I(\pid_side.un1_pid_prereg_79 ));
    LocalMux I__19467 (
            .O(N__82042),
            .I(\pid_side.un1_pid_prereg_79 ));
    InMux I__19466 (
            .O(N__82035),
            .I(N__82032));
    LocalMux I__19465 (
            .O(N__82032),
            .I(N__82029));
    Odrv4 I__19464 (
            .O(N__82029),
            .I(\pid_side.N_5_0 ));
    CascadeMux I__19463 (
            .O(N__82026),
            .I(\pid_side.N_3_i_1_cascade_ ));
    InMux I__19462 (
            .O(N__82023),
            .I(N__82018));
    InMux I__19461 (
            .O(N__82022),
            .I(N__82015));
    InMux I__19460 (
            .O(N__82021),
            .I(N__82012));
    LocalMux I__19459 (
            .O(N__82018),
            .I(N__82009));
    LocalMux I__19458 (
            .O(N__82015),
            .I(N__82006));
    LocalMux I__19457 (
            .O(N__82012),
            .I(N__82003));
    Span4Mux_v I__19456 (
            .O(N__82009),
            .I(N__82000));
    Span4Mux_h I__19455 (
            .O(N__82006),
            .I(N__81997));
    Span4Mux_v I__19454 (
            .O(N__82003),
            .I(N__81994));
    Span4Mux_h I__19453 (
            .O(N__82000),
            .I(N__81989));
    Span4Mux_h I__19452 (
            .O(N__81997),
            .I(N__81989));
    Odrv4 I__19451 (
            .O(N__81994),
            .I(\pid_side.error_i_reg_esr_RNIO6NRZ0Z_14 ));
    Odrv4 I__19450 (
            .O(N__81989),
            .I(\pid_side.error_i_reg_esr_RNIO6NRZ0Z_14 ));
    InMux I__19449 (
            .O(N__81984),
            .I(N__81979));
    InMux I__19448 (
            .O(N__81983),
            .I(N__81976));
    InMux I__19447 (
            .O(N__81982),
            .I(N__81972));
    LocalMux I__19446 (
            .O(N__81979),
            .I(N__81969));
    LocalMux I__19445 (
            .O(N__81976),
            .I(N__81966));
    InMux I__19444 (
            .O(N__81975),
            .I(N__81963));
    LocalMux I__19443 (
            .O(N__81972),
            .I(N__81960));
    Span4Mux_v I__19442 (
            .O(N__81969),
            .I(N__81957));
    Span4Mux_v I__19441 (
            .O(N__81966),
            .I(N__81952));
    LocalMux I__19440 (
            .O(N__81963),
            .I(N__81952));
    Span4Mux_v I__19439 (
            .O(N__81960),
            .I(N__81949));
    Span4Mux_h I__19438 (
            .O(N__81957),
            .I(N__81944));
    Span4Mux_v I__19437 (
            .O(N__81952),
            .I(N__81944));
    Odrv4 I__19436 (
            .O(N__81949),
            .I(\pid_side.error_i_reg_esr_RNIM3MRZ0Z_13 ));
    Odrv4 I__19435 (
            .O(N__81944),
            .I(\pid_side.error_i_reg_esr_RNIM3MRZ0Z_13 ));
    CascadeMux I__19434 (
            .O(N__81939),
            .I(\pid_side.error_d_reg_prev_esr_RNIQTGL4Z0Z_12_cascade_ ));
    InMux I__19433 (
            .O(N__81936),
            .I(N__81933));
    LocalMux I__19432 (
            .O(N__81933),
            .I(\pid_side.error_d_reg_prev_esr_RNI6P1R3Z0Z_12 ));
    InMux I__19431 (
            .O(N__81930),
            .I(N__81927));
    LocalMux I__19430 (
            .O(N__81927),
            .I(N__81923));
    InMux I__19429 (
            .O(N__81926),
            .I(N__81920));
    Span4Mux_h I__19428 (
            .O(N__81923),
            .I(N__81915));
    LocalMux I__19427 (
            .O(N__81920),
            .I(N__81915));
    Span4Mux_h I__19426 (
            .O(N__81915),
            .I(N__81912));
    Span4Mux_v I__19425 (
            .O(N__81912),
            .I(N__81909));
    Odrv4 I__19424 (
            .O(N__81909),
            .I(\pid_side.un1_pid_prereg_0_axb_14 ));
    InMux I__19423 (
            .O(N__81906),
            .I(N__81903));
    LocalMux I__19422 (
            .O(N__81903),
            .I(N__81897));
    InMux I__19421 (
            .O(N__81902),
            .I(N__81894));
    InMux I__19420 (
            .O(N__81901),
            .I(N__81889));
    InMux I__19419 (
            .O(N__81900),
            .I(N__81889));
    Odrv4 I__19418 (
            .O(N__81897),
            .I(\pid_side.error_d_reg_prev_fastZ0Z_12 ));
    LocalMux I__19417 (
            .O(N__81894),
            .I(\pid_side.error_d_reg_prev_fastZ0Z_12 ));
    LocalMux I__19416 (
            .O(N__81889),
            .I(\pid_side.error_d_reg_prev_fastZ0Z_12 ));
    CascadeMux I__19415 (
            .O(N__81882),
            .I(\pid_side.g1_1_cascade_ ));
    InMux I__19414 (
            .O(N__81879),
            .I(N__81876));
    LocalMux I__19413 (
            .O(N__81876),
            .I(N__81873));
    Odrv4 I__19412 (
            .O(N__81873),
            .I(\pid_side.g0_3_2 ));
    InMux I__19411 (
            .O(N__81870),
            .I(N__81866));
    InMux I__19410 (
            .O(N__81869),
            .I(N__81861));
    LocalMux I__19409 (
            .O(N__81866),
            .I(N__81858));
    InMux I__19408 (
            .O(N__81865),
            .I(N__81853));
    InMux I__19407 (
            .O(N__81864),
            .I(N__81853));
    LocalMux I__19406 (
            .O(N__81861),
            .I(\pid_side.error_d_reg_fastZ0Z_12 ));
    Odrv4 I__19405 (
            .O(N__81858),
            .I(\pid_side.error_d_reg_fastZ0Z_12 ));
    LocalMux I__19404 (
            .O(N__81853),
            .I(\pid_side.error_d_reg_fastZ0Z_12 ));
    CascadeMux I__19403 (
            .O(N__81846),
            .I(\pid_side.N_2398_i_cascade_ ));
    InMux I__19402 (
            .O(N__81843),
            .I(N__81837));
    InMux I__19401 (
            .O(N__81842),
            .I(N__81837));
    LocalMux I__19400 (
            .O(N__81837),
            .I(N__81834));
    Odrv4 I__19399 (
            .O(N__81834),
            .I(\pid_side.error_p_reg_esr_RNIL0VP1Z0Z_12 ));
    InMux I__19398 (
            .O(N__81831),
            .I(N__81820));
    InMux I__19397 (
            .O(N__81830),
            .I(N__81820));
    InMux I__19396 (
            .O(N__81829),
            .I(N__81820));
    InMux I__19395 (
            .O(N__81828),
            .I(N__81815));
    InMux I__19394 (
            .O(N__81827),
            .I(N__81815));
    LocalMux I__19393 (
            .O(N__81820),
            .I(\pid_side.error_d_reg_prevZ0Z_11 ));
    LocalMux I__19392 (
            .O(N__81815),
            .I(\pid_side.error_d_reg_prevZ0Z_11 ));
    InMux I__19391 (
            .O(N__81810),
            .I(N__81807));
    LocalMux I__19390 (
            .O(N__81807),
            .I(\pid_side.N_2398_i ));
    CascadeMux I__19389 (
            .O(N__81804),
            .I(\pid_side.un1_pid_prereg_79_cascade_ ));
    CascadeMux I__19388 (
            .O(N__81801),
            .I(\pid_side.un1_pid_prereg_167_0_1_cascade_ ));
    InMux I__19387 (
            .O(N__81798),
            .I(N__81795));
    LocalMux I__19386 (
            .O(N__81795),
            .I(\pid_side.un1_pid_prereg_167_0 ));
    InMux I__19385 (
            .O(N__81792),
            .I(N__81789));
    LocalMux I__19384 (
            .O(N__81789),
            .I(N__81786));
    Odrv4 I__19383 (
            .O(N__81786),
            .I(\pid_side.g0_19_1_1 ));
    InMux I__19382 (
            .O(N__81783),
            .I(N__81780));
    LocalMux I__19381 (
            .O(N__81780),
            .I(\pid_side.g0_19_1 ));
    InMux I__19380 (
            .O(N__81777),
            .I(N__81770));
    InMux I__19379 (
            .O(N__81776),
            .I(N__81770));
    InMux I__19378 (
            .O(N__81775),
            .I(N__81767));
    LocalMux I__19377 (
            .O(N__81770),
            .I(N__81764));
    LocalMux I__19376 (
            .O(N__81767),
            .I(N__81761));
    Span4Mux_h I__19375 (
            .O(N__81764),
            .I(N__81758));
    Odrv12 I__19374 (
            .O(N__81761),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_2_c_RNI3PMN ));
    Odrv4 I__19373 (
            .O(N__81758),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_2_c_RNI3PMN ));
    CascadeMux I__19372 (
            .O(N__81753),
            .I(\pid_side.error_p_reg_esr_RNIFEEQ_0Z0Z_3_cascade_ ));
    CascadeMux I__19371 (
            .O(N__81750),
            .I(N__81747));
    InMux I__19370 (
            .O(N__81747),
            .I(N__81744));
    LocalMux I__19369 (
            .O(N__81744),
            .I(N__81741));
    Span4Mux_v I__19368 (
            .O(N__81741),
            .I(N__81738));
    Odrv4 I__19367 (
            .O(N__81738),
            .I(\pid_side.error_p_reg_esr_RNI7U286Z0Z_2 ));
    InMux I__19366 (
            .O(N__81735),
            .I(N__81731));
    InMux I__19365 (
            .O(N__81734),
            .I(N__81728));
    LocalMux I__19364 (
            .O(N__81731),
            .I(N__81725));
    LocalMux I__19363 (
            .O(N__81728),
            .I(N__81722));
    Span4Mux_h I__19362 (
            .O(N__81725),
            .I(N__81719));
    Span4Mux_h I__19361 (
            .O(N__81722),
            .I(N__81716));
    Odrv4 I__19360 (
            .O(N__81719),
            .I(\pid_side.error_d_reg_prev_esr_RNIKAJO_0Z0Z_19 ));
    Odrv4 I__19359 (
            .O(N__81716),
            .I(\pid_side.error_d_reg_prev_esr_RNIKAJO_0Z0Z_19 ));
    InMux I__19358 (
            .O(N__81711),
            .I(N__81705));
    InMux I__19357 (
            .O(N__81710),
            .I(N__81705));
    LocalMux I__19356 (
            .O(N__81705),
            .I(\pid_side.error_d_reg_prevZ0Z_19 ));
    InMux I__19355 (
            .O(N__81702),
            .I(N__81699));
    LocalMux I__19354 (
            .O(N__81699),
            .I(N__81695));
    InMux I__19353 (
            .O(N__81698),
            .I(N__81692));
    Span4Mux_v I__19352 (
            .O(N__81695),
            .I(N__81687));
    LocalMux I__19351 (
            .O(N__81692),
            .I(N__81687));
    Odrv4 I__19350 (
            .O(N__81687),
            .I(\pid_side.error_d_reg_prev_esr_RNIKAJOZ0Z_19 ));
    InMux I__19349 (
            .O(N__81684),
            .I(N__81681));
    LocalMux I__19348 (
            .O(N__81681),
            .I(N__81678));
    Span4Mux_h I__19347 (
            .O(N__81678),
            .I(N__81675));
    Odrv4 I__19346 (
            .O(N__81675),
            .I(\pid_side.g0_1_0 ));
    InMux I__19345 (
            .O(N__81672),
            .I(N__81666));
    InMux I__19344 (
            .O(N__81671),
            .I(N__81666));
    LocalMux I__19343 (
            .O(N__81666),
            .I(N__81663));
    Span4Mux_h I__19342 (
            .O(N__81663),
            .I(N__81660));
    Odrv4 I__19341 (
            .O(N__81660),
            .I(\pid_side.error_d_reg_prev_esr_RNISHIO_1Z0Z_11 ));
    InMux I__19340 (
            .O(N__81657),
            .I(N__81654));
    LocalMux I__19339 (
            .O(N__81654),
            .I(N__81650));
    InMux I__19338 (
            .O(N__81653),
            .I(N__81647));
    Span4Mux_v I__19337 (
            .O(N__81650),
            .I(N__81642));
    LocalMux I__19336 (
            .O(N__81647),
            .I(N__81642));
    Odrv4 I__19335 (
            .O(N__81642),
            .I(\pid_side.error_d_reg_prev_esr_RNISKLO_0Z0Z_20 ));
    InMux I__19334 (
            .O(N__81639),
            .I(N__81636));
    LocalMux I__19333 (
            .O(N__81636),
            .I(N__81633));
    Span4Mux_v I__19332 (
            .O(N__81633),
            .I(N__81630));
    Odrv4 I__19331 (
            .O(N__81630),
            .I(\pid_side.O_2_13 ));
    InMux I__19330 (
            .O(N__81627),
            .I(N__81623));
    CascadeMux I__19329 (
            .O(N__81626),
            .I(N__81620));
    LocalMux I__19328 (
            .O(N__81623),
            .I(N__81616));
    InMux I__19327 (
            .O(N__81620),
            .I(N__81611));
    InMux I__19326 (
            .O(N__81619),
            .I(N__81611));
    Odrv12 I__19325 (
            .O(N__81616),
            .I(\pid_side.error_p_regZ0Z_10 ));
    LocalMux I__19324 (
            .O(N__81611),
            .I(\pid_side.error_p_regZ0Z_10 ));
    InMux I__19323 (
            .O(N__81606),
            .I(N__81602));
    InMux I__19322 (
            .O(N__81605),
            .I(N__81599));
    LocalMux I__19321 (
            .O(N__81602),
            .I(N__81596));
    LocalMux I__19320 (
            .O(N__81599),
            .I(N__81593));
    Odrv4 I__19319 (
            .O(N__81596),
            .I(\pid_side.error_p_reg_esr_RNIG7MC2_0Z0Z_5 ));
    Odrv12 I__19318 (
            .O(N__81593),
            .I(\pid_side.error_p_reg_esr_RNIG7MC2_0Z0Z_5 ));
    CascadeMux I__19317 (
            .O(N__81588),
            .I(\pid_side.error_p_reg_esr_RNIFEEQZ0Z_3_cascade_ ));
    CascadeMux I__19316 (
            .O(N__81585),
            .I(N__81582));
    InMux I__19315 (
            .O(N__81582),
            .I(N__81579));
    LocalMux I__19314 (
            .O(N__81579),
            .I(N__81576));
    Span4Mux_v I__19313 (
            .O(N__81576),
            .I(N__81573));
    Span4Mux_h I__19312 (
            .O(N__81573),
            .I(N__81570));
    Odrv4 I__19311 (
            .O(N__81570),
            .I(\pid_side.error_p_reg_esr_RNIN4BP4Z0Z_3 ));
    InMux I__19310 (
            .O(N__81567),
            .I(N__81564));
    LocalMux I__19309 (
            .O(N__81564),
            .I(N__81560));
    InMux I__19308 (
            .O(N__81563),
            .I(N__81557));
    Odrv12 I__19307 (
            .O(N__81560),
            .I(\pid_side.error_p_regZ0Z_4 ));
    LocalMux I__19306 (
            .O(N__81557),
            .I(\pid_side.error_p_regZ0Z_4 ));
    InMux I__19305 (
            .O(N__81552),
            .I(N__81549));
    LocalMux I__19304 (
            .O(N__81549),
            .I(N__81545));
    InMux I__19303 (
            .O(N__81548),
            .I(N__81542));
    Span4Mux_v I__19302 (
            .O(N__81545),
            .I(N__81537));
    LocalMux I__19301 (
            .O(N__81542),
            .I(N__81537));
    Span4Mux_h I__19300 (
            .O(N__81537),
            .I(N__81534));
    Odrv4 I__19299 (
            .O(N__81534),
            .I(\pid_side.error_d_reg_prevZ0Z_4 ));
    InMux I__19298 (
            .O(N__81531),
            .I(N__81528));
    LocalMux I__19297 (
            .O(N__81528),
            .I(N__81525));
    Span4Mux_h I__19296 (
            .O(N__81525),
            .I(N__81521));
    InMux I__19295 (
            .O(N__81524),
            .I(N__81517));
    Span4Mux_h I__19294 (
            .O(N__81521),
            .I(N__81514));
    InMux I__19293 (
            .O(N__81520),
            .I(N__81511));
    LocalMux I__19292 (
            .O(N__81517),
            .I(N__81508));
    Odrv4 I__19291 (
            .O(N__81514),
            .I(\pid_side.error_d_regZ0Z_4 ));
    LocalMux I__19290 (
            .O(N__81511),
            .I(\pid_side.error_d_regZ0Z_4 ));
    Odrv4 I__19289 (
            .O(N__81508),
            .I(\pid_side.error_d_regZ0Z_4 ));
    InMux I__19288 (
            .O(N__81501),
            .I(N__81498));
    LocalMux I__19287 (
            .O(N__81498),
            .I(N__81495));
    Odrv4 I__19286 (
            .O(N__81495),
            .I(\pid_side.error_p_reg_esr_RNIIHEQ_0Z0Z_4 ));
    InMux I__19285 (
            .O(N__81492),
            .I(N__81489));
    LocalMux I__19284 (
            .O(N__81489),
            .I(\pid_side.error_p_reg_esr_RNIFEEQZ0Z_3 ));
    CascadeMux I__19283 (
            .O(N__81486),
            .I(\pid_side.error_p_reg_esr_RNIIHEQ_0Z0Z_4_cascade_ ));
    InMux I__19282 (
            .O(N__81483),
            .I(N__81478));
    InMux I__19281 (
            .O(N__81482),
            .I(N__81473));
    InMux I__19280 (
            .O(N__81481),
            .I(N__81473));
    LocalMux I__19279 (
            .O(N__81478),
            .I(N__81470));
    LocalMux I__19278 (
            .O(N__81473),
            .I(N__81467));
    Odrv4 I__19277 (
            .O(N__81470),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_3_c_RNI6TNN ));
    Odrv12 I__19276 (
            .O(N__81467),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_3_c_RNI6TNN ));
    InMux I__19275 (
            .O(N__81462),
            .I(N__81459));
    LocalMux I__19274 (
            .O(N__81459),
            .I(N__81456));
    Span4Mux_h I__19273 (
            .O(N__81456),
            .I(N__81453));
    Span4Mux_h I__19272 (
            .O(N__81453),
            .I(N__81450));
    Odrv4 I__19271 (
            .O(N__81450),
            .I(\pid_side.error_p_reg_esr_RNI5G8P4Z0Z_3 ));
    CascadeMux I__19270 (
            .O(N__81447),
            .I(N__81444));
    InMux I__19269 (
            .O(N__81444),
            .I(N__81441));
    LocalMux I__19268 (
            .O(N__81441),
            .I(N__81437));
    InMux I__19267 (
            .O(N__81440),
            .I(N__81434));
    Span4Mux_h I__19266 (
            .O(N__81437),
            .I(N__81431));
    LocalMux I__19265 (
            .O(N__81434),
            .I(\pid_side.error_p_reg_esr_RNIUIJC2Z0Z_2 ));
    Odrv4 I__19264 (
            .O(N__81431),
            .I(\pid_side.error_p_reg_esr_RNIUIJC2Z0Z_2 ));
    CascadeMux I__19263 (
            .O(N__81426),
            .I(N__81423));
    InMux I__19262 (
            .O(N__81423),
            .I(N__81417));
    InMux I__19261 (
            .O(N__81422),
            .I(N__81417));
    LocalMux I__19260 (
            .O(N__81417),
            .I(\pid_side.error_d_reg_prevZ0Z_3 ));
    InMux I__19259 (
            .O(N__81414),
            .I(N__81408));
    InMux I__19258 (
            .O(N__81413),
            .I(N__81408));
    LocalMux I__19257 (
            .O(N__81408),
            .I(N__81405));
    Odrv4 I__19256 (
            .O(N__81405),
            .I(\pid_side.error_p_regZ0Z_3 ));
    InMux I__19255 (
            .O(N__81402),
            .I(N__81399));
    LocalMux I__19254 (
            .O(N__81399),
            .I(\pid_side.error_p_reg_esr_RNIFEEQ_0Z0Z_3 ));
    InMux I__19253 (
            .O(N__81396),
            .I(N__81393));
    LocalMux I__19252 (
            .O(N__81393),
            .I(N__81390));
    Span4Mux_h I__19251 (
            .O(N__81390),
            .I(N__81387));
    Span4Mux_v I__19250 (
            .O(N__81387),
            .I(N__81384));
    Odrv4 I__19249 (
            .O(N__81384),
            .I(\pid_side.O_1_7 ));
    InMux I__19248 (
            .O(N__81381),
            .I(N__81377));
    InMux I__19247 (
            .O(N__81380),
            .I(N__81374));
    LocalMux I__19246 (
            .O(N__81377),
            .I(N__81371));
    LocalMux I__19245 (
            .O(N__81374),
            .I(N__81368));
    Span12Mux_h I__19244 (
            .O(N__81371),
            .I(N__81362));
    Span12Mux_h I__19243 (
            .O(N__81368),
            .I(N__81359));
    InMux I__19242 (
            .O(N__81367),
            .I(N__81352));
    InMux I__19241 (
            .O(N__81366),
            .I(N__81352));
    InMux I__19240 (
            .O(N__81365),
            .I(N__81352));
    Odrv12 I__19239 (
            .O(N__81362),
            .I(\pid_side.error_d_regZ0Z_5 ));
    Odrv12 I__19238 (
            .O(N__81359),
            .I(\pid_side.error_d_regZ0Z_5 ));
    LocalMux I__19237 (
            .O(N__81352),
            .I(\pid_side.error_d_regZ0Z_5 ));
    InMux I__19236 (
            .O(N__81345),
            .I(N__81342));
    LocalMux I__19235 (
            .O(N__81342),
            .I(N__81339));
    Span4Mux_h I__19234 (
            .O(N__81339),
            .I(N__81336));
    Odrv4 I__19233 (
            .O(N__81336),
            .I(\pid_side.O_2_6 ));
    InMux I__19232 (
            .O(N__81333),
            .I(N__81330));
    LocalMux I__19231 (
            .O(N__81330),
            .I(N__81327));
    Span4Mux_h I__19230 (
            .O(N__81327),
            .I(N__81324));
    Odrv4 I__19229 (
            .O(N__81324),
            .I(\pid_side.O_1_4 ));
    InMux I__19228 (
            .O(N__81321),
            .I(N__81318));
    LocalMux I__19227 (
            .O(N__81318),
            .I(N__81315));
    Span4Mux_h I__19226 (
            .O(N__81315),
            .I(N__81312));
    Odrv4 I__19225 (
            .O(N__81312),
            .I(\pid_side.O_1_12 ));
    InMux I__19224 (
            .O(N__81309),
            .I(N__81303));
    InMux I__19223 (
            .O(N__81308),
            .I(N__81303));
    LocalMux I__19222 (
            .O(N__81303),
            .I(N__81296));
    InMux I__19221 (
            .O(N__81302),
            .I(N__81287));
    InMux I__19220 (
            .O(N__81301),
            .I(N__81287));
    InMux I__19219 (
            .O(N__81300),
            .I(N__81287));
    InMux I__19218 (
            .O(N__81299),
            .I(N__81287));
    Odrv12 I__19217 (
            .O(N__81296),
            .I(\pid_side.error_d_regZ0Z_10 ));
    LocalMux I__19216 (
            .O(N__81287),
            .I(\pid_side.error_d_regZ0Z_10 ));
    InMux I__19215 (
            .O(N__81282),
            .I(N__81279));
    LocalMux I__19214 (
            .O(N__81279),
            .I(N__81276));
    Span4Mux_h I__19213 (
            .O(N__81276),
            .I(N__81273));
    Odrv4 I__19212 (
            .O(N__81273),
            .I(\pid_side.O_1_8 ));
    InMux I__19211 (
            .O(N__81270),
            .I(N__81258));
    InMux I__19210 (
            .O(N__81269),
            .I(N__81258));
    InMux I__19209 (
            .O(N__81268),
            .I(N__81258));
    InMux I__19208 (
            .O(N__81267),
            .I(N__81258));
    LocalMux I__19207 (
            .O(N__81258),
            .I(N__81255));
    Span4Mux_h I__19206 (
            .O(N__81255),
            .I(N__81252));
    Span4Mux_h I__19205 (
            .O(N__81252),
            .I(N__81249));
    Odrv4 I__19204 (
            .O(N__81249),
            .I(\pid_side.error_d_regZ0Z_6 ));
    InMux I__19203 (
            .O(N__81246),
            .I(N__81243));
    LocalMux I__19202 (
            .O(N__81243),
            .I(N__81240));
    Span4Mux_h I__19201 (
            .O(N__81240),
            .I(N__81237));
    Odrv4 I__19200 (
            .O(N__81237),
            .I(\pid_side.O_1_9 ));
    InMux I__19199 (
            .O(N__81234),
            .I(N__81230));
    InMux I__19198 (
            .O(N__81233),
            .I(N__81225));
    LocalMux I__19197 (
            .O(N__81230),
            .I(N__81222));
    InMux I__19196 (
            .O(N__81229),
            .I(N__81217));
    InMux I__19195 (
            .O(N__81228),
            .I(N__81217));
    LocalMux I__19194 (
            .O(N__81225),
            .I(N__81214));
    Span4Mux_h I__19193 (
            .O(N__81222),
            .I(N__81211));
    LocalMux I__19192 (
            .O(N__81217),
            .I(N__81208));
    Span4Mux_h I__19191 (
            .O(N__81214),
            .I(N__81205));
    Span4Mux_h I__19190 (
            .O(N__81211),
            .I(N__81202));
    Span4Mux_h I__19189 (
            .O(N__81208),
            .I(N__81199));
    Span4Mux_h I__19188 (
            .O(N__81205),
            .I(N__81196));
    Span4Mux_h I__19187 (
            .O(N__81202),
            .I(N__81193));
    Span4Mux_h I__19186 (
            .O(N__81199),
            .I(N__81188));
    Span4Mux_v I__19185 (
            .O(N__81196),
            .I(N__81188));
    Odrv4 I__19184 (
            .O(N__81193),
            .I(\pid_side.error_d_regZ0Z_7 ));
    Odrv4 I__19183 (
            .O(N__81188),
            .I(\pid_side.error_d_regZ0Z_7 ));
    InMux I__19182 (
            .O(N__81183),
            .I(N__81180));
    LocalMux I__19181 (
            .O(N__81180),
            .I(N__81177));
    Span4Mux_h I__19180 (
            .O(N__81177),
            .I(N__81174));
    Odrv4 I__19179 (
            .O(N__81174),
            .I(\pid_side.O_1_10 ));
    CascadeMux I__19178 (
            .O(N__81171),
            .I(N__81166));
    CascadeMux I__19177 (
            .O(N__81170),
            .I(N__81163));
    InMux I__19176 (
            .O(N__81169),
            .I(N__81153));
    InMux I__19175 (
            .O(N__81166),
            .I(N__81153));
    InMux I__19174 (
            .O(N__81163),
            .I(N__81153));
    InMux I__19173 (
            .O(N__81162),
            .I(N__81153));
    LocalMux I__19172 (
            .O(N__81153),
            .I(N__81150));
    Span4Mux_h I__19171 (
            .O(N__81150),
            .I(N__81147));
    Span4Mux_h I__19170 (
            .O(N__81147),
            .I(N__81144));
    Odrv4 I__19169 (
            .O(N__81144),
            .I(\pid_side.error_d_regZ0Z_8 ));
    InMux I__19168 (
            .O(N__81141),
            .I(N__81138));
    LocalMux I__19167 (
            .O(N__81138),
            .I(N__81135));
    Span4Mux_h I__19166 (
            .O(N__81135),
            .I(N__81132));
    Odrv4 I__19165 (
            .O(N__81132),
            .I(\pid_side.O_1_11 ));
    InMux I__19164 (
            .O(N__81129),
            .I(N__81120));
    InMux I__19163 (
            .O(N__81128),
            .I(N__81120));
    InMux I__19162 (
            .O(N__81127),
            .I(N__81120));
    LocalMux I__19161 (
            .O(N__81120),
            .I(N__81115));
    InMux I__19160 (
            .O(N__81119),
            .I(N__81110));
    InMux I__19159 (
            .O(N__81118),
            .I(N__81110));
    Odrv4 I__19158 (
            .O(N__81115),
            .I(\pid_side.error_d_regZ0Z_9 ));
    LocalMux I__19157 (
            .O(N__81110),
            .I(\pid_side.error_d_regZ0Z_9 ));
    InMux I__19156 (
            .O(N__81105),
            .I(N__81102));
    LocalMux I__19155 (
            .O(N__81102),
            .I(N__81099));
    Span4Mux_h I__19154 (
            .O(N__81099),
            .I(N__81096));
    Odrv4 I__19153 (
            .O(N__81096),
            .I(\pid_side.O_2_4 ));
    CascadeMux I__19152 (
            .O(N__81093),
            .I(\pid_side.N_2405_0_0_0_cascade_ ));
    CascadeMux I__19151 (
            .O(N__81090),
            .I(\pid_side.g0_2_0_cascade_ ));
    InMux I__19150 (
            .O(N__81087),
            .I(N__81084));
    LocalMux I__19149 (
            .O(N__81084),
            .I(\pid_side.error_d_reg_prev_esr_RNIQ0PB4Z0Z_12 ));
    InMux I__19148 (
            .O(N__81081),
            .I(N__81078));
    LocalMux I__19147 (
            .O(N__81078),
            .I(\pid_side.N_4_1_0_1 ));
    InMux I__19146 (
            .O(N__81075),
            .I(N__81072));
    LocalMux I__19145 (
            .O(N__81072),
            .I(N__81068));
    InMux I__19144 (
            .O(N__81071),
            .I(N__81064));
    Span4Mux_v I__19143 (
            .O(N__81068),
            .I(N__81061));
    CascadeMux I__19142 (
            .O(N__81067),
            .I(N__81054));
    LocalMux I__19141 (
            .O(N__81064),
            .I(N__81051));
    Span4Mux_s0_h I__19140 (
            .O(N__81061),
            .I(N__81048));
    InMux I__19139 (
            .O(N__81060),
            .I(N__81044));
    InMux I__19138 (
            .O(N__81059),
            .I(N__81041));
    InMux I__19137 (
            .O(N__81058),
            .I(N__81038));
    InMux I__19136 (
            .O(N__81057),
            .I(N__81035));
    InMux I__19135 (
            .O(N__81054),
            .I(N__81032));
    Span4Mux_v I__19134 (
            .O(N__81051),
            .I(N__81027));
    Span4Mux_h I__19133 (
            .O(N__81048),
            .I(N__81027));
    InMux I__19132 (
            .O(N__81047),
            .I(N__81024));
    LocalMux I__19131 (
            .O(N__81044),
            .I(N__81021));
    LocalMux I__19130 (
            .O(N__81041),
            .I(N__81018));
    LocalMux I__19129 (
            .O(N__81038),
            .I(N__81015));
    LocalMux I__19128 (
            .O(N__81035),
            .I(N__81012));
    LocalMux I__19127 (
            .O(N__81032),
            .I(N__81009));
    Span4Mux_h I__19126 (
            .O(N__81027),
            .I(N__81004));
    LocalMux I__19125 (
            .O(N__81024),
            .I(N__81004));
    Span12Mux_s0_h I__19124 (
            .O(N__81021),
            .I(N__81001));
    Span4Mux_h I__19123 (
            .O(N__81018),
            .I(N__80998));
    Span4Mux_h I__19122 (
            .O(N__81015),
            .I(N__80989));
    Span4Mux_h I__19121 (
            .O(N__81012),
            .I(N__80989));
    Span4Mux_h I__19120 (
            .O(N__81009),
            .I(N__80989));
    Span4Mux_h I__19119 (
            .O(N__81004),
            .I(N__80989));
    Odrv12 I__19118 (
            .O(N__81001),
            .I(drone_H_disp_side_0));
    Odrv4 I__19117 (
            .O(N__80998),
            .I(drone_H_disp_side_0));
    Odrv4 I__19116 (
            .O(N__80989),
            .I(drone_H_disp_side_0));
    InMux I__19115 (
            .O(N__80982),
            .I(N__80977));
    InMux I__19114 (
            .O(N__80981),
            .I(N__80968));
    CascadeMux I__19113 (
            .O(N__80980),
            .I(N__80965));
    LocalMux I__19112 (
            .O(N__80977),
            .I(N__80956));
    InMux I__19111 (
            .O(N__80976),
            .I(N__80953));
    InMux I__19110 (
            .O(N__80975),
            .I(N__80948));
    InMux I__19109 (
            .O(N__80974),
            .I(N__80948));
    CascadeMux I__19108 (
            .O(N__80973),
            .I(N__80945));
    CascadeMux I__19107 (
            .O(N__80972),
            .I(N__80940));
    CascadeMux I__19106 (
            .O(N__80971),
            .I(N__80935));
    LocalMux I__19105 (
            .O(N__80968),
            .I(N__80932));
    InMux I__19104 (
            .O(N__80965),
            .I(N__80924));
    InMux I__19103 (
            .O(N__80964),
            .I(N__80924));
    InMux I__19102 (
            .O(N__80963),
            .I(N__80924));
    InMux I__19101 (
            .O(N__80962),
            .I(N__80919));
    InMux I__19100 (
            .O(N__80961),
            .I(N__80919));
    InMux I__19099 (
            .O(N__80960),
            .I(N__80914));
    InMux I__19098 (
            .O(N__80959),
            .I(N__80914));
    Span4Mux_v I__19097 (
            .O(N__80956),
            .I(N__80907));
    LocalMux I__19096 (
            .O(N__80953),
            .I(N__80907));
    LocalMux I__19095 (
            .O(N__80948),
            .I(N__80907));
    InMux I__19094 (
            .O(N__80945),
            .I(N__80904));
    InMux I__19093 (
            .O(N__80944),
            .I(N__80899));
    InMux I__19092 (
            .O(N__80943),
            .I(N__80899));
    InMux I__19091 (
            .O(N__80940),
            .I(N__80896));
    InMux I__19090 (
            .O(N__80939),
            .I(N__80893));
    InMux I__19089 (
            .O(N__80938),
            .I(N__80888));
    InMux I__19088 (
            .O(N__80935),
            .I(N__80888));
    Span4Mux_h I__19087 (
            .O(N__80932),
            .I(N__80885));
    CascadeMux I__19086 (
            .O(N__80931),
            .I(N__80882));
    LocalMux I__19085 (
            .O(N__80924),
            .I(N__80879));
    LocalMux I__19084 (
            .O(N__80919),
            .I(N__80876));
    LocalMux I__19083 (
            .O(N__80914),
            .I(N__80871));
    Span4Mux_v I__19082 (
            .O(N__80907),
            .I(N__80871));
    LocalMux I__19081 (
            .O(N__80904),
            .I(N__80868));
    LocalMux I__19080 (
            .O(N__80899),
            .I(N__80865));
    LocalMux I__19079 (
            .O(N__80896),
            .I(N__80858));
    LocalMux I__19078 (
            .O(N__80893),
            .I(N__80858));
    LocalMux I__19077 (
            .O(N__80888),
            .I(N__80858));
    Span4Mux_h I__19076 (
            .O(N__80885),
            .I(N__80854));
    InMux I__19075 (
            .O(N__80882),
            .I(N__80851));
    Span4Mux_v I__19074 (
            .O(N__80879),
            .I(N__80846));
    Span4Mux_h I__19073 (
            .O(N__80876),
            .I(N__80846));
    Span4Mux_h I__19072 (
            .O(N__80871),
            .I(N__80843));
    Span4Mux_v I__19071 (
            .O(N__80868),
            .I(N__80840));
    Span4Mux_h I__19070 (
            .O(N__80865),
            .I(N__80835));
    Span4Mux_v I__19069 (
            .O(N__80858),
            .I(N__80835));
    InMux I__19068 (
            .O(N__80857),
            .I(N__80832));
    Sp12to4 I__19067 (
            .O(N__80854),
            .I(N__80829));
    LocalMux I__19066 (
            .O(N__80851),
            .I(N__80826));
    Span4Mux_h I__19065 (
            .O(N__80846),
            .I(N__80823));
    Span4Mux_v I__19064 (
            .O(N__80843),
            .I(N__80820));
    Span4Mux_h I__19063 (
            .O(N__80840),
            .I(N__80817));
    Span4Mux_h I__19062 (
            .O(N__80835),
            .I(N__80814));
    LocalMux I__19061 (
            .O(N__80832),
            .I(N__80809));
    Span12Mux_s11_v I__19060 (
            .O(N__80829),
            .I(N__80809));
    Odrv12 I__19059 (
            .O(N__80826),
            .I(xy_ki_1_rep2));
    Odrv4 I__19058 (
            .O(N__80823),
            .I(xy_ki_1_rep2));
    Odrv4 I__19057 (
            .O(N__80820),
            .I(xy_ki_1_rep2));
    Odrv4 I__19056 (
            .O(N__80817),
            .I(xy_ki_1_rep2));
    Odrv4 I__19055 (
            .O(N__80814),
            .I(xy_ki_1_rep2));
    Odrv12 I__19054 (
            .O(N__80809),
            .I(xy_ki_1_rep2));
    CascadeMux I__19053 (
            .O(N__80796),
            .I(N__80788));
    InMux I__19052 (
            .O(N__80795),
            .I(N__80781));
    InMux I__19051 (
            .O(N__80794),
            .I(N__80781));
    InMux I__19050 (
            .O(N__80793),
            .I(N__80775));
    InMux I__19049 (
            .O(N__80792),
            .I(N__80771));
    InMux I__19048 (
            .O(N__80791),
            .I(N__80768));
    InMux I__19047 (
            .O(N__80788),
            .I(N__80759));
    InMux I__19046 (
            .O(N__80787),
            .I(N__80759));
    InMux I__19045 (
            .O(N__80786),
            .I(N__80756));
    LocalMux I__19044 (
            .O(N__80781),
            .I(N__80751));
    InMux I__19043 (
            .O(N__80780),
            .I(N__80748));
    InMux I__19042 (
            .O(N__80779),
            .I(N__80745));
    InMux I__19041 (
            .O(N__80778),
            .I(N__80742));
    LocalMux I__19040 (
            .O(N__80775),
            .I(N__80739));
    CascadeMux I__19039 (
            .O(N__80774),
            .I(N__80735));
    LocalMux I__19038 (
            .O(N__80771),
            .I(N__80732));
    LocalMux I__19037 (
            .O(N__80768),
            .I(N__80729));
    InMux I__19036 (
            .O(N__80767),
            .I(N__80726));
    CascadeMux I__19035 (
            .O(N__80766),
            .I(N__80722));
    InMux I__19034 (
            .O(N__80765),
            .I(N__80718));
    InMux I__19033 (
            .O(N__80764),
            .I(N__80715));
    LocalMux I__19032 (
            .O(N__80759),
            .I(N__80710));
    LocalMux I__19031 (
            .O(N__80756),
            .I(N__80710));
    InMux I__19030 (
            .O(N__80755),
            .I(N__80705));
    InMux I__19029 (
            .O(N__80754),
            .I(N__80705));
    Span4Mux_h I__19028 (
            .O(N__80751),
            .I(N__80699));
    LocalMux I__19027 (
            .O(N__80748),
            .I(N__80694));
    LocalMux I__19026 (
            .O(N__80745),
            .I(N__80694));
    LocalMux I__19025 (
            .O(N__80742),
            .I(N__80689));
    Span4Mux_v I__19024 (
            .O(N__80739),
            .I(N__80689));
    InMux I__19023 (
            .O(N__80738),
            .I(N__80686));
    InMux I__19022 (
            .O(N__80735),
            .I(N__80683));
    Span4Mux_v I__19021 (
            .O(N__80732),
            .I(N__80680));
    Span4Mux_v I__19020 (
            .O(N__80729),
            .I(N__80675));
    LocalMux I__19019 (
            .O(N__80726),
            .I(N__80675));
    InMux I__19018 (
            .O(N__80725),
            .I(N__80670));
    InMux I__19017 (
            .O(N__80722),
            .I(N__80670));
    InMux I__19016 (
            .O(N__80721),
            .I(N__80667));
    LocalMux I__19015 (
            .O(N__80718),
            .I(N__80664));
    LocalMux I__19014 (
            .O(N__80715),
            .I(N__80659));
    Span4Mux_v I__19013 (
            .O(N__80710),
            .I(N__80659));
    LocalMux I__19012 (
            .O(N__80705),
            .I(N__80656));
    InMux I__19011 (
            .O(N__80704),
            .I(N__80649));
    InMux I__19010 (
            .O(N__80703),
            .I(N__80649));
    InMux I__19009 (
            .O(N__80702),
            .I(N__80649));
    Span4Mux_v I__19008 (
            .O(N__80699),
            .I(N__80646));
    Span4Mux_h I__19007 (
            .O(N__80694),
            .I(N__80639));
    Span4Mux_v I__19006 (
            .O(N__80689),
            .I(N__80639));
    LocalMux I__19005 (
            .O(N__80686),
            .I(N__80639));
    LocalMux I__19004 (
            .O(N__80683),
            .I(xy_ki_0));
    Odrv4 I__19003 (
            .O(N__80680),
            .I(xy_ki_0));
    Odrv4 I__19002 (
            .O(N__80675),
            .I(xy_ki_0));
    LocalMux I__19001 (
            .O(N__80670),
            .I(xy_ki_0));
    LocalMux I__19000 (
            .O(N__80667),
            .I(xy_ki_0));
    Odrv12 I__18999 (
            .O(N__80664),
            .I(xy_ki_0));
    Odrv4 I__18998 (
            .O(N__80659),
            .I(xy_ki_0));
    Odrv4 I__18997 (
            .O(N__80656),
            .I(xy_ki_0));
    LocalMux I__18996 (
            .O(N__80649),
            .I(xy_ki_0));
    Odrv4 I__18995 (
            .O(N__80646),
            .I(xy_ki_0));
    Odrv4 I__18994 (
            .O(N__80639),
            .I(xy_ki_0));
    CascadeMux I__18993 (
            .O(N__80616),
            .I(N__80604));
    InMux I__18992 (
            .O(N__80615),
            .I(N__80600));
    InMux I__18991 (
            .O(N__80614),
            .I(N__80596));
    InMux I__18990 (
            .O(N__80613),
            .I(N__80591));
    InMux I__18989 (
            .O(N__80612),
            .I(N__80586));
    InMux I__18988 (
            .O(N__80611),
            .I(N__80586));
    InMux I__18987 (
            .O(N__80610),
            .I(N__80583));
    InMux I__18986 (
            .O(N__80609),
            .I(N__80580));
    InMux I__18985 (
            .O(N__80608),
            .I(N__80577));
    InMux I__18984 (
            .O(N__80607),
            .I(N__80572));
    InMux I__18983 (
            .O(N__80604),
            .I(N__80572));
    InMux I__18982 (
            .O(N__80603),
            .I(N__80569));
    LocalMux I__18981 (
            .O(N__80600),
            .I(N__80564));
    InMux I__18980 (
            .O(N__80599),
            .I(N__80561));
    LocalMux I__18979 (
            .O(N__80596),
            .I(N__80558));
    CascadeMux I__18978 (
            .O(N__80595),
            .I(N__80555));
    InMux I__18977 (
            .O(N__80594),
            .I(N__80551));
    LocalMux I__18976 (
            .O(N__80591),
            .I(N__80542));
    LocalMux I__18975 (
            .O(N__80586),
            .I(N__80542));
    LocalMux I__18974 (
            .O(N__80583),
            .I(N__80542));
    LocalMux I__18973 (
            .O(N__80580),
            .I(N__80542));
    LocalMux I__18972 (
            .O(N__80577),
            .I(N__80539));
    LocalMux I__18971 (
            .O(N__80572),
            .I(N__80529));
    LocalMux I__18970 (
            .O(N__80569),
            .I(N__80526));
    InMux I__18969 (
            .O(N__80568),
            .I(N__80523));
    CascadeMux I__18968 (
            .O(N__80567),
            .I(N__80516));
    Span4Mux_h I__18967 (
            .O(N__80564),
            .I(N__80512));
    LocalMux I__18966 (
            .O(N__80561),
            .I(N__80507));
    Span4Mux_v I__18965 (
            .O(N__80558),
            .I(N__80507));
    InMux I__18964 (
            .O(N__80555),
            .I(N__80502));
    InMux I__18963 (
            .O(N__80554),
            .I(N__80502));
    LocalMux I__18962 (
            .O(N__80551),
            .I(N__80497));
    Span4Mux_v I__18961 (
            .O(N__80542),
            .I(N__80497));
    Span4Mux_v I__18960 (
            .O(N__80539),
            .I(N__80494));
    InMux I__18959 (
            .O(N__80538),
            .I(N__80491));
    InMux I__18958 (
            .O(N__80537),
            .I(N__80484));
    InMux I__18957 (
            .O(N__80536),
            .I(N__80484));
    InMux I__18956 (
            .O(N__80535),
            .I(N__80484));
    InMux I__18955 (
            .O(N__80534),
            .I(N__80479));
    InMux I__18954 (
            .O(N__80533),
            .I(N__80479));
    InMux I__18953 (
            .O(N__80532),
            .I(N__80476));
    Span4Mux_h I__18952 (
            .O(N__80529),
            .I(N__80472));
    Span12Mux_s11_h I__18951 (
            .O(N__80526),
            .I(N__80467));
    LocalMux I__18950 (
            .O(N__80523),
            .I(N__80467));
    InMux I__18949 (
            .O(N__80522),
            .I(N__80460));
    InMux I__18948 (
            .O(N__80521),
            .I(N__80460));
    InMux I__18947 (
            .O(N__80520),
            .I(N__80460));
    InMux I__18946 (
            .O(N__80519),
            .I(N__80453));
    InMux I__18945 (
            .O(N__80516),
            .I(N__80453));
    InMux I__18944 (
            .O(N__80515),
            .I(N__80453));
    Sp12to4 I__18943 (
            .O(N__80512),
            .I(N__80450));
    Span4Mux_v I__18942 (
            .O(N__80507),
            .I(N__80441));
    LocalMux I__18941 (
            .O(N__80502),
            .I(N__80441));
    Span4Mux_v I__18940 (
            .O(N__80497),
            .I(N__80441));
    Span4Mux_h I__18939 (
            .O(N__80494),
            .I(N__80441));
    LocalMux I__18938 (
            .O(N__80491),
            .I(N__80436));
    LocalMux I__18937 (
            .O(N__80484),
            .I(N__80436));
    LocalMux I__18936 (
            .O(N__80479),
            .I(N__80431));
    LocalMux I__18935 (
            .O(N__80476),
            .I(N__80431));
    InMux I__18934 (
            .O(N__80475),
            .I(N__80428));
    Sp12to4 I__18933 (
            .O(N__80472),
            .I(N__80423));
    Span12Mux_s7_v I__18932 (
            .O(N__80467),
            .I(N__80423));
    LocalMux I__18931 (
            .O(N__80460),
            .I(N__80418));
    LocalMux I__18930 (
            .O(N__80453),
            .I(N__80418));
    Span12Mux_v I__18929 (
            .O(N__80450),
            .I(N__80413));
    Sp12to4 I__18928 (
            .O(N__80441),
            .I(N__80413));
    Span4Mux_v I__18927 (
            .O(N__80436),
            .I(N__80408));
    Span4Mux_h I__18926 (
            .O(N__80431),
            .I(N__80408));
    LocalMux I__18925 (
            .O(N__80428),
            .I(xy_ki_2_rep2));
    Odrv12 I__18924 (
            .O(N__80423),
            .I(xy_ki_2_rep2));
    Odrv4 I__18923 (
            .O(N__80418),
            .I(xy_ki_2_rep2));
    Odrv12 I__18922 (
            .O(N__80413),
            .I(xy_ki_2_rep2));
    Odrv4 I__18921 (
            .O(N__80408),
            .I(xy_ki_2_rep2));
    CascadeMux I__18920 (
            .O(N__80397),
            .I(N__80391));
    CascadeMux I__18919 (
            .O(N__80396),
            .I(N__80387));
    CascadeMux I__18918 (
            .O(N__80395),
            .I(N__80384));
    InMux I__18917 (
            .O(N__80394),
            .I(N__80379));
    InMux I__18916 (
            .O(N__80391),
            .I(N__80372));
    InMux I__18915 (
            .O(N__80390),
            .I(N__80372));
    InMux I__18914 (
            .O(N__80387),
            .I(N__80369));
    InMux I__18913 (
            .O(N__80384),
            .I(N__80366));
    CascadeMux I__18912 (
            .O(N__80383),
            .I(N__80360));
    InMux I__18911 (
            .O(N__80382),
            .I(N__80357));
    LocalMux I__18910 (
            .O(N__80379),
            .I(N__80354));
    InMux I__18909 (
            .O(N__80378),
            .I(N__80351));
    InMux I__18908 (
            .O(N__80377),
            .I(N__80348));
    LocalMux I__18907 (
            .O(N__80372),
            .I(N__80344));
    LocalMux I__18906 (
            .O(N__80369),
            .I(N__80341));
    LocalMux I__18905 (
            .O(N__80366),
            .I(N__80335));
    InMux I__18904 (
            .O(N__80365),
            .I(N__80330));
    InMux I__18903 (
            .O(N__80364),
            .I(N__80330));
    InMux I__18902 (
            .O(N__80363),
            .I(N__80327));
    InMux I__18901 (
            .O(N__80360),
            .I(N__80324));
    LocalMux I__18900 (
            .O(N__80357),
            .I(N__80321));
    Span4Mux_v I__18899 (
            .O(N__80354),
            .I(N__80318));
    LocalMux I__18898 (
            .O(N__80351),
            .I(N__80313));
    LocalMux I__18897 (
            .O(N__80348),
            .I(N__80313));
    InMux I__18896 (
            .O(N__80347),
            .I(N__80310));
    Span4Mux_v I__18895 (
            .O(N__80344),
            .I(N__80305));
    Span4Mux_v I__18894 (
            .O(N__80341),
            .I(N__80305));
    CascadeMux I__18893 (
            .O(N__80340),
            .I(N__80301));
    InMux I__18892 (
            .O(N__80339),
            .I(N__80298));
    InMux I__18891 (
            .O(N__80338),
            .I(N__80295));
    Span4Mux_v I__18890 (
            .O(N__80335),
            .I(N__80288));
    LocalMux I__18889 (
            .O(N__80330),
            .I(N__80288));
    LocalMux I__18888 (
            .O(N__80327),
            .I(N__80288));
    LocalMux I__18887 (
            .O(N__80324),
            .I(N__80284));
    Span4Mux_h I__18886 (
            .O(N__80321),
            .I(N__80281));
    Span4Mux_v I__18885 (
            .O(N__80318),
            .I(N__80278));
    Span4Mux_h I__18884 (
            .O(N__80313),
            .I(N__80275));
    LocalMux I__18883 (
            .O(N__80310),
            .I(N__80270));
    Span4Mux_v I__18882 (
            .O(N__80305),
            .I(N__80270));
    InMux I__18881 (
            .O(N__80304),
            .I(N__80267));
    InMux I__18880 (
            .O(N__80301),
            .I(N__80264));
    LocalMux I__18879 (
            .O(N__80298),
            .I(N__80261));
    LocalMux I__18878 (
            .O(N__80295),
            .I(N__80256));
    Span4Mux_v I__18877 (
            .O(N__80288),
            .I(N__80256));
    InMux I__18876 (
            .O(N__80287),
            .I(N__80253));
    Span12Mux_v I__18875 (
            .O(N__80284),
            .I(N__80250));
    Span4Mux_h I__18874 (
            .O(N__80281),
            .I(N__80239));
    Span4Mux_h I__18873 (
            .O(N__80278),
            .I(N__80239));
    Span4Mux_h I__18872 (
            .O(N__80275),
            .I(N__80239));
    Span4Mux_h I__18871 (
            .O(N__80270),
            .I(N__80239));
    LocalMux I__18870 (
            .O(N__80267),
            .I(N__80239));
    LocalMux I__18869 (
            .O(N__80264),
            .I(N__80230));
    Span4Mux_v I__18868 (
            .O(N__80261),
            .I(N__80230));
    Span4Mux_v I__18867 (
            .O(N__80256),
            .I(N__80230));
    LocalMux I__18866 (
            .O(N__80253),
            .I(N__80230));
    Odrv12 I__18865 (
            .O(N__80250),
            .I(xy_ki_3_rep1));
    Odrv4 I__18864 (
            .O(N__80239),
            .I(xy_ki_3_rep1));
    Odrv4 I__18863 (
            .O(N__80230),
            .I(xy_ki_3_rep1));
    InMux I__18862 (
            .O(N__80223),
            .I(N__80217));
    InMux I__18861 (
            .O(N__80222),
            .I(N__80217));
    LocalMux I__18860 (
            .O(N__80217),
            .I(N__80214));
    Span4Mux_h I__18859 (
            .O(N__80214),
            .I(N__80210));
    InMux I__18858 (
            .O(N__80213),
            .I(N__80207));
    Span4Mux_v I__18857 (
            .O(N__80210),
            .I(N__80202));
    LocalMux I__18856 (
            .O(N__80207),
            .I(N__80202));
    Span4Mux_h I__18855 (
            .O(N__80202),
            .I(N__80198));
    InMux I__18854 (
            .O(N__80201),
            .I(N__80195));
    Odrv4 I__18853 (
            .O(N__80198),
            .I(\pid_side.m0_0_03 ));
    LocalMux I__18852 (
            .O(N__80195),
            .I(\pid_side.m0_0_03 ));
    InMux I__18851 (
            .O(N__80190),
            .I(N__80187));
    LocalMux I__18850 (
            .O(N__80187),
            .I(N__80184));
    Span4Mux_v I__18849 (
            .O(N__80184),
            .I(N__80181));
    Odrv4 I__18848 (
            .O(N__80181),
            .I(\pid_side.m0_2_03 ));
    InMux I__18847 (
            .O(N__80178),
            .I(N__80175));
    LocalMux I__18846 (
            .O(N__80175),
            .I(N__80172));
    Odrv12 I__18845 (
            .O(N__80172),
            .I(\pid_side.O_2_7 ));
    InMux I__18844 (
            .O(N__80169),
            .I(N__80166));
    LocalMux I__18843 (
            .O(N__80166),
            .I(N__80163));
    Span4Mux_h I__18842 (
            .O(N__80163),
            .I(N__80160));
    Odrv4 I__18841 (
            .O(N__80160),
            .I(\pid_side.O_2_12 ));
    InMux I__18840 (
            .O(N__80157),
            .I(N__80151));
    InMux I__18839 (
            .O(N__80156),
            .I(N__80151));
    LocalMux I__18838 (
            .O(N__80151),
            .I(N__80148));
    Span4Mux_h I__18837 (
            .O(N__80148),
            .I(N__80145));
    Span4Mux_h I__18836 (
            .O(N__80145),
            .I(N__80142));
    Odrv4 I__18835 (
            .O(N__80142),
            .I(\pid_side.error_p_regZ0Z_9 ));
    InMux I__18834 (
            .O(N__80139),
            .I(N__80136));
    LocalMux I__18833 (
            .O(N__80136),
            .I(N__80133));
    Span12Mux_s10_v I__18832 (
            .O(N__80133),
            .I(N__80130));
    Odrv12 I__18831 (
            .O(N__80130),
            .I(\pid_side.O_2_8 ));
    CascadeMux I__18830 (
            .O(N__80127),
            .I(N__80123));
    InMux I__18829 (
            .O(N__80126),
            .I(N__80118));
    InMux I__18828 (
            .O(N__80123),
            .I(N__80118));
    LocalMux I__18827 (
            .O(N__80118),
            .I(\pid_side.error_p_regZ0Z_5 ));
    InMux I__18826 (
            .O(N__80115),
            .I(N__80112));
    LocalMux I__18825 (
            .O(N__80112),
            .I(N__80108));
    CascadeMux I__18824 (
            .O(N__80111),
            .I(N__80105));
    Span4Mux_v I__18823 (
            .O(N__80108),
            .I(N__80101));
    InMux I__18822 (
            .O(N__80105),
            .I(N__80096));
    InMux I__18821 (
            .O(N__80104),
            .I(N__80096));
    Odrv4 I__18820 (
            .O(N__80101),
            .I(\pid_side.error_d_reg_prev_esr_RNI73UC2_0Z0Z_14 ));
    LocalMux I__18819 (
            .O(N__80096),
            .I(\pid_side.error_d_reg_prev_esr_RNI73UC2_0Z0Z_14 ));
    InMux I__18818 (
            .O(N__80091),
            .I(N__80088));
    LocalMux I__18817 (
            .O(N__80088),
            .I(N__80085));
    Span4Mux_h I__18816 (
            .O(N__80085),
            .I(N__80082));
    Odrv4 I__18815 (
            .O(N__80082),
            .I(\pid_side.error_d_reg_prev_esr_RNI0UI8JZ0Z_12 ));
    InMux I__18814 (
            .O(N__80079),
            .I(N__80076));
    LocalMux I__18813 (
            .O(N__80076),
            .I(N__80073));
    Odrv12 I__18812 (
            .O(N__80073),
            .I(\pid_side.error_d_reg_prev_esr_RNI5RIO_0Z0Z_14 ));
    CascadeMux I__18811 (
            .O(N__80070),
            .I(\pid_side.un1_pid_prereg_97_cascade_ ));
    CascadeMux I__18810 (
            .O(N__80067),
            .I(N__80064));
    InMux I__18809 (
            .O(N__80064),
            .I(N__80061));
    LocalMux I__18808 (
            .O(N__80061),
            .I(N__80058));
    Span4Mux_v I__18807 (
            .O(N__80058),
            .I(N__80053));
    InMux I__18806 (
            .O(N__80057),
            .I(N__80048));
    InMux I__18805 (
            .O(N__80056),
            .I(N__80048));
    Odrv4 I__18804 (
            .O(N__80053),
            .I(\pid_side.error_d_reg_prev_esr_RNI45PU7Z0Z_12 ));
    LocalMux I__18803 (
            .O(N__80048),
            .I(\pid_side.error_d_reg_prev_esr_RNI45PU7Z0Z_12 ));
    InMux I__18802 (
            .O(N__80043),
            .I(N__80040));
    LocalMux I__18801 (
            .O(N__80040),
            .I(\pid_side.error_d_reg_fast_esr_RNIPHKNZ0Z_12 ));
    InMux I__18800 (
            .O(N__80037),
            .I(N__80034));
    LocalMux I__18799 (
            .O(N__80034),
            .I(\pid_side.error_d_reg_fast_esr_RNIPEC11Z0Z_12 ));
    CascadeMux I__18798 (
            .O(N__80031),
            .I(\pid_side.error_d_reg_fast_esr_RNIEIJH2Z0Z_12_cascade_ ));
    CascadeMux I__18797 (
            .O(N__80028),
            .I(\pid_side.g1_2_1_cascade_ ));
    CascadeMux I__18796 (
            .O(N__80025),
            .I(\pid_side.g1_3_cascade_ ));
    CascadeMux I__18795 (
            .O(N__80022),
            .I(N__80019));
    InMux I__18794 (
            .O(N__80019),
            .I(N__80016));
    LocalMux I__18793 (
            .O(N__80016),
            .I(N__80012));
    InMux I__18792 (
            .O(N__80015),
            .I(N__80009));
    Span4Mux_h I__18791 (
            .O(N__80012),
            .I(N__80006));
    LocalMux I__18790 (
            .O(N__80009),
            .I(\pid_side.error_p_reg_esr_RNILLRS8Z0Z_12 ));
    Odrv4 I__18789 (
            .O(N__80006),
            .I(\pid_side.error_p_reg_esr_RNILLRS8Z0Z_12 ));
    CascadeMux I__18788 (
            .O(N__80001),
            .I(N__79987));
    CascadeMux I__18787 (
            .O(N__80000),
            .I(N__79970));
    CascadeMux I__18786 (
            .O(N__79999),
            .I(N__79938));
    InMux I__18785 (
            .O(N__79998),
            .I(N__79912));
    InMux I__18784 (
            .O(N__79997),
            .I(N__79909));
    InMux I__18783 (
            .O(N__79996),
            .I(N__79904));
    InMux I__18782 (
            .O(N__79995),
            .I(N__79904));
    InMux I__18781 (
            .O(N__79994),
            .I(N__79901));
    InMux I__18780 (
            .O(N__79993),
            .I(N__79896));
    InMux I__18779 (
            .O(N__79992),
            .I(N__79896));
    InMux I__18778 (
            .O(N__79991),
            .I(N__79893));
    InMux I__18777 (
            .O(N__79990),
            .I(N__79888));
    InMux I__18776 (
            .O(N__79987),
            .I(N__79888));
    InMux I__18775 (
            .O(N__79986),
            .I(N__79885));
    InMux I__18774 (
            .O(N__79985),
            .I(N__79882));
    InMux I__18773 (
            .O(N__79984),
            .I(N__79879));
    InMux I__18772 (
            .O(N__79983),
            .I(N__79876));
    InMux I__18771 (
            .O(N__79982),
            .I(N__79871));
    InMux I__18770 (
            .O(N__79981),
            .I(N__79871));
    InMux I__18769 (
            .O(N__79980),
            .I(N__79864));
    InMux I__18768 (
            .O(N__79979),
            .I(N__79864));
    InMux I__18767 (
            .O(N__79978),
            .I(N__79864));
    InMux I__18766 (
            .O(N__79977),
            .I(N__79857));
    InMux I__18765 (
            .O(N__79976),
            .I(N__79857));
    InMux I__18764 (
            .O(N__79975),
            .I(N__79857));
    InMux I__18763 (
            .O(N__79974),
            .I(N__79850));
    InMux I__18762 (
            .O(N__79973),
            .I(N__79850));
    InMux I__18761 (
            .O(N__79970),
            .I(N__79850));
    InMux I__18760 (
            .O(N__79969),
            .I(N__79845));
    InMux I__18759 (
            .O(N__79968),
            .I(N__79845));
    InMux I__18758 (
            .O(N__79967),
            .I(N__79842));
    InMux I__18757 (
            .O(N__79966),
            .I(N__79839));
    InMux I__18756 (
            .O(N__79965),
            .I(N__79836));
    InMux I__18755 (
            .O(N__79964),
            .I(N__79831));
    InMux I__18754 (
            .O(N__79963),
            .I(N__79831));
    InMux I__18753 (
            .O(N__79962),
            .I(N__79826));
    InMux I__18752 (
            .O(N__79961),
            .I(N__79826));
    InMux I__18751 (
            .O(N__79960),
            .I(N__79823));
    InMux I__18750 (
            .O(N__79959),
            .I(N__79820));
    InMux I__18749 (
            .O(N__79958),
            .I(N__79813));
    InMux I__18748 (
            .O(N__79957),
            .I(N__79813));
    InMux I__18747 (
            .O(N__79956),
            .I(N__79813));
    InMux I__18746 (
            .O(N__79955),
            .I(N__79810));
    InMux I__18745 (
            .O(N__79954),
            .I(N__79805));
    InMux I__18744 (
            .O(N__79953),
            .I(N__79805));
    InMux I__18743 (
            .O(N__79952),
            .I(N__79800));
    InMux I__18742 (
            .O(N__79951),
            .I(N__79800));
    InMux I__18741 (
            .O(N__79950),
            .I(N__79793));
    InMux I__18740 (
            .O(N__79949),
            .I(N__79793));
    InMux I__18739 (
            .O(N__79948),
            .I(N__79793));
    InMux I__18738 (
            .O(N__79947),
            .I(N__79784));
    InMux I__18737 (
            .O(N__79946),
            .I(N__79784));
    InMux I__18736 (
            .O(N__79945),
            .I(N__79784));
    InMux I__18735 (
            .O(N__79944),
            .I(N__79784));
    InMux I__18734 (
            .O(N__79943),
            .I(N__79779));
    InMux I__18733 (
            .O(N__79942),
            .I(N__79779));
    InMux I__18732 (
            .O(N__79941),
            .I(N__79776));
    InMux I__18731 (
            .O(N__79938),
            .I(N__79771));
    InMux I__18730 (
            .O(N__79937),
            .I(N__79771));
    InMux I__18729 (
            .O(N__79936),
            .I(N__79768));
    InMux I__18728 (
            .O(N__79935),
            .I(N__79765));
    InMux I__18727 (
            .O(N__79934),
            .I(N__79762));
    InMux I__18726 (
            .O(N__79933),
            .I(N__79759));
    InMux I__18725 (
            .O(N__79932),
            .I(N__79752));
    InMux I__18724 (
            .O(N__79931),
            .I(N__79752));
    InMux I__18723 (
            .O(N__79930),
            .I(N__79752));
    InMux I__18722 (
            .O(N__79929),
            .I(N__79747));
    InMux I__18721 (
            .O(N__79928),
            .I(N__79747));
    InMux I__18720 (
            .O(N__79927),
            .I(N__79740));
    InMux I__18719 (
            .O(N__79926),
            .I(N__79740));
    InMux I__18718 (
            .O(N__79925),
            .I(N__79740));
    InMux I__18717 (
            .O(N__79924),
            .I(N__79737));
    InMux I__18716 (
            .O(N__79923),
            .I(N__79732));
    InMux I__18715 (
            .O(N__79922),
            .I(N__79732));
    InMux I__18714 (
            .O(N__79921),
            .I(N__79725));
    InMux I__18713 (
            .O(N__79920),
            .I(N__79725));
    InMux I__18712 (
            .O(N__79919),
            .I(N__79725));
    InMux I__18711 (
            .O(N__79918),
            .I(N__79722));
    InMux I__18710 (
            .O(N__79917),
            .I(N__79719));
    InMux I__18709 (
            .O(N__79916),
            .I(N__79716));
    InMux I__18708 (
            .O(N__79915),
            .I(N__79713));
    LocalMux I__18707 (
            .O(N__79912),
            .I(N__79553));
    LocalMux I__18706 (
            .O(N__79909),
            .I(N__79550));
    LocalMux I__18705 (
            .O(N__79904),
            .I(N__79547));
    LocalMux I__18704 (
            .O(N__79901),
            .I(N__79544));
    LocalMux I__18703 (
            .O(N__79896),
            .I(N__79541));
    LocalMux I__18702 (
            .O(N__79893),
            .I(N__79538));
    LocalMux I__18701 (
            .O(N__79888),
            .I(N__79535));
    LocalMux I__18700 (
            .O(N__79885),
            .I(N__79532));
    LocalMux I__18699 (
            .O(N__79882),
            .I(N__79529));
    LocalMux I__18698 (
            .O(N__79879),
            .I(N__79526));
    LocalMux I__18697 (
            .O(N__79876),
            .I(N__79523));
    LocalMux I__18696 (
            .O(N__79871),
            .I(N__79520));
    LocalMux I__18695 (
            .O(N__79864),
            .I(N__79517));
    LocalMux I__18694 (
            .O(N__79857),
            .I(N__79514));
    LocalMux I__18693 (
            .O(N__79850),
            .I(N__79511));
    LocalMux I__18692 (
            .O(N__79845),
            .I(N__79508));
    LocalMux I__18691 (
            .O(N__79842),
            .I(N__79505));
    LocalMux I__18690 (
            .O(N__79839),
            .I(N__79502));
    LocalMux I__18689 (
            .O(N__79836),
            .I(N__79499));
    LocalMux I__18688 (
            .O(N__79831),
            .I(N__79496));
    LocalMux I__18687 (
            .O(N__79826),
            .I(N__79493));
    LocalMux I__18686 (
            .O(N__79823),
            .I(N__79490));
    LocalMux I__18685 (
            .O(N__79820),
            .I(N__79487));
    LocalMux I__18684 (
            .O(N__79813),
            .I(N__79484));
    LocalMux I__18683 (
            .O(N__79810),
            .I(N__79481));
    LocalMux I__18682 (
            .O(N__79805),
            .I(N__79478));
    LocalMux I__18681 (
            .O(N__79800),
            .I(N__79475));
    LocalMux I__18680 (
            .O(N__79793),
            .I(N__79472));
    LocalMux I__18679 (
            .O(N__79784),
            .I(N__79469));
    LocalMux I__18678 (
            .O(N__79779),
            .I(N__79466));
    LocalMux I__18677 (
            .O(N__79776),
            .I(N__79463));
    LocalMux I__18676 (
            .O(N__79771),
            .I(N__79460));
    LocalMux I__18675 (
            .O(N__79768),
            .I(N__79457));
    LocalMux I__18674 (
            .O(N__79765),
            .I(N__79454));
    LocalMux I__18673 (
            .O(N__79762),
            .I(N__79451));
    LocalMux I__18672 (
            .O(N__79759),
            .I(N__79448));
    LocalMux I__18671 (
            .O(N__79752),
            .I(N__79445));
    LocalMux I__18670 (
            .O(N__79747),
            .I(N__79442));
    LocalMux I__18669 (
            .O(N__79740),
            .I(N__79439));
    LocalMux I__18668 (
            .O(N__79737),
            .I(N__79436));
    LocalMux I__18667 (
            .O(N__79732),
            .I(N__79433));
    LocalMux I__18666 (
            .O(N__79725),
            .I(N__79430));
    LocalMux I__18665 (
            .O(N__79722),
            .I(N__79427));
    LocalMux I__18664 (
            .O(N__79719),
            .I(N__79424));
    LocalMux I__18663 (
            .O(N__79716),
            .I(N__79421));
    LocalMux I__18662 (
            .O(N__79713),
            .I(N__79418));
    SRMux I__18661 (
            .O(N__79712),
            .I(N__79011));
    SRMux I__18660 (
            .O(N__79711),
            .I(N__79011));
    SRMux I__18659 (
            .O(N__79710),
            .I(N__79011));
    SRMux I__18658 (
            .O(N__79709),
            .I(N__79011));
    SRMux I__18657 (
            .O(N__79708),
            .I(N__79011));
    SRMux I__18656 (
            .O(N__79707),
            .I(N__79011));
    SRMux I__18655 (
            .O(N__79706),
            .I(N__79011));
    SRMux I__18654 (
            .O(N__79705),
            .I(N__79011));
    SRMux I__18653 (
            .O(N__79704),
            .I(N__79011));
    SRMux I__18652 (
            .O(N__79703),
            .I(N__79011));
    SRMux I__18651 (
            .O(N__79702),
            .I(N__79011));
    SRMux I__18650 (
            .O(N__79701),
            .I(N__79011));
    SRMux I__18649 (
            .O(N__79700),
            .I(N__79011));
    SRMux I__18648 (
            .O(N__79699),
            .I(N__79011));
    SRMux I__18647 (
            .O(N__79698),
            .I(N__79011));
    SRMux I__18646 (
            .O(N__79697),
            .I(N__79011));
    SRMux I__18645 (
            .O(N__79696),
            .I(N__79011));
    SRMux I__18644 (
            .O(N__79695),
            .I(N__79011));
    SRMux I__18643 (
            .O(N__79694),
            .I(N__79011));
    SRMux I__18642 (
            .O(N__79693),
            .I(N__79011));
    SRMux I__18641 (
            .O(N__79692),
            .I(N__79011));
    SRMux I__18640 (
            .O(N__79691),
            .I(N__79011));
    SRMux I__18639 (
            .O(N__79690),
            .I(N__79011));
    SRMux I__18638 (
            .O(N__79689),
            .I(N__79011));
    SRMux I__18637 (
            .O(N__79688),
            .I(N__79011));
    SRMux I__18636 (
            .O(N__79687),
            .I(N__79011));
    SRMux I__18635 (
            .O(N__79686),
            .I(N__79011));
    SRMux I__18634 (
            .O(N__79685),
            .I(N__79011));
    SRMux I__18633 (
            .O(N__79684),
            .I(N__79011));
    SRMux I__18632 (
            .O(N__79683),
            .I(N__79011));
    SRMux I__18631 (
            .O(N__79682),
            .I(N__79011));
    SRMux I__18630 (
            .O(N__79681),
            .I(N__79011));
    SRMux I__18629 (
            .O(N__79680),
            .I(N__79011));
    SRMux I__18628 (
            .O(N__79679),
            .I(N__79011));
    SRMux I__18627 (
            .O(N__79678),
            .I(N__79011));
    SRMux I__18626 (
            .O(N__79677),
            .I(N__79011));
    SRMux I__18625 (
            .O(N__79676),
            .I(N__79011));
    SRMux I__18624 (
            .O(N__79675),
            .I(N__79011));
    SRMux I__18623 (
            .O(N__79674),
            .I(N__79011));
    SRMux I__18622 (
            .O(N__79673),
            .I(N__79011));
    SRMux I__18621 (
            .O(N__79672),
            .I(N__79011));
    SRMux I__18620 (
            .O(N__79671),
            .I(N__79011));
    SRMux I__18619 (
            .O(N__79670),
            .I(N__79011));
    SRMux I__18618 (
            .O(N__79669),
            .I(N__79011));
    SRMux I__18617 (
            .O(N__79668),
            .I(N__79011));
    SRMux I__18616 (
            .O(N__79667),
            .I(N__79011));
    SRMux I__18615 (
            .O(N__79666),
            .I(N__79011));
    SRMux I__18614 (
            .O(N__79665),
            .I(N__79011));
    SRMux I__18613 (
            .O(N__79664),
            .I(N__79011));
    SRMux I__18612 (
            .O(N__79663),
            .I(N__79011));
    SRMux I__18611 (
            .O(N__79662),
            .I(N__79011));
    SRMux I__18610 (
            .O(N__79661),
            .I(N__79011));
    SRMux I__18609 (
            .O(N__79660),
            .I(N__79011));
    SRMux I__18608 (
            .O(N__79659),
            .I(N__79011));
    SRMux I__18607 (
            .O(N__79658),
            .I(N__79011));
    SRMux I__18606 (
            .O(N__79657),
            .I(N__79011));
    SRMux I__18605 (
            .O(N__79656),
            .I(N__79011));
    SRMux I__18604 (
            .O(N__79655),
            .I(N__79011));
    SRMux I__18603 (
            .O(N__79654),
            .I(N__79011));
    SRMux I__18602 (
            .O(N__79653),
            .I(N__79011));
    SRMux I__18601 (
            .O(N__79652),
            .I(N__79011));
    SRMux I__18600 (
            .O(N__79651),
            .I(N__79011));
    SRMux I__18599 (
            .O(N__79650),
            .I(N__79011));
    SRMux I__18598 (
            .O(N__79649),
            .I(N__79011));
    SRMux I__18597 (
            .O(N__79648),
            .I(N__79011));
    SRMux I__18596 (
            .O(N__79647),
            .I(N__79011));
    SRMux I__18595 (
            .O(N__79646),
            .I(N__79011));
    SRMux I__18594 (
            .O(N__79645),
            .I(N__79011));
    SRMux I__18593 (
            .O(N__79644),
            .I(N__79011));
    SRMux I__18592 (
            .O(N__79643),
            .I(N__79011));
    SRMux I__18591 (
            .O(N__79642),
            .I(N__79011));
    SRMux I__18590 (
            .O(N__79641),
            .I(N__79011));
    SRMux I__18589 (
            .O(N__79640),
            .I(N__79011));
    SRMux I__18588 (
            .O(N__79639),
            .I(N__79011));
    SRMux I__18587 (
            .O(N__79638),
            .I(N__79011));
    SRMux I__18586 (
            .O(N__79637),
            .I(N__79011));
    SRMux I__18585 (
            .O(N__79636),
            .I(N__79011));
    SRMux I__18584 (
            .O(N__79635),
            .I(N__79011));
    SRMux I__18583 (
            .O(N__79634),
            .I(N__79011));
    SRMux I__18582 (
            .O(N__79633),
            .I(N__79011));
    SRMux I__18581 (
            .O(N__79632),
            .I(N__79011));
    SRMux I__18580 (
            .O(N__79631),
            .I(N__79011));
    SRMux I__18579 (
            .O(N__79630),
            .I(N__79011));
    SRMux I__18578 (
            .O(N__79629),
            .I(N__79011));
    SRMux I__18577 (
            .O(N__79628),
            .I(N__79011));
    SRMux I__18576 (
            .O(N__79627),
            .I(N__79011));
    SRMux I__18575 (
            .O(N__79626),
            .I(N__79011));
    SRMux I__18574 (
            .O(N__79625),
            .I(N__79011));
    SRMux I__18573 (
            .O(N__79624),
            .I(N__79011));
    SRMux I__18572 (
            .O(N__79623),
            .I(N__79011));
    SRMux I__18571 (
            .O(N__79622),
            .I(N__79011));
    SRMux I__18570 (
            .O(N__79621),
            .I(N__79011));
    SRMux I__18569 (
            .O(N__79620),
            .I(N__79011));
    SRMux I__18568 (
            .O(N__79619),
            .I(N__79011));
    SRMux I__18567 (
            .O(N__79618),
            .I(N__79011));
    SRMux I__18566 (
            .O(N__79617),
            .I(N__79011));
    SRMux I__18565 (
            .O(N__79616),
            .I(N__79011));
    SRMux I__18564 (
            .O(N__79615),
            .I(N__79011));
    SRMux I__18563 (
            .O(N__79614),
            .I(N__79011));
    SRMux I__18562 (
            .O(N__79613),
            .I(N__79011));
    SRMux I__18561 (
            .O(N__79612),
            .I(N__79011));
    SRMux I__18560 (
            .O(N__79611),
            .I(N__79011));
    SRMux I__18559 (
            .O(N__79610),
            .I(N__79011));
    SRMux I__18558 (
            .O(N__79609),
            .I(N__79011));
    SRMux I__18557 (
            .O(N__79608),
            .I(N__79011));
    SRMux I__18556 (
            .O(N__79607),
            .I(N__79011));
    SRMux I__18555 (
            .O(N__79606),
            .I(N__79011));
    SRMux I__18554 (
            .O(N__79605),
            .I(N__79011));
    SRMux I__18553 (
            .O(N__79604),
            .I(N__79011));
    SRMux I__18552 (
            .O(N__79603),
            .I(N__79011));
    SRMux I__18551 (
            .O(N__79602),
            .I(N__79011));
    SRMux I__18550 (
            .O(N__79601),
            .I(N__79011));
    SRMux I__18549 (
            .O(N__79600),
            .I(N__79011));
    SRMux I__18548 (
            .O(N__79599),
            .I(N__79011));
    SRMux I__18547 (
            .O(N__79598),
            .I(N__79011));
    SRMux I__18546 (
            .O(N__79597),
            .I(N__79011));
    SRMux I__18545 (
            .O(N__79596),
            .I(N__79011));
    SRMux I__18544 (
            .O(N__79595),
            .I(N__79011));
    SRMux I__18543 (
            .O(N__79594),
            .I(N__79011));
    SRMux I__18542 (
            .O(N__79593),
            .I(N__79011));
    SRMux I__18541 (
            .O(N__79592),
            .I(N__79011));
    SRMux I__18540 (
            .O(N__79591),
            .I(N__79011));
    SRMux I__18539 (
            .O(N__79590),
            .I(N__79011));
    SRMux I__18538 (
            .O(N__79589),
            .I(N__79011));
    SRMux I__18537 (
            .O(N__79588),
            .I(N__79011));
    SRMux I__18536 (
            .O(N__79587),
            .I(N__79011));
    SRMux I__18535 (
            .O(N__79586),
            .I(N__79011));
    SRMux I__18534 (
            .O(N__79585),
            .I(N__79011));
    SRMux I__18533 (
            .O(N__79584),
            .I(N__79011));
    SRMux I__18532 (
            .O(N__79583),
            .I(N__79011));
    SRMux I__18531 (
            .O(N__79582),
            .I(N__79011));
    SRMux I__18530 (
            .O(N__79581),
            .I(N__79011));
    SRMux I__18529 (
            .O(N__79580),
            .I(N__79011));
    SRMux I__18528 (
            .O(N__79579),
            .I(N__79011));
    SRMux I__18527 (
            .O(N__79578),
            .I(N__79011));
    SRMux I__18526 (
            .O(N__79577),
            .I(N__79011));
    SRMux I__18525 (
            .O(N__79576),
            .I(N__79011));
    SRMux I__18524 (
            .O(N__79575),
            .I(N__79011));
    SRMux I__18523 (
            .O(N__79574),
            .I(N__79011));
    SRMux I__18522 (
            .O(N__79573),
            .I(N__79011));
    SRMux I__18521 (
            .O(N__79572),
            .I(N__79011));
    SRMux I__18520 (
            .O(N__79571),
            .I(N__79011));
    SRMux I__18519 (
            .O(N__79570),
            .I(N__79011));
    SRMux I__18518 (
            .O(N__79569),
            .I(N__79011));
    SRMux I__18517 (
            .O(N__79568),
            .I(N__79011));
    SRMux I__18516 (
            .O(N__79567),
            .I(N__79011));
    SRMux I__18515 (
            .O(N__79566),
            .I(N__79011));
    SRMux I__18514 (
            .O(N__79565),
            .I(N__79011));
    SRMux I__18513 (
            .O(N__79564),
            .I(N__79011));
    SRMux I__18512 (
            .O(N__79563),
            .I(N__79011));
    SRMux I__18511 (
            .O(N__79562),
            .I(N__79011));
    SRMux I__18510 (
            .O(N__79561),
            .I(N__79011));
    SRMux I__18509 (
            .O(N__79560),
            .I(N__79011));
    SRMux I__18508 (
            .O(N__79559),
            .I(N__79011));
    SRMux I__18507 (
            .O(N__79558),
            .I(N__79011));
    SRMux I__18506 (
            .O(N__79557),
            .I(N__79011));
    SRMux I__18505 (
            .O(N__79556),
            .I(N__79011));
    Glb2LocalMux I__18504 (
            .O(N__79553),
            .I(N__79011));
    Glb2LocalMux I__18503 (
            .O(N__79550),
            .I(N__79011));
    Glb2LocalMux I__18502 (
            .O(N__79547),
            .I(N__79011));
    Glb2LocalMux I__18501 (
            .O(N__79544),
            .I(N__79011));
    Glb2LocalMux I__18500 (
            .O(N__79541),
            .I(N__79011));
    Glb2LocalMux I__18499 (
            .O(N__79538),
            .I(N__79011));
    Glb2LocalMux I__18498 (
            .O(N__79535),
            .I(N__79011));
    Glb2LocalMux I__18497 (
            .O(N__79532),
            .I(N__79011));
    Glb2LocalMux I__18496 (
            .O(N__79529),
            .I(N__79011));
    Glb2LocalMux I__18495 (
            .O(N__79526),
            .I(N__79011));
    Glb2LocalMux I__18494 (
            .O(N__79523),
            .I(N__79011));
    Glb2LocalMux I__18493 (
            .O(N__79520),
            .I(N__79011));
    Glb2LocalMux I__18492 (
            .O(N__79517),
            .I(N__79011));
    Glb2LocalMux I__18491 (
            .O(N__79514),
            .I(N__79011));
    Glb2LocalMux I__18490 (
            .O(N__79511),
            .I(N__79011));
    Glb2LocalMux I__18489 (
            .O(N__79508),
            .I(N__79011));
    Glb2LocalMux I__18488 (
            .O(N__79505),
            .I(N__79011));
    Glb2LocalMux I__18487 (
            .O(N__79502),
            .I(N__79011));
    Glb2LocalMux I__18486 (
            .O(N__79499),
            .I(N__79011));
    Glb2LocalMux I__18485 (
            .O(N__79496),
            .I(N__79011));
    Glb2LocalMux I__18484 (
            .O(N__79493),
            .I(N__79011));
    Glb2LocalMux I__18483 (
            .O(N__79490),
            .I(N__79011));
    Glb2LocalMux I__18482 (
            .O(N__79487),
            .I(N__79011));
    Glb2LocalMux I__18481 (
            .O(N__79484),
            .I(N__79011));
    Glb2LocalMux I__18480 (
            .O(N__79481),
            .I(N__79011));
    Glb2LocalMux I__18479 (
            .O(N__79478),
            .I(N__79011));
    Glb2LocalMux I__18478 (
            .O(N__79475),
            .I(N__79011));
    Glb2LocalMux I__18477 (
            .O(N__79472),
            .I(N__79011));
    Glb2LocalMux I__18476 (
            .O(N__79469),
            .I(N__79011));
    Glb2LocalMux I__18475 (
            .O(N__79466),
            .I(N__79011));
    Glb2LocalMux I__18474 (
            .O(N__79463),
            .I(N__79011));
    Glb2LocalMux I__18473 (
            .O(N__79460),
            .I(N__79011));
    Glb2LocalMux I__18472 (
            .O(N__79457),
            .I(N__79011));
    Glb2LocalMux I__18471 (
            .O(N__79454),
            .I(N__79011));
    Glb2LocalMux I__18470 (
            .O(N__79451),
            .I(N__79011));
    Glb2LocalMux I__18469 (
            .O(N__79448),
            .I(N__79011));
    Glb2LocalMux I__18468 (
            .O(N__79445),
            .I(N__79011));
    Glb2LocalMux I__18467 (
            .O(N__79442),
            .I(N__79011));
    Glb2LocalMux I__18466 (
            .O(N__79439),
            .I(N__79011));
    Glb2LocalMux I__18465 (
            .O(N__79436),
            .I(N__79011));
    Glb2LocalMux I__18464 (
            .O(N__79433),
            .I(N__79011));
    Glb2LocalMux I__18463 (
            .O(N__79430),
            .I(N__79011));
    Glb2LocalMux I__18462 (
            .O(N__79427),
            .I(N__79011));
    Glb2LocalMux I__18461 (
            .O(N__79424),
            .I(N__79011));
    Glb2LocalMux I__18460 (
            .O(N__79421),
            .I(N__79011));
    Glb2LocalMux I__18459 (
            .O(N__79418),
            .I(N__79011));
    GlobalMux I__18458 (
            .O(N__79011),
            .I(N__79008));
    gio2CtrlBuf I__18457 (
            .O(N__79008),
            .I(reset_system_g));
    InMux I__18456 (
            .O(N__79005),
            .I(N__79002));
    LocalMux I__18455 (
            .O(N__79002),
            .I(N__78999));
    Span4Mux_h I__18454 (
            .O(N__78999),
            .I(N__78996));
    Odrv4 I__18453 (
            .O(N__78996),
            .I(\pid_side.error_d_reg_prev_esr_RNI5RIOZ0Z_14 ));
    CascadeMux I__18452 (
            .O(N__78993),
            .I(\pid_side.error_d_reg_prev_esr_RNI5RIOZ0Z_14_cascade_ ));
    InMux I__18451 (
            .O(N__78990),
            .I(N__78986));
    InMux I__18450 (
            .O(N__78989),
            .I(N__78983));
    LocalMux I__18449 (
            .O(N__78986),
            .I(N__78979));
    LocalMux I__18448 (
            .O(N__78983),
            .I(N__78976));
    InMux I__18447 (
            .O(N__78982),
            .I(N__78973));
    Span4Mux_v I__18446 (
            .O(N__78979),
            .I(N__78968));
    Span4Mux_h I__18445 (
            .O(N__78976),
            .I(N__78968));
    LocalMux I__18444 (
            .O(N__78973),
            .I(\pid_side.error_i_reg_esr_RNIQ9ORZ0Z_15 ));
    Odrv4 I__18443 (
            .O(N__78968),
            .I(\pid_side.error_i_reg_esr_RNIQ9ORZ0Z_15 ));
    InMux I__18442 (
            .O(N__78963),
            .I(N__78960));
    LocalMux I__18441 (
            .O(N__78960),
            .I(N__78956));
    InMux I__18440 (
            .O(N__78959),
            .I(N__78953));
    Odrv4 I__18439 (
            .O(N__78956),
            .I(\pid_side.error_d_reg_prev_esr_RNI8UIO_0Z0Z_15 ));
    LocalMux I__18438 (
            .O(N__78953),
            .I(\pid_side.error_d_reg_prev_esr_RNI8UIO_0Z0Z_15 ));
    InMux I__18437 (
            .O(N__78948),
            .I(N__78942));
    InMux I__18436 (
            .O(N__78947),
            .I(N__78942));
    LocalMux I__18435 (
            .O(N__78942),
            .I(\pid_side.error_d_reg_prevZ0Z_15 ));
    InMux I__18434 (
            .O(N__78939),
            .I(N__78933));
    InMux I__18433 (
            .O(N__78938),
            .I(N__78933));
    LocalMux I__18432 (
            .O(N__78933),
            .I(N__78930));
    Odrv4 I__18431 (
            .O(N__78930),
            .I(\pid_side.error_d_reg_prev_esr_RNI8UIOZ0Z_15 ));
    InMux I__18430 (
            .O(N__78927),
            .I(N__78924));
    LocalMux I__18429 (
            .O(N__78924),
            .I(N__78921));
    Span4Mux_h I__18428 (
            .O(N__78921),
            .I(N__78918));
    Odrv4 I__18427 (
            .O(N__78918),
            .I(\pid_side.error_d_reg_prev_esr_RNIB8NBAZ0Z_12 ));
    CascadeMux I__18426 (
            .O(N__78915),
            .I(\pid_side.error_p_reg_esr_RNI4O091_0Z0Z_10_cascade_ ));
    InMux I__18425 (
            .O(N__78912),
            .I(N__78909));
    LocalMux I__18424 (
            .O(N__78909),
            .I(\pid_side.error_p_reg_esr_RNI4O091Z0Z_10 ));
    CascadeMux I__18423 (
            .O(N__78906),
            .I(\pid_side.error_d_reg_prev_esr_RNIV62K2Z0Z_10_cascade_ ));
    InMux I__18422 (
            .O(N__78903),
            .I(N__78900));
    LocalMux I__18421 (
            .O(N__78900),
            .I(N__78897));
    Span4Mux_v I__18420 (
            .O(N__78897),
            .I(N__78892));
    InMux I__18419 (
            .O(N__78896),
            .I(N__78889));
    InMux I__18418 (
            .O(N__78895),
            .I(N__78886));
    Span4Mux_h I__18417 (
            .O(N__78892),
            .I(N__78881));
    LocalMux I__18416 (
            .O(N__78889),
            .I(N__78881));
    LocalMux I__18415 (
            .O(N__78886),
            .I(\pid_side.error_d_reg_prev_esr_RNID3GT3_0Z0Z_10 ));
    Odrv4 I__18414 (
            .O(N__78881),
            .I(\pid_side.error_d_reg_prev_esr_RNID3GT3_0Z0Z_10 ));
    InMux I__18413 (
            .O(N__78876),
            .I(N__78871));
    InMux I__18412 (
            .O(N__78875),
            .I(N__78867));
    InMux I__18411 (
            .O(N__78874),
            .I(N__78864));
    LocalMux I__18410 (
            .O(N__78871),
            .I(N__78861));
    InMux I__18409 (
            .O(N__78870),
            .I(N__78858));
    LocalMux I__18408 (
            .O(N__78867),
            .I(N__78855));
    LocalMux I__18407 (
            .O(N__78864),
            .I(N__78852));
    Span4Mux_v I__18406 (
            .O(N__78861),
            .I(N__78849));
    LocalMux I__18405 (
            .O(N__78858),
            .I(N__78846));
    Span4Mux_v I__18404 (
            .O(N__78855),
            .I(N__78841));
    Span4Mux_v I__18403 (
            .O(N__78852),
            .I(N__78841));
    Span4Mux_h I__18402 (
            .O(N__78849),
            .I(N__78836));
    Span4Mux_v I__18401 (
            .O(N__78846),
            .I(N__78836));
    Odrv4 I__18400 (
            .O(N__78841),
            .I(\pid_side.error_i_reg_esr_RNIGRJRZ0Z_11 ));
    Odrv4 I__18399 (
            .O(N__78836),
            .I(\pid_side.error_i_reg_esr_RNIGRJRZ0Z_11 ));
    CascadeMux I__18398 (
            .O(N__78831),
            .I(\pid_side.un1_pid_prereg_153_0_cascade_ ));
    InMux I__18397 (
            .O(N__78828),
            .I(N__78825));
    LocalMux I__18396 (
            .O(N__78825),
            .I(N__78822));
    Odrv4 I__18395 (
            .O(N__78822),
            .I(\pid_side.error_d_reg_prev_esr_RNII28CBZ0Z_10 ));
    CascadeMux I__18394 (
            .O(N__78819),
            .I(N__78816));
    InMux I__18393 (
            .O(N__78816),
            .I(N__78807));
    InMux I__18392 (
            .O(N__78815),
            .I(N__78807));
    InMux I__18391 (
            .O(N__78814),
            .I(N__78807));
    LocalMux I__18390 (
            .O(N__78807),
            .I(N__78803));
    InMux I__18389 (
            .O(N__78806),
            .I(N__78800));
    Odrv4 I__18388 (
            .O(N__78803),
            .I(\pid_side.error_d_reg_prevZ0Z_10 ));
    LocalMux I__18387 (
            .O(N__78800),
            .I(\pid_side.error_d_reg_prevZ0Z_10 ));
    InMux I__18386 (
            .O(N__78795),
            .I(N__78792));
    LocalMux I__18385 (
            .O(N__78792),
            .I(\pid_side.error_d_reg_prev_esr_RNIV62K2Z0Z_10 ));
    InMux I__18384 (
            .O(N__78789),
            .I(N__78786));
    LocalMux I__18383 (
            .O(N__78786),
            .I(\pid_side.error_d_reg_prev_esr_RNID3GT3Z0Z_10 ));
    InMux I__18382 (
            .O(N__78783),
            .I(N__78778));
    InMux I__18381 (
            .O(N__78782),
            .I(N__78773));
    InMux I__18380 (
            .O(N__78781),
            .I(N__78773));
    LocalMux I__18379 (
            .O(N__78778),
            .I(N__78770));
    LocalMux I__18378 (
            .O(N__78773),
            .I(N__78767));
    Span4Mux_v I__18377 (
            .O(N__78770),
            .I(N__78762));
    Span4Mux_h I__18376 (
            .O(N__78767),
            .I(N__78762));
    Odrv4 I__18375 (
            .O(N__78762),
            .I(\pid_side.error_i_reg_esr_RNIJVKRZ0Z_12 ));
    InMux I__18374 (
            .O(N__78759),
            .I(N__78756));
    LocalMux I__18373 (
            .O(N__78756),
            .I(N__78753));
    Span4Mux_h I__18372 (
            .O(N__78753),
            .I(N__78749));
    InMux I__18371 (
            .O(N__78752),
            .I(N__78746));
    Odrv4 I__18370 (
            .O(N__78749),
            .I(\pid_side.error_d_reg_prev_esr_RNISSNM4Z0Z_12 ));
    LocalMux I__18369 (
            .O(N__78746),
            .I(\pid_side.error_d_reg_prev_esr_RNISSNM4Z0Z_12 ));
    CascadeMux I__18368 (
            .O(N__78741),
            .I(\pid_side.error_d_reg_prev_esr_RNID3GT3Z0Z_10_cascade_ ));
    CascadeMux I__18367 (
            .O(N__78738),
            .I(N__78735));
    InMux I__18366 (
            .O(N__78735),
            .I(N__78732));
    LocalMux I__18365 (
            .O(N__78732),
            .I(N__78729));
    Odrv4 I__18364 (
            .O(N__78729),
            .I(\pid_side.error_d_reg_prev_esr_RNIH0S9BZ0Z_10 ));
    InMux I__18363 (
            .O(N__78726),
            .I(N__78723));
    LocalMux I__18362 (
            .O(N__78723),
            .I(N__78720));
    Span4Mux_v I__18361 (
            .O(N__78720),
            .I(N__78717));
    Span4Mux_h I__18360 (
            .O(N__78717),
            .I(N__78714));
    Odrv4 I__18359 (
            .O(N__78714),
            .I(\pid_side.O_1_6 ));
    CEMux I__18358 (
            .O(N__78711),
            .I(N__78707));
    CEMux I__18357 (
            .O(N__78710),
            .I(N__78704));
    LocalMux I__18356 (
            .O(N__78707),
            .I(N__78700));
    LocalMux I__18355 (
            .O(N__78704),
            .I(N__78697));
    CEMux I__18354 (
            .O(N__78703),
            .I(N__78694));
    Span4Mux_v I__18353 (
            .O(N__78700),
            .I(N__78691));
    Span4Mux_h I__18352 (
            .O(N__78697),
            .I(N__78687));
    LocalMux I__18351 (
            .O(N__78694),
            .I(N__78684));
    Span4Mux_h I__18350 (
            .O(N__78691),
            .I(N__78681));
    CEMux I__18349 (
            .O(N__78690),
            .I(N__78678));
    Span4Mux_h I__18348 (
            .O(N__78687),
            .I(N__78675));
    Span4Mux_v I__18347 (
            .O(N__78684),
            .I(N__78672));
    Span4Mux_h I__18346 (
            .O(N__78681),
            .I(N__78667));
    LocalMux I__18345 (
            .O(N__78678),
            .I(N__78667));
    Span4Mux_h I__18344 (
            .O(N__78675),
            .I(N__78663));
    Span4Mux_v I__18343 (
            .O(N__78672),
            .I(N__78660));
    Span4Mux_v I__18342 (
            .O(N__78667),
            .I(N__78657));
    CEMux I__18341 (
            .O(N__78666),
            .I(N__78654));
    Span4Mux_h I__18340 (
            .O(N__78663),
            .I(N__78651));
    Span4Mux_h I__18339 (
            .O(N__78660),
            .I(N__78646));
    Span4Mux_v I__18338 (
            .O(N__78657),
            .I(N__78646));
    LocalMux I__18337 (
            .O(N__78654),
            .I(N__78643));
    Odrv4 I__18336 (
            .O(N__78651),
            .I(\Commands_frame_decoder.source_xy_ki_1_sqmuxa_0 ));
    Odrv4 I__18335 (
            .O(N__78646),
            .I(\Commands_frame_decoder.source_xy_ki_1_sqmuxa_0 ));
    Odrv4 I__18334 (
            .O(N__78643),
            .I(\Commands_frame_decoder.source_xy_ki_1_sqmuxa_0 ));
    CascadeMux I__18333 (
            .O(N__78636),
            .I(\pid_side.error_p_reg_esr_RNI76TK1_0Z0Z_5_cascade_ ));
    CascadeMux I__18332 (
            .O(N__78633),
            .I(N__78630));
    InMux I__18331 (
            .O(N__78630),
            .I(N__78627));
    LocalMux I__18330 (
            .O(N__78627),
            .I(N__78624));
    Odrv12 I__18329 (
            .O(N__78624),
            .I(\pid_side.error_p_reg_esr_RNIG7MC2Z0Z_5 ));
    InMux I__18328 (
            .O(N__78621),
            .I(N__78618));
    LocalMux I__18327 (
            .O(N__78618),
            .I(\pid_side.error_p_reg_esr_RNIIHEQZ0Z_4 ));
    CascadeMux I__18326 (
            .O(N__78615),
            .I(\pid_side.error_p_reg_esr_RNIIHEQZ0Z_4_cascade_ ));
    InMux I__18325 (
            .O(N__78612),
            .I(N__78602));
    InMux I__18324 (
            .O(N__78611),
            .I(N__78602));
    InMux I__18323 (
            .O(N__78610),
            .I(N__78602));
    InMux I__18322 (
            .O(N__78609),
            .I(N__78599));
    LocalMux I__18321 (
            .O(N__78602),
            .I(N__78596));
    LocalMux I__18320 (
            .O(N__78599),
            .I(\pid_side.error_d_reg_prevZ0Z_5 ));
    Odrv12 I__18319 (
            .O(N__78596),
            .I(\pid_side.error_d_reg_prevZ0Z_5 ));
    InMux I__18318 (
            .O(N__78591),
            .I(N__78588));
    LocalMux I__18317 (
            .O(N__78588),
            .I(N__78585));
    Span4Mux_h I__18316 (
            .O(N__78585),
            .I(N__78581));
    CascadeMux I__18315 (
            .O(N__78584),
            .I(N__78578));
    Span4Mux_h I__18314 (
            .O(N__78581),
            .I(N__78575));
    InMux I__18313 (
            .O(N__78578),
            .I(N__78572));
    Odrv4 I__18312 (
            .O(N__78575),
            .I(\pid_side.error_p_regZ0Z_6 ));
    LocalMux I__18311 (
            .O(N__78572),
            .I(\pid_side.error_p_regZ0Z_6 ));
    InMux I__18310 (
            .O(N__78567),
            .I(N__78564));
    LocalMux I__18309 (
            .O(N__78564),
            .I(N__78561));
    Span4Mux_h I__18308 (
            .O(N__78561),
            .I(N__78558));
    Span4Mux_h I__18307 (
            .O(N__78558),
            .I(N__78555));
    Odrv4 I__18306 (
            .O(N__78555),
            .I(\pid_side.N_2362_i ));
    InMux I__18305 (
            .O(N__78552),
            .I(N__78549));
    LocalMux I__18304 (
            .O(N__78549),
            .I(N__78546));
    Odrv4 I__18303 (
            .O(N__78546),
            .I(\pid_side.error_p_reg_esr_RNIIFTC1_0Z0Z_6 ));
    CascadeMux I__18302 (
            .O(N__78543),
            .I(\pid_side.error_p_reg_esr_RNIIFTC1_0Z0Z_6_cascade_ ));
    InMux I__18301 (
            .O(N__78540),
            .I(N__78535));
    InMux I__18300 (
            .O(N__78539),
            .I(N__78532));
    InMux I__18299 (
            .O(N__78538),
            .I(N__78529));
    LocalMux I__18298 (
            .O(N__78535),
            .I(N__78524));
    LocalMux I__18297 (
            .O(N__78532),
            .I(N__78524));
    LocalMux I__18296 (
            .O(N__78529),
            .I(N__78521));
    Span4Mux_h I__18295 (
            .O(N__78524),
            .I(N__78518));
    Odrv12 I__18294 (
            .O(N__78521),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_5_c_RNIC5QN ));
    Odrv4 I__18293 (
            .O(N__78518),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_5_c_RNIC5QN ));
    InMux I__18292 (
            .O(N__78513),
            .I(N__78507));
    InMux I__18291 (
            .O(N__78512),
            .I(N__78500));
    InMux I__18290 (
            .O(N__78511),
            .I(N__78500));
    InMux I__18289 (
            .O(N__78510),
            .I(N__78500));
    LocalMux I__18288 (
            .O(N__78507),
            .I(N__78497));
    LocalMux I__18287 (
            .O(N__78500),
            .I(N__78494));
    Span4Mux_v I__18286 (
            .O(N__78497),
            .I(N__78489));
    Span4Mux_h I__18285 (
            .O(N__78494),
            .I(N__78489));
    Odrv4 I__18284 (
            .O(N__78489),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_4_c_RNI91PN ));
    InMux I__18283 (
            .O(N__78486),
            .I(N__78482));
    InMux I__18282 (
            .O(N__78485),
            .I(N__78479));
    LocalMux I__18281 (
            .O(N__78482),
            .I(\pid_side.error_p_reg_esr_RNI76TK1_0Z0Z_5 ));
    LocalMux I__18280 (
            .O(N__78479),
            .I(\pid_side.error_p_reg_esr_RNI76TK1_0Z0Z_5 ));
    CascadeMux I__18279 (
            .O(N__78474),
            .I(\pid_side.un1_pid_prereg_66_0_cascade_ ));
    InMux I__18278 (
            .O(N__78471),
            .I(N__78468));
    LocalMux I__18277 (
            .O(N__78468),
            .I(N__78464));
    InMux I__18276 (
            .O(N__78467),
            .I(N__78461));
    Odrv4 I__18275 (
            .O(N__78464),
            .I(\pid_side.error_p_reg_esr_RNI76TK1Z0Z_5 ));
    LocalMux I__18274 (
            .O(N__78461),
            .I(\pid_side.error_p_reg_esr_RNI76TK1Z0Z_5 ));
    InMux I__18273 (
            .O(N__78456),
            .I(N__78453));
    LocalMux I__18272 (
            .O(N__78453),
            .I(N__78450));
    Odrv4 I__18271 (
            .O(N__78450),
            .I(\pid_side.error_p_reg_esr_RNIL2B66Z0Z_5 ));
    CascadeMux I__18270 (
            .O(N__78447),
            .I(N__78443));
    InMux I__18269 (
            .O(N__78446),
            .I(N__78436));
    InMux I__18268 (
            .O(N__78443),
            .I(N__78436));
    InMux I__18267 (
            .O(N__78442),
            .I(N__78431));
    InMux I__18266 (
            .O(N__78441),
            .I(N__78431));
    LocalMux I__18265 (
            .O(N__78436),
            .I(N__78428));
    LocalMux I__18264 (
            .O(N__78431),
            .I(\pid_side.error_d_reg_prevZ0Z_9 ));
    Odrv4 I__18263 (
            .O(N__78428),
            .I(\pid_side.error_d_reg_prevZ0Z_9 ));
    CascadeMux I__18262 (
            .O(N__78423),
            .I(N__78420));
    InMux I__18261 (
            .O(N__78420),
            .I(N__78412));
    CascadeMux I__18260 (
            .O(N__78419),
            .I(N__78408));
    InMux I__18259 (
            .O(N__78418),
            .I(N__78404));
    CascadeMux I__18258 (
            .O(N__78417),
            .I(N__78400));
    CascadeMux I__18257 (
            .O(N__78416),
            .I(N__78396));
    CascadeMux I__18256 (
            .O(N__78415),
            .I(N__78393));
    LocalMux I__18255 (
            .O(N__78412),
            .I(N__78390));
    InMux I__18254 (
            .O(N__78411),
            .I(N__78385));
    InMux I__18253 (
            .O(N__78408),
            .I(N__78385));
    CascadeMux I__18252 (
            .O(N__78407),
            .I(N__78382));
    LocalMux I__18251 (
            .O(N__78404),
            .I(N__78377));
    InMux I__18250 (
            .O(N__78403),
            .I(N__78374));
    InMux I__18249 (
            .O(N__78400),
            .I(N__78369));
    InMux I__18248 (
            .O(N__78399),
            .I(N__78366));
    InMux I__18247 (
            .O(N__78396),
            .I(N__78361));
    InMux I__18246 (
            .O(N__78393),
            .I(N__78361));
    Span4Mux_v I__18245 (
            .O(N__78390),
            .I(N__78354));
    LocalMux I__18244 (
            .O(N__78385),
            .I(N__78354));
    InMux I__18243 (
            .O(N__78382),
            .I(N__78351));
    CascadeMux I__18242 (
            .O(N__78381),
            .I(N__78348));
    InMux I__18241 (
            .O(N__78380),
            .I(N__78344));
    Span4Mux_v I__18240 (
            .O(N__78377),
            .I(N__78341));
    LocalMux I__18239 (
            .O(N__78374),
            .I(N__78338));
    CascadeMux I__18238 (
            .O(N__78373),
            .I(N__78335));
    CascadeMux I__18237 (
            .O(N__78372),
            .I(N__78331));
    LocalMux I__18236 (
            .O(N__78369),
            .I(N__78325));
    LocalMux I__18235 (
            .O(N__78366),
            .I(N__78325));
    LocalMux I__18234 (
            .O(N__78361),
            .I(N__78322));
    InMux I__18233 (
            .O(N__78360),
            .I(N__78317));
    InMux I__18232 (
            .O(N__78359),
            .I(N__78317));
    Span4Mux_h I__18231 (
            .O(N__78354),
            .I(N__78314));
    LocalMux I__18230 (
            .O(N__78351),
            .I(N__78311));
    InMux I__18229 (
            .O(N__78348),
            .I(N__78306));
    InMux I__18228 (
            .O(N__78347),
            .I(N__78306));
    LocalMux I__18227 (
            .O(N__78344),
            .I(N__78303));
    Span4Mux_v I__18226 (
            .O(N__78341),
            .I(N__78298));
    Span4Mux_h I__18225 (
            .O(N__78338),
            .I(N__78298));
    InMux I__18224 (
            .O(N__78335),
            .I(N__78293));
    InMux I__18223 (
            .O(N__78334),
            .I(N__78293));
    InMux I__18222 (
            .O(N__78331),
            .I(N__78288));
    InMux I__18221 (
            .O(N__78330),
            .I(N__78288));
    Span4Mux_v I__18220 (
            .O(N__78325),
            .I(N__78281));
    Span4Mux_v I__18219 (
            .O(N__78322),
            .I(N__78281));
    LocalMux I__18218 (
            .O(N__78317),
            .I(N__78281));
    Span4Mux_v I__18217 (
            .O(N__78314),
            .I(N__78278));
    Span4Mux_h I__18216 (
            .O(N__78311),
            .I(N__78271));
    LocalMux I__18215 (
            .O(N__78306),
            .I(N__78271));
    Span4Mux_h I__18214 (
            .O(N__78303),
            .I(N__78271));
    Span4Mux_h I__18213 (
            .O(N__78298),
            .I(N__78266));
    LocalMux I__18212 (
            .O(N__78293),
            .I(N__78266));
    LocalMux I__18211 (
            .O(N__78288),
            .I(N__78259));
    Span4Mux_h I__18210 (
            .O(N__78281),
            .I(N__78259));
    Span4Mux_h I__18209 (
            .O(N__78278),
            .I(N__78259));
    Odrv4 I__18208 (
            .O(N__78271),
            .I(xy_ki_0_rep2));
    Odrv4 I__18207 (
            .O(N__78266),
            .I(xy_ki_0_rep2));
    Odrv4 I__18206 (
            .O(N__78259),
            .I(xy_ki_0_rep2));
    InMux I__18205 (
            .O(N__78252),
            .I(N__78240));
    InMux I__18204 (
            .O(N__78251),
            .I(N__78235));
    InMux I__18203 (
            .O(N__78250),
            .I(N__78235));
    InMux I__18202 (
            .O(N__78249),
            .I(N__78232));
    InMux I__18201 (
            .O(N__78248),
            .I(N__78227));
    InMux I__18200 (
            .O(N__78247),
            .I(N__78227));
    InMux I__18199 (
            .O(N__78246),
            .I(N__78222));
    InMux I__18198 (
            .O(N__78245),
            .I(N__78222));
    InMux I__18197 (
            .O(N__78244),
            .I(N__78210));
    InMux I__18196 (
            .O(N__78243),
            .I(N__78205));
    LocalMux I__18195 (
            .O(N__78240),
            .I(N__78194));
    LocalMux I__18194 (
            .O(N__78235),
            .I(N__78194));
    LocalMux I__18193 (
            .O(N__78232),
            .I(N__78194));
    LocalMux I__18192 (
            .O(N__78227),
            .I(N__78194));
    LocalMux I__18191 (
            .O(N__78222),
            .I(N__78194));
    InMux I__18190 (
            .O(N__78221),
            .I(N__78191));
    InMux I__18189 (
            .O(N__78220),
            .I(N__78188));
    InMux I__18188 (
            .O(N__78219),
            .I(N__78185));
    InMux I__18187 (
            .O(N__78218),
            .I(N__78180));
    InMux I__18186 (
            .O(N__78217),
            .I(N__78180));
    InMux I__18185 (
            .O(N__78216),
            .I(N__78173));
    InMux I__18184 (
            .O(N__78215),
            .I(N__78173));
    InMux I__18183 (
            .O(N__78214),
            .I(N__78173));
    InMux I__18182 (
            .O(N__78213),
            .I(N__78170));
    LocalMux I__18181 (
            .O(N__78210),
            .I(N__78167));
    InMux I__18180 (
            .O(N__78209),
            .I(N__78163));
    InMux I__18179 (
            .O(N__78208),
            .I(N__78160));
    LocalMux I__18178 (
            .O(N__78205),
            .I(N__78157));
    Span4Mux_v I__18177 (
            .O(N__78194),
            .I(N__78152));
    LocalMux I__18176 (
            .O(N__78191),
            .I(N__78152));
    LocalMux I__18175 (
            .O(N__78188),
            .I(N__78143));
    LocalMux I__18174 (
            .O(N__78185),
            .I(N__78143));
    LocalMux I__18173 (
            .O(N__78180),
            .I(N__78143));
    LocalMux I__18172 (
            .O(N__78173),
            .I(N__78143));
    LocalMux I__18171 (
            .O(N__78170),
            .I(N__78140));
    Span4Mux_v I__18170 (
            .O(N__78167),
            .I(N__78137));
    InMux I__18169 (
            .O(N__78166),
            .I(N__78134));
    LocalMux I__18168 (
            .O(N__78163),
            .I(N__78131));
    LocalMux I__18167 (
            .O(N__78160),
            .I(N__78126));
    Span4Mux_h I__18166 (
            .O(N__78157),
            .I(N__78126));
    Span4Mux_h I__18165 (
            .O(N__78152),
            .I(N__78121));
    Span4Mux_h I__18164 (
            .O(N__78143),
            .I(N__78121));
    Span12Mux_v I__18163 (
            .O(N__78140),
            .I(N__78118));
    Odrv4 I__18162 (
            .O(N__78137),
            .I(xy_ki_fast_0));
    LocalMux I__18161 (
            .O(N__78134),
            .I(xy_ki_fast_0));
    Odrv4 I__18160 (
            .O(N__78131),
            .I(xy_ki_fast_0));
    Odrv4 I__18159 (
            .O(N__78126),
            .I(xy_ki_fast_0));
    Odrv4 I__18158 (
            .O(N__78121),
            .I(xy_ki_fast_0));
    Odrv12 I__18157 (
            .O(N__78118),
            .I(xy_ki_fast_0));
    CascadeMux I__18156 (
            .O(N__78105),
            .I(N__78100));
    CascadeMux I__18155 (
            .O(N__78104),
            .I(N__78094));
    CascadeMux I__18154 (
            .O(N__78103),
            .I(N__78086));
    InMux I__18153 (
            .O(N__78100),
            .I(N__78079));
    CascadeMux I__18152 (
            .O(N__78099),
            .I(N__78076));
    CascadeMux I__18151 (
            .O(N__78098),
            .I(N__78073));
    CascadeMux I__18150 (
            .O(N__78097),
            .I(N__78068));
    InMux I__18149 (
            .O(N__78094),
            .I(N__78065));
    CascadeMux I__18148 (
            .O(N__78093),
            .I(N__78062));
    CascadeMux I__18147 (
            .O(N__78092),
            .I(N__78058));
    InMux I__18146 (
            .O(N__78091),
            .I(N__78054));
    InMux I__18145 (
            .O(N__78090),
            .I(N__78047));
    InMux I__18144 (
            .O(N__78089),
            .I(N__78047));
    InMux I__18143 (
            .O(N__78086),
            .I(N__78047));
    CascadeMux I__18142 (
            .O(N__78085),
            .I(N__78042));
    CascadeMux I__18141 (
            .O(N__78084),
            .I(N__78036));
    CascadeMux I__18140 (
            .O(N__78083),
            .I(N__78032));
    InMux I__18139 (
            .O(N__78082),
            .I(N__78029));
    LocalMux I__18138 (
            .O(N__78079),
            .I(N__78026));
    InMux I__18137 (
            .O(N__78076),
            .I(N__78023));
    InMux I__18136 (
            .O(N__78073),
            .I(N__78018));
    InMux I__18135 (
            .O(N__78072),
            .I(N__78018));
    InMux I__18134 (
            .O(N__78071),
            .I(N__78015));
    InMux I__18133 (
            .O(N__78068),
            .I(N__78012));
    LocalMux I__18132 (
            .O(N__78065),
            .I(N__78009));
    InMux I__18131 (
            .O(N__78062),
            .I(N__78006));
    InMux I__18130 (
            .O(N__78061),
            .I(N__78001));
    InMux I__18129 (
            .O(N__78058),
            .I(N__78001));
    InMux I__18128 (
            .O(N__78057),
            .I(N__77998));
    LocalMux I__18127 (
            .O(N__78054),
            .I(N__77993));
    LocalMux I__18126 (
            .O(N__78047),
            .I(N__77993));
    InMux I__18125 (
            .O(N__78046),
            .I(N__77988));
    InMux I__18124 (
            .O(N__78045),
            .I(N__77988));
    InMux I__18123 (
            .O(N__78042),
            .I(N__77983));
    InMux I__18122 (
            .O(N__78041),
            .I(N__77983));
    InMux I__18121 (
            .O(N__78040),
            .I(N__77976));
    InMux I__18120 (
            .O(N__78039),
            .I(N__77976));
    InMux I__18119 (
            .O(N__78036),
            .I(N__77976));
    InMux I__18118 (
            .O(N__78035),
            .I(N__77971));
    InMux I__18117 (
            .O(N__78032),
            .I(N__77971));
    LocalMux I__18116 (
            .O(N__78029),
            .I(N__77964));
    Span4Mux_v I__18115 (
            .O(N__78026),
            .I(N__77964));
    LocalMux I__18114 (
            .O(N__78023),
            .I(N__77964));
    LocalMux I__18113 (
            .O(N__78018),
            .I(N__77961));
    LocalMux I__18112 (
            .O(N__78015),
            .I(N__77956));
    LocalMux I__18111 (
            .O(N__78012),
            .I(N__77956));
    Span4Mux_h I__18110 (
            .O(N__78009),
            .I(N__77953));
    LocalMux I__18109 (
            .O(N__78006),
            .I(N__77948));
    LocalMux I__18108 (
            .O(N__78001),
            .I(N__77948));
    LocalMux I__18107 (
            .O(N__77998),
            .I(N__77940));
    Span4Mux_v I__18106 (
            .O(N__77993),
            .I(N__77940));
    LocalMux I__18105 (
            .O(N__77988),
            .I(N__77940));
    LocalMux I__18104 (
            .O(N__77983),
            .I(N__77937));
    LocalMux I__18103 (
            .O(N__77976),
            .I(N__77930));
    LocalMux I__18102 (
            .O(N__77971),
            .I(N__77930));
    Span4Mux_h I__18101 (
            .O(N__77964),
            .I(N__77930));
    Span4Mux_v I__18100 (
            .O(N__77961),
            .I(N__77921));
    Span4Mux_v I__18099 (
            .O(N__77956),
            .I(N__77921));
    Span4Mux_v I__18098 (
            .O(N__77953),
            .I(N__77921));
    Span4Mux_h I__18097 (
            .O(N__77948),
            .I(N__77921));
    InMux I__18096 (
            .O(N__77947),
            .I(N__77918));
    Span4Mux_h I__18095 (
            .O(N__77940),
            .I(N__77915));
    Odrv4 I__18094 (
            .O(N__77937),
            .I(xy_ki_1_rep1));
    Odrv4 I__18093 (
            .O(N__77930),
            .I(xy_ki_1_rep1));
    Odrv4 I__18092 (
            .O(N__77921),
            .I(xy_ki_1_rep1));
    LocalMux I__18091 (
            .O(N__77918),
            .I(xy_ki_1_rep1));
    Odrv4 I__18090 (
            .O(N__77915),
            .I(xy_ki_1_rep1));
    CascadeMux I__18089 (
            .O(N__77904),
            .I(N__77898));
    InMux I__18088 (
            .O(N__77903),
            .I(N__77893));
    InMux I__18087 (
            .O(N__77902),
            .I(N__77886));
    InMux I__18086 (
            .O(N__77901),
            .I(N__77881));
    InMux I__18085 (
            .O(N__77898),
            .I(N__77881));
    CascadeMux I__18084 (
            .O(N__77897),
            .I(N__77878));
    CascadeMux I__18083 (
            .O(N__77896),
            .I(N__77875));
    LocalMux I__18082 (
            .O(N__77893),
            .I(N__77871));
    InMux I__18081 (
            .O(N__77892),
            .I(N__77868));
    InMux I__18080 (
            .O(N__77891),
            .I(N__77863));
    InMux I__18079 (
            .O(N__77890),
            .I(N__77863));
    InMux I__18078 (
            .O(N__77889),
            .I(N__77860));
    LocalMux I__18077 (
            .O(N__77886),
            .I(N__77855));
    LocalMux I__18076 (
            .O(N__77881),
            .I(N__77855));
    InMux I__18075 (
            .O(N__77878),
            .I(N__77850));
    InMux I__18074 (
            .O(N__77875),
            .I(N__77850));
    InMux I__18073 (
            .O(N__77874),
            .I(N__77846));
    Span4Mux_h I__18072 (
            .O(N__77871),
            .I(N__77841));
    LocalMux I__18071 (
            .O(N__77868),
            .I(N__77841));
    LocalMux I__18070 (
            .O(N__77863),
            .I(N__77838));
    LocalMux I__18069 (
            .O(N__77860),
            .I(N__77835));
    Span4Mux_v I__18068 (
            .O(N__77855),
            .I(N__77830));
    LocalMux I__18067 (
            .O(N__77850),
            .I(N__77830));
    CascadeMux I__18066 (
            .O(N__77849),
            .I(N__77827));
    LocalMux I__18065 (
            .O(N__77846),
            .I(N__77824));
    Span4Mux_v I__18064 (
            .O(N__77841),
            .I(N__77821));
    Span4Mux_h I__18063 (
            .O(N__77838),
            .I(N__77818));
    Span4Mux_v I__18062 (
            .O(N__77835),
            .I(N__77813));
    Span4Mux_h I__18061 (
            .O(N__77830),
            .I(N__77813));
    InMux I__18060 (
            .O(N__77827),
            .I(N__77810));
    Odrv12 I__18059 (
            .O(N__77824),
            .I(xy_ki_fast_1));
    Odrv4 I__18058 (
            .O(N__77821),
            .I(xy_ki_fast_1));
    Odrv4 I__18057 (
            .O(N__77818),
            .I(xy_ki_fast_1));
    Odrv4 I__18056 (
            .O(N__77813),
            .I(xy_ki_fast_1));
    LocalMux I__18055 (
            .O(N__77810),
            .I(xy_ki_fast_1));
    InMux I__18054 (
            .O(N__77799),
            .I(N__77796));
    LocalMux I__18053 (
            .O(N__77796),
            .I(N__77791));
    InMux I__18052 (
            .O(N__77795),
            .I(N__77788));
    CascadeMux I__18051 (
            .O(N__77794),
            .I(N__77784));
    Span4Mux_h I__18050 (
            .O(N__77791),
            .I(N__77774));
    LocalMux I__18049 (
            .O(N__77788),
            .I(N__77774));
    InMux I__18048 (
            .O(N__77787),
            .I(N__77771));
    InMux I__18047 (
            .O(N__77784),
            .I(N__77768));
    InMux I__18046 (
            .O(N__77783),
            .I(N__77764));
    CascadeMux I__18045 (
            .O(N__77782),
            .I(N__77756));
    CascadeMux I__18044 (
            .O(N__77781),
            .I(N__77752));
    InMux I__18043 (
            .O(N__77780),
            .I(N__77748));
    CascadeMux I__18042 (
            .O(N__77779),
            .I(N__77744));
    Span4Mux_h I__18041 (
            .O(N__77774),
            .I(N__77740));
    LocalMux I__18040 (
            .O(N__77771),
            .I(N__77731));
    LocalMux I__18039 (
            .O(N__77768),
            .I(N__77731));
    InMux I__18038 (
            .O(N__77767),
            .I(N__77728));
    LocalMux I__18037 (
            .O(N__77764),
            .I(N__77725));
    InMux I__18036 (
            .O(N__77763),
            .I(N__77720));
    InMux I__18035 (
            .O(N__77762),
            .I(N__77720));
    InMux I__18034 (
            .O(N__77761),
            .I(N__77715));
    InMux I__18033 (
            .O(N__77760),
            .I(N__77715));
    InMux I__18032 (
            .O(N__77759),
            .I(N__77710));
    InMux I__18031 (
            .O(N__77756),
            .I(N__77710));
    InMux I__18030 (
            .O(N__77755),
            .I(N__77705));
    InMux I__18029 (
            .O(N__77752),
            .I(N__77705));
    InMux I__18028 (
            .O(N__77751),
            .I(N__77700));
    LocalMux I__18027 (
            .O(N__77748),
            .I(N__77695));
    InMux I__18026 (
            .O(N__77747),
            .I(N__77688));
    InMux I__18025 (
            .O(N__77744),
            .I(N__77688));
    InMux I__18024 (
            .O(N__77743),
            .I(N__77688));
    Sp12to4 I__18023 (
            .O(N__77740),
            .I(N__77684));
    InMux I__18022 (
            .O(N__77739),
            .I(N__77678));
    InMux I__18021 (
            .O(N__77738),
            .I(N__77675));
    InMux I__18020 (
            .O(N__77737),
            .I(N__77670));
    InMux I__18019 (
            .O(N__77736),
            .I(N__77670));
    Span4Mux_v I__18018 (
            .O(N__77731),
            .I(N__77667));
    LocalMux I__18017 (
            .O(N__77728),
            .I(N__77662));
    Span4Mux_h I__18016 (
            .O(N__77725),
            .I(N__77662));
    LocalMux I__18015 (
            .O(N__77720),
            .I(N__77653));
    LocalMux I__18014 (
            .O(N__77715),
            .I(N__77653));
    LocalMux I__18013 (
            .O(N__77710),
            .I(N__77653));
    LocalMux I__18012 (
            .O(N__77705),
            .I(N__77653));
    InMux I__18011 (
            .O(N__77704),
            .I(N__77650));
    InMux I__18010 (
            .O(N__77703),
            .I(N__77647));
    LocalMux I__18009 (
            .O(N__77700),
            .I(N__77644));
    InMux I__18008 (
            .O(N__77699),
            .I(N__77639));
    InMux I__18007 (
            .O(N__77698),
            .I(N__77639));
    Span4Mux_h I__18006 (
            .O(N__77695),
            .I(N__77634));
    LocalMux I__18005 (
            .O(N__77688),
            .I(N__77634));
    InMux I__18004 (
            .O(N__77687),
            .I(N__77631));
    Span12Mux_v I__18003 (
            .O(N__77684),
            .I(N__77628));
    InMux I__18002 (
            .O(N__77683),
            .I(N__77621));
    InMux I__18001 (
            .O(N__77682),
            .I(N__77621));
    InMux I__18000 (
            .O(N__77681),
            .I(N__77621));
    LocalMux I__17999 (
            .O(N__77678),
            .I(N__77608));
    LocalMux I__17998 (
            .O(N__77675),
            .I(N__77608));
    LocalMux I__17997 (
            .O(N__77670),
            .I(N__77608));
    Span4Mux_h I__17996 (
            .O(N__77667),
            .I(N__77608));
    Span4Mux_v I__17995 (
            .O(N__77662),
            .I(N__77608));
    Span4Mux_v I__17994 (
            .O(N__77653),
            .I(N__77608));
    LocalMux I__17993 (
            .O(N__77650),
            .I(N__77599));
    LocalMux I__17992 (
            .O(N__77647),
            .I(N__77599));
    Span4Mux_v I__17991 (
            .O(N__77644),
            .I(N__77599));
    LocalMux I__17990 (
            .O(N__77639),
            .I(N__77599));
    Odrv4 I__17989 (
            .O(N__77634),
            .I(xy_ki_2_rep1));
    LocalMux I__17988 (
            .O(N__77631),
            .I(xy_ki_2_rep1));
    Odrv12 I__17987 (
            .O(N__77628),
            .I(xy_ki_2_rep1));
    LocalMux I__17986 (
            .O(N__77621),
            .I(xy_ki_2_rep1));
    Odrv4 I__17985 (
            .O(N__77608),
            .I(xy_ki_2_rep1));
    Odrv4 I__17984 (
            .O(N__77599),
            .I(xy_ki_2_rep1));
    InMux I__17983 (
            .O(N__77586),
            .I(N__77582));
    InMux I__17982 (
            .O(N__77585),
            .I(N__77579));
    LocalMux I__17981 (
            .O(N__77582),
            .I(N__77575));
    LocalMux I__17980 (
            .O(N__77579),
            .I(N__77567));
    InMux I__17979 (
            .O(N__77578),
            .I(N__77564));
    Span4Mux_v I__17978 (
            .O(N__77575),
            .I(N__77561));
    InMux I__17977 (
            .O(N__77574),
            .I(N__77558));
    InMux I__17976 (
            .O(N__77573),
            .I(N__77555));
    InMux I__17975 (
            .O(N__77572),
            .I(N__77550));
    InMux I__17974 (
            .O(N__77571),
            .I(N__77550));
    InMux I__17973 (
            .O(N__77570),
            .I(N__77543));
    Span4Mux_v I__17972 (
            .O(N__77567),
            .I(N__77538));
    LocalMux I__17971 (
            .O(N__77564),
            .I(N__77538));
    Span4Mux_h I__17970 (
            .O(N__77561),
            .I(N__77531));
    LocalMux I__17969 (
            .O(N__77558),
            .I(N__77531));
    LocalMux I__17968 (
            .O(N__77555),
            .I(N__77531));
    LocalMux I__17967 (
            .O(N__77550),
            .I(N__77528));
    InMux I__17966 (
            .O(N__77549),
            .I(N__77524));
    InMux I__17965 (
            .O(N__77548),
            .I(N__77521));
    InMux I__17964 (
            .O(N__77547),
            .I(N__77517));
    InMux I__17963 (
            .O(N__77546),
            .I(N__77514));
    LocalMux I__17962 (
            .O(N__77543),
            .I(N__77511));
    Span4Mux_v I__17961 (
            .O(N__77538),
            .I(N__77507));
    Span4Mux_v I__17960 (
            .O(N__77531),
            .I(N__77504));
    Span4Mux_v I__17959 (
            .O(N__77528),
            .I(N__77501));
    CascadeMux I__17958 (
            .O(N__77527),
            .I(N__77495));
    LocalMux I__17957 (
            .O(N__77524),
            .I(N__77492));
    LocalMux I__17956 (
            .O(N__77521),
            .I(N__77489));
    InMux I__17955 (
            .O(N__77520),
            .I(N__77486));
    LocalMux I__17954 (
            .O(N__77517),
            .I(N__77483));
    LocalMux I__17953 (
            .O(N__77514),
            .I(N__77480));
    Span4Mux_v I__17952 (
            .O(N__77511),
            .I(N__77477));
    InMux I__17951 (
            .O(N__77510),
            .I(N__77474));
    Sp12to4 I__17950 (
            .O(N__77507),
            .I(N__77467));
    Sp12to4 I__17949 (
            .O(N__77504),
            .I(N__77467));
    Sp12to4 I__17948 (
            .O(N__77501),
            .I(N__77467));
    InMux I__17947 (
            .O(N__77500),
            .I(N__77460));
    InMux I__17946 (
            .O(N__77499),
            .I(N__77460));
    InMux I__17945 (
            .O(N__77498),
            .I(N__77460));
    InMux I__17944 (
            .O(N__77495),
            .I(N__77456));
    Span4Mux_v I__17943 (
            .O(N__77492),
            .I(N__77453));
    Span4Mux_h I__17942 (
            .O(N__77489),
            .I(N__77450));
    LocalMux I__17941 (
            .O(N__77486),
            .I(N__77445));
    Span12Mux_v I__17940 (
            .O(N__77483),
            .I(N__77445));
    Span4Mux_v I__17939 (
            .O(N__77480),
            .I(N__77438));
    Span4Mux_v I__17938 (
            .O(N__77477),
            .I(N__77438));
    LocalMux I__17937 (
            .O(N__77474),
            .I(N__77438));
    Span12Mux_h I__17936 (
            .O(N__77467),
            .I(N__77435));
    LocalMux I__17935 (
            .O(N__77460),
            .I(N__77432));
    InMux I__17934 (
            .O(N__77459),
            .I(N__77429));
    LocalMux I__17933 (
            .O(N__77456),
            .I(uart_pc_data_2));
    Odrv4 I__17932 (
            .O(N__77453),
            .I(uart_pc_data_2));
    Odrv4 I__17931 (
            .O(N__77450),
            .I(uart_pc_data_2));
    Odrv12 I__17930 (
            .O(N__77445),
            .I(uart_pc_data_2));
    Odrv4 I__17929 (
            .O(N__77438),
            .I(uart_pc_data_2));
    Odrv12 I__17928 (
            .O(N__77435),
            .I(uart_pc_data_2));
    Odrv4 I__17927 (
            .O(N__77432),
            .I(uart_pc_data_2));
    LocalMux I__17926 (
            .O(N__77429),
            .I(uart_pc_data_2));
    CascadeMux I__17925 (
            .O(N__77412),
            .I(N__77407));
    InMux I__17924 (
            .O(N__77411),
            .I(N__77398));
    CascadeMux I__17923 (
            .O(N__77410),
            .I(N__77395));
    InMux I__17922 (
            .O(N__77407),
            .I(N__77387));
    InMux I__17921 (
            .O(N__77406),
            .I(N__77387));
    InMux I__17920 (
            .O(N__77405),
            .I(N__77383));
    InMux I__17919 (
            .O(N__77404),
            .I(N__77380));
    InMux I__17918 (
            .O(N__77403),
            .I(N__77377));
    InMux I__17917 (
            .O(N__77402),
            .I(N__77372));
    InMux I__17916 (
            .O(N__77401),
            .I(N__77372));
    LocalMux I__17915 (
            .O(N__77398),
            .I(N__77369));
    InMux I__17914 (
            .O(N__77395),
            .I(N__77366));
    InMux I__17913 (
            .O(N__77394),
            .I(N__77363));
    InMux I__17912 (
            .O(N__77393),
            .I(N__77360));
    InMux I__17911 (
            .O(N__77392),
            .I(N__77357));
    LocalMux I__17910 (
            .O(N__77387),
            .I(N__77354));
    InMux I__17909 (
            .O(N__77386),
            .I(N__77351));
    LocalMux I__17908 (
            .O(N__77383),
            .I(N__77348));
    LocalMux I__17907 (
            .O(N__77380),
            .I(N__77345));
    LocalMux I__17906 (
            .O(N__77377),
            .I(N__77342));
    LocalMux I__17905 (
            .O(N__77372),
            .I(N__77339));
    Span4Mux_h I__17904 (
            .O(N__77369),
            .I(N__77334));
    LocalMux I__17903 (
            .O(N__77366),
            .I(N__77334));
    LocalMux I__17902 (
            .O(N__77363),
            .I(N__77331));
    LocalMux I__17901 (
            .O(N__77360),
            .I(N__77328));
    LocalMux I__17900 (
            .O(N__77357),
            .I(N__77323));
    Span4Mux_h I__17899 (
            .O(N__77354),
            .I(N__77323));
    LocalMux I__17898 (
            .O(N__77351),
            .I(N__77320));
    Span4Mux_v I__17897 (
            .O(N__77348),
            .I(N__77315));
    Span4Mux_v I__17896 (
            .O(N__77345),
            .I(N__77315));
    Span4Mux_h I__17895 (
            .O(N__77342),
            .I(N__77310));
    Span4Mux_h I__17894 (
            .O(N__77339),
            .I(N__77310));
    Span4Mux_v I__17893 (
            .O(N__77334),
            .I(N__77301));
    Span4Mux_h I__17892 (
            .O(N__77331),
            .I(N__77301));
    Span4Mux_v I__17891 (
            .O(N__77328),
            .I(N__77301));
    Span4Mux_v I__17890 (
            .O(N__77323),
            .I(N__77301));
    Odrv12 I__17889 (
            .O(N__77320),
            .I(xy_ki_fast_2));
    Odrv4 I__17888 (
            .O(N__77315),
            .I(xy_ki_fast_2));
    Odrv4 I__17887 (
            .O(N__77310),
            .I(xy_ki_fast_2));
    Odrv4 I__17886 (
            .O(N__77301),
            .I(xy_ki_fast_2));
    InMux I__17885 (
            .O(N__77292),
            .I(N__77289));
    LocalMux I__17884 (
            .O(N__77289),
            .I(N__77286));
    Span12Mux_s10_v I__17883 (
            .O(N__77286),
            .I(N__77283));
    Odrv12 I__17882 (
            .O(N__77283),
            .I(\pid_side.O_2_9 ));
    InMux I__17881 (
            .O(N__77280),
            .I(N__77276));
    InMux I__17880 (
            .O(N__77279),
            .I(N__77273));
    LocalMux I__17879 (
            .O(N__77276),
            .I(N__77270));
    LocalMux I__17878 (
            .O(N__77273),
            .I(N__77267));
    Span4Mux_v I__17877 (
            .O(N__77270),
            .I(N__77264));
    Span4Mux_s2_h I__17876 (
            .O(N__77267),
            .I(N__77259));
    Span4Mux_h I__17875 (
            .O(N__77264),
            .I(N__77255));
    InMux I__17874 (
            .O(N__77263),
            .I(N__77252));
    InMux I__17873 (
            .O(N__77262),
            .I(N__77249));
    Span4Mux_h I__17872 (
            .O(N__77259),
            .I(N__77246));
    InMux I__17871 (
            .O(N__77258),
            .I(N__77243));
    Span4Mux_h I__17870 (
            .O(N__77255),
            .I(N__77240));
    LocalMux I__17869 (
            .O(N__77252),
            .I(N__77237));
    LocalMux I__17868 (
            .O(N__77249),
            .I(N__77234));
    Span4Mux_v I__17867 (
            .O(N__77246),
            .I(N__77227));
    LocalMux I__17866 (
            .O(N__77243),
            .I(N__77227));
    Span4Mux_h I__17865 (
            .O(N__77240),
            .I(N__77220));
    Span4Mux_v I__17864 (
            .O(N__77237),
            .I(N__77220));
    Span4Mux_v I__17863 (
            .O(N__77234),
            .I(N__77220));
    InMux I__17862 (
            .O(N__77233),
            .I(N__77215));
    InMux I__17861 (
            .O(N__77232),
            .I(N__77215));
    Span4Mux_h I__17860 (
            .O(N__77227),
            .I(N__77212));
    Odrv4 I__17859 (
            .O(N__77220),
            .I(drone_H_disp_front_0));
    LocalMux I__17858 (
            .O(N__77215),
            .I(drone_H_disp_front_0));
    Odrv4 I__17857 (
            .O(N__77212),
            .I(drone_H_disp_front_0));
    InMux I__17856 (
            .O(N__77205),
            .I(N__77201));
    InMux I__17855 (
            .O(N__77204),
            .I(N__77198));
    LocalMux I__17854 (
            .O(N__77201),
            .I(N__77195));
    LocalMux I__17853 (
            .O(N__77198),
            .I(N__77192));
    Span4Mux_h I__17852 (
            .O(N__77195),
            .I(N__77189));
    Span4Mux_s1_h I__17851 (
            .O(N__77192),
            .I(N__77186));
    Span4Mux_v I__17850 (
            .O(N__77189),
            .I(N__77182));
    Span4Mux_h I__17849 (
            .O(N__77186),
            .I(N__77179));
    InMux I__17848 (
            .O(N__77185),
            .I(N__77176));
    Span4Mux_h I__17847 (
            .O(N__77182),
            .I(N__77172));
    Span4Mux_h I__17846 (
            .O(N__77179),
            .I(N__77167));
    LocalMux I__17845 (
            .O(N__77176),
            .I(N__77167));
    InMux I__17844 (
            .O(N__77175),
            .I(N__77163));
    Span4Mux_h I__17843 (
            .O(N__77172),
            .I(N__77158));
    Span4Mux_v I__17842 (
            .O(N__77167),
            .I(N__77158));
    InMux I__17841 (
            .O(N__77166),
            .I(N__77155));
    LocalMux I__17840 (
            .O(N__77163),
            .I(N__77152));
    Odrv4 I__17839 (
            .O(N__77158),
            .I(\pid_front.error_1 ));
    LocalMux I__17838 (
            .O(N__77155),
            .I(\pid_front.error_1 ));
    Odrv12 I__17837 (
            .O(N__77152),
            .I(\pid_front.error_1 ));
    InMux I__17836 (
            .O(N__77145),
            .I(N__77142));
    LocalMux I__17835 (
            .O(N__77142),
            .I(N__77139));
    Sp12to4 I__17834 (
            .O(N__77139),
            .I(N__77135));
    InMux I__17833 (
            .O(N__77138),
            .I(N__77132));
    Span12Mux_v I__17832 (
            .O(N__77135),
            .I(N__77129));
    LocalMux I__17831 (
            .O(N__77132),
            .I(N__77126));
    Span12Mux_h I__17830 (
            .O(N__77129),
            .I(N__77120));
    Span12Mux_s7_v I__17829 (
            .O(N__77126),
            .I(N__77120));
    InMux I__17828 (
            .O(N__77125),
            .I(N__77115));
    Span12Mux_h I__17827 (
            .O(N__77120),
            .I(N__77112));
    InMux I__17826 (
            .O(N__77119),
            .I(N__77109));
    InMux I__17825 (
            .O(N__77118),
            .I(N__77106));
    LocalMux I__17824 (
            .O(N__77115),
            .I(N__77103));
    Odrv12 I__17823 (
            .O(N__77112),
            .I(\pid_front.error_2 ));
    LocalMux I__17822 (
            .O(N__77109),
            .I(\pid_front.error_2 ));
    LocalMux I__17821 (
            .O(N__77106),
            .I(\pid_front.error_2 ));
    Odrv12 I__17820 (
            .O(N__77103),
            .I(\pid_front.error_2 ));
    CascadeMux I__17819 (
            .O(N__77094),
            .I(\pid_front.m14_0_ns_1_cascade_ ));
    InMux I__17818 (
            .O(N__77091),
            .I(N__77087));
    InMux I__17817 (
            .O(N__77090),
            .I(N__77084));
    LocalMux I__17816 (
            .O(N__77087),
            .I(N__77081));
    LocalMux I__17815 (
            .O(N__77084),
            .I(N__77078));
    Span4Mux_h I__17814 (
            .O(N__77081),
            .I(N__77075));
    Span4Mux_s1_h I__17813 (
            .O(N__77078),
            .I(N__77072));
    Span4Mux_v I__17812 (
            .O(N__77075),
            .I(N__77068));
    Span4Mux_h I__17811 (
            .O(N__77072),
            .I(N__77064));
    InMux I__17810 (
            .O(N__77071),
            .I(N__77061));
    Span4Mux_h I__17809 (
            .O(N__77068),
            .I(N__77057));
    InMux I__17808 (
            .O(N__77067),
            .I(N__77054));
    Span4Mux_v I__17807 (
            .O(N__77064),
            .I(N__77049));
    LocalMux I__17806 (
            .O(N__77061),
            .I(N__77049));
    InMux I__17805 (
            .O(N__77060),
            .I(N__77046));
    Span4Mux_h I__17804 (
            .O(N__77057),
            .I(N__77039));
    LocalMux I__17803 (
            .O(N__77054),
            .I(N__77039));
    Span4Mux_h I__17802 (
            .O(N__77049),
            .I(N__77039));
    LocalMux I__17801 (
            .O(N__77046),
            .I(\pid_front.error_3 ));
    Odrv4 I__17800 (
            .O(N__77039),
            .I(\pid_front.error_3 ));
    CascadeMux I__17799 (
            .O(N__77034),
            .I(\pid_front.N_15_1_cascade_ ));
    CascadeMux I__17798 (
            .O(N__77031),
            .I(N__77026));
    CascadeMux I__17797 (
            .O(N__77030),
            .I(N__77019));
    CascadeMux I__17796 (
            .O(N__77029),
            .I(N__77015));
    InMux I__17795 (
            .O(N__77026),
            .I(N__77009));
    InMux I__17794 (
            .O(N__77025),
            .I(N__77006));
    InMux I__17793 (
            .O(N__77024),
            .I(N__76999));
    InMux I__17792 (
            .O(N__77023),
            .I(N__76994));
    InMux I__17791 (
            .O(N__77022),
            .I(N__76994));
    InMux I__17790 (
            .O(N__77019),
            .I(N__76991));
    CascadeMux I__17789 (
            .O(N__77018),
            .I(N__76987));
    InMux I__17788 (
            .O(N__77015),
            .I(N__76981));
    CascadeMux I__17787 (
            .O(N__77014),
            .I(N__76976));
    InMux I__17786 (
            .O(N__77013),
            .I(N__76971));
    InMux I__17785 (
            .O(N__77012),
            .I(N__76971));
    LocalMux I__17784 (
            .O(N__77009),
            .I(N__76968));
    LocalMux I__17783 (
            .O(N__77006),
            .I(N__76965));
    InMux I__17782 (
            .O(N__77005),
            .I(N__76962));
    CascadeMux I__17781 (
            .O(N__77004),
            .I(N__76956));
    InMux I__17780 (
            .O(N__77003),
            .I(N__76950));
    CascadeMux I__17779 (
            .O(N__77002),
            .I(N__76947));
    LocalMux I__17778 (
            .O(N__76999),
            .I(N__76934));
    LocalMux I__17777 (
            .O(N__76994),
            .I(N__76934));
    LocalMux I__17776 (
            .O(N__76991),
            .I(N__76934));
    InMux I__17775 (
            .O(N__76990),
            .I(N__76931));
    InMux I__17774 (
            .O(N__76987),
            .I(N__76926));
    InMux I__17773 (
            .O(N__76986),
            .I(N__76926));
    InMux I__17772 (
            .O(N__76985),
            .I(N__76923));
    CascadeMux I__17771 (
            .O(N__76984),
            .I(N__76920));
    LocalMux I__17770 (
            .O(N__76981),
            .I(N__76917));
    InMux I__17769 (
            .O(N__76980),
            .I(N__76914));
    InMux I__17768 (
            .O(N__76979),
            .I(N__76910));
    InMux I__17767 (
            .O(N__76976),
            .I(N__76907));
    LocalMux I__17766 (
            .O(N__76971),
            .I(N__76904));
    Span4Mux_v I__17765 (
            .O(N__76968),
            .I(N__76897));
    Span4Mux_h I__17764 (
            .O(N__76965),
            .I(N__76897));
    LocalMux I__17763 (
            .O(N__76962),
            .I(N__76897));
    InMux I__17762 (
            .O(N__76961),
            .I(N__76886));
    InMux I__17761 (
            .O(N__76960),
            .I(N__76886));
    InMux I__17760 (
            .O(N__76959),
            .I(N__76886));
    InMux I__17759 (
            .O(N__76956),
            .I(N__76886));
    InMux I__17758 (
            .O(N__76955),
            .I(N__76886));
    InMux I__17757 (
            .O(N__76954),
            .I(N__76879));
    InMux I__17756 (
            .O(N__76953),
            .I(N__76879));
    LocalMux I__17755 (
            .O(N__76950),
            .I(N__76876));
    InMux I__17754 (
            .O(N__76947),
            .I(N__76873));
    InMux I__17753 (
            .O(N__76946),
            .I(N__76870));
    InMux I__17752 (
            .O(N__76945),
            .I(N__76865));
    InMux I__17751 (
            .O(N__76944),
            .I(N__76860));
    InMux I__17750 (
            .O(N__76943),
            .I(N__76857));
    CascadeMux I__17749 (
            .O(N__76942),
            .I(N__76854));
    CascadeMux I__17748 (
            .O(N__76941),
            .I(N__76850));
    Span4Mux_v I__17747 (
            .O(N__76934),
            .I(N__76841));
    LocalMux I__17746 (
            .O(N__76931),
            .I(N__76841));
    LocalMux I__17745 (
            .O(N__76926),
            .I(N__76841));
    LocalMux I__17744 (
            .O(N__76923),
            .I(N__76841));
    InMux I__17743 (
            .O(N__76920),
            .I(N__76837));
    Span4Mux_h I__17742 (
            .O(N__76917),
            .I(N__76832));
    LocalMux I__17741 (
            .O(N__76914),
            .I(N__76832));
    InMux I__17740 (
            .O(N__76913),
            .I(N__76829));
    LocalMux I__17739 (
            .O(N__76910),
            .I(N__76818));
    LocalMux I__17738 (
            .O(N__76907),
            .I(N__76818));
    Span4Mux_h I__17737 (
            .O(N__76904),
            .I(N__76818));
    Span4Mux_v I__17736 (
            .O(N__76897),
            .I(N__76818));
    LocalMux I__17735 (
            .O(N__76886),
            .I(N__76818));
    InMux I__17734 (
            .O(N__76885),
            .I(N__76813));
    InMux I__17733 (
            .O(N__76884),
            .I(N__76813));
    LocalMux I__17732 (
            .O(N__76879),
            .I(N__76808));
    Span4Mux_h I__17731 (
            .O(N__76876),
            .I(N__76808));
    LocalMux I__17730 (
            .O(N__76873),
            .I(N__76805));
    LocalMux I__17729 (
            .O(N__76870),
            .I(N__76802));
    InMux I__17728 (
            .O(N__76869),
            .I(N__76799));
    InMux I__17727 (
            .O(N__76868),
            .I(N__76796));
    LocalMux I__17726 (
            .O(N__76865),
            .I(N__76793));
    InMux I__17725 (
            .O(N__76864),
            .I(N__76790));
    InMux I__17724 (
            .O(N__76863),
            .I(N__76785));
    LocalMux I__17723 (
            .O(N__76860),
            .I(N__76780));
    LocalMux I__17722 (
            .O(N__76857),
            .I(N__76780));
    InMux I__17721 (
            .O(N__76854),
            .I(N__76773));
    InMux I__17720 (
            .O(N__76853),
            .I(N__76773));
    InMux I__17719 (
            .O(N__76850),
            .I(N__76773));
    Span4Mux_h I__17718 (
            .O(N__76841),
            .I(N__76770));
    InMux I__17717 (
            .O(N__76840),
            .I(N__76767));
    LocalMux I__17716 (
            .O(N__76837),
            .I(N__76756));
    Span4Mux_v I__17715 (
            .O(N__76832),
            .I(N__76756));
    LocalMux I__17714 (
            .O(N__76829),
            .I(N__76756));
    Span4Mux_v I__17713 (
            .O(N__76818),
            .I(N__76756));
    LocalMux I__17712 (
            .O(N__76813),
            .I(N__76756));
    Span4Mux_h I__17711 (
            .O(N__76808),
            .I(N__76753));
    Span4Mux_h I__17710 (
            .O(N__76805),
            .I(N__76750));
    Span4Mux_v I__17709 (
            .O(N__76802),
            .I(N__76747));
    LocalMux I__17708 (
            .O(N__76799),
            .I(N__76742));
    LocalMux I__17707 (
            .O(N__76796),
            .I(N__76742));
    Span4Mux_v I__17706 (
            .O(N__76793),
            .I(N__76737));
    LocalMux I__17705 (
            .O(N__76790),
            .I(N__76737));
    InMux I__17704 (
            .O(N__76789),
            .I(N__76732));
    InMux I__17703 (
            .O(N__76788),
            .I(N__76732));
    LocalMux I__17702 (
            .O(N__76785),
            .I(N__76727));
    Span4Mux_v I__17701 (
            .O(N__76780),
            .I(N__76727));
    LocalMux I__17700 (
            .O(N__76773),
            .I(N__76724));
    Span4Mux_h I__17699 (
            .O(N__76770),
            .I(N__76721));
    LocalMux I__17698 (
            .O(N__76767),
            .I(N__76716));
    Span4Mux_v I__17697 (
            .O(N__76756),
            .I(N__76716));
    Span4Mux_h I__17696 (
            .O(N__76753),
            .I(N__76711));
    Span4Mux_h I__17695 (
            .O(N__76750),
            .I(N__76711));
    Span4Mux_h I__17694 (
            .O(N__76747),
            .I(N__76706));
    Span4Mux_v I__17693 (
            .O(N__76742),
            .I(N__76706));
    Span4Mux_v I__17692 (
            .O(N__76737),
            .I(N__76701));
    LocalMux I__17691 (
            .O(N__76732),
            .I(N__76701));
    Span4Mux_h I__17690 (
            .O(N__76727),
            .I(N__76696));
    Span4Mux_h I__17689 (
            .O(N__76724),
            .I(N__76696));
    Span4Mux_h I__17688 (
            .O(N__76721),
            .I(N__76693));
    Span4Mux_v I__17687 (
            .O(N__76716),
            .I(N__76690));
    Sp12to4 I__17686 (
            .O(N__76711),
            .I(N__76687));
    Span4Mux_h I__17685 (
            .O(N__76706),
            .I(N__76684));
    Span4Mux_h I__17684 (
            .O(N__76701),
            .I(N__76681));
    Span4Mux_h I__17683 (
            .O(N__76696),
            .I(N__76676));
    Span4Mux_v I__17682 (
            .O(N__76693),
            .I(N__76676));
    Sp12to4 I__17681 (
            .O(N__76690),
            .I(N__76673));
    Span12Mux_v I__17680 (
            .O(N__76687),
            .I(N__76670));
    Odrv4 I__17679 (
            .O(N__76684),
            .I(xy_ki_4));
    Odrv4 I__17678 (
            .O(N__76681),
            .I(xy_ki_4));
    Odrv4 I__17677 (
            .O(N__76676),
            .I(xy_ki_4));
    Odrv12 I__17676 (
            .O(N__76673),
            .I(xy_ki_4));
    Odrv12 I__17675 (
            .O(N__76670),
            .I(xy_ki_4));
    InMux I__17674 (
            .O(N__76659),
            .I(N__76652));
    InMux I__17673 (
            .O(N__76658),
            .I(N__76643));
    InMux I__17672 (
            .O(N__76657),
            .I(N__76643));
    InMux I__17671 (
            .O(N__76656),
            .I(N__76643));
    InMux I__17670 (
            .O(N__76655),
            .I(N__76643));
    LocalMux I__17669 (
            .O(N__76652),
            .I(N__76632));
    LocalMux I__17668 (
            .O(N__76643),
            .I(N__76632));
    InMux I__17667 (
            .O(N__76642),
            .I(N__76625));
    InMux I__17666 (
            .O(N__76641),
            .I(N__76619));
    InMux I__17665 (
            .O(N__76640),
            .I(N__76619));
    InMux I__17664 (
            .O(N__76639),
            .I(N__76612));
    InMux I__17663 (
            .O(N__76638),
            .I(N__76606));
    InMux I__17662 (
            .O(N__76637),
            .I(N__76606));
    Span4Mux_h I__17661 (
            .O(N__76632),
            .I(N__76602));
    InMux I__17660 (
            .O(N__76631),
            .I(N__76597));
    InMux I__17659 (
            .O(N__76630),
            .I(N__76597));
    InMux I__17658 (
            .O(N__76629),
            .I(N__76594));
    InMux I__17657 (
            .O(N__76628),
            .I(N__76591));
    LocalMux I__17656 (
            .O(N__76625),
            .I(N__76588));
    InMux I__17655 (
            .O(N__76624),
            .I(N__76585));
    LocalMux I__17654 (
            .O(N__76619),
            .I(N__76582));
    InMux I__17653 (
            .O(N__76618),
            .I(N__76578));
    InMux I__17652 (
            .O(N__76617),
            .I(N__76573));
    InMux I__17651 (
            .O(N__76616),
            .I(N__76573));
    InMux I__17650 (
            .O(N__76615),
            .I(N__76569));
    LocalMux I__17649 (
            .O(N__76612),
            .I(N__76566));
    InMux I__17648 (
            .O(N__76611),
            .I(N__76563));
    LocalMux I__17647 (
            .O(N__76606),
            .I(N__76560));
    InMux I__17646 (
            .O(N__76605),
            .I(N__76554));
    Span4Mux_v I__17645 (
            .O(N__76602),
            .I(N__76541));
    LocalMux I__17644 (
            .O(N__76597),
            .I(N__76536));
    LocalMux I__17643 (
            .O(N__76594),
            .I(N__76536));
    LocalMux I__17642 (
            .O(N__76591),
            .I(N__76526));
    Span4Mux_v I__17641 (
            .O(N__76588),
            .I(N__76526));
    LocalMux I__17640 (
            .O(N__76585),
            .I(N__76526));
    Span4Mux_h I__17639 (
            .O(N__76582),
            .I(N__76526));
    InMux I__17638 (
            .O(N__76581),
            .I(N__76523));
    LocalMux I__17637 (
            .O(N__76578),
            .I(N__76518));
    LocalMux I__17636 (
            .O(N__76573),
            .I(N__76518));
    InMux I__17635 (
            .O(N__76572),
            .I(N__76515));
    LocalMux I__17634 (
            .O(N__76569),
            .I(N__76510));
    Span4Mux_h I__17633 (
            .O(N__76566),
            .I(N__76507));
    LocalMux I__17632 (
            .O(N__76563),
            .I(N__76504));
    Span4Mux_h I__17631 (
            .O(N__76560),
            .I(N__76501));
    InMux I__17630 (
            .O(N__76559),
            .I(N__76496));
    InMux I__17629 (
            .O(N__76558),
            .I(N__76496));
    InMux I__17628 (
            .O(N__76557),
            .I(N__76493));
    LocalMux I__17627 (
            .O(N__76554),
            .I(N__76490));
    InMux I__17626 (
            .O(N__76553),
            .I(N__76487));
    InMux I__17625 (
            .O(N__76552),
            .I(N__76484));
    InMux I__17624 (
            .O(N__76551),
            .I(N__76473));
    InMux I__17623 (
            .O(N__76550),
            .I(N__76473));
    InMux I__17622 (
            .O(N__76549),
            .I(N__76473));
    InMux I__17621 (
            .O(N__76548),
            .I(N__76473));
    InMux I__17620 (
            .O(N__76547),
            .I(N__76473));
    InMux I__17619 (
            .O(N__76546),
            .I(N__76466));
    InMux I__17618 (
            .O(N__76545),
            .I(N__76466));
    InMux I__17617 (
            .O(N__76544),
            .I(N__76466));
    Span4Mux_h I__17616 (
            .O(N__76541),
            .I(N__76461));
    Span4Mux_h I__17615 (
            .O(N__76536),
            .I(N__76461));
    InMux I__17614 (
            .O(N__76535),
            .I(N__76458));
    Span4Mux_v I__17613 (
            .O(N__76526),
            .I(N__76455));
    LocalMux I__17612 (
            .O(N__76523),
            .I(N__76450));
    Span4Mux_h I__17611 (
            .O(N__76518),
            .I(N__76450));
    LocalMux I__17610 (
            .O(N__76515),
            .I(N__76447));
    InMux I__17609 (
            .O(N__76514),
            .I(N__76444));
    InMux I__17608 (
            .O(N__76513),
            .I(N__76441));
    Span4Mux_v I__17607 (
            .O(N__76510),
            .I(N__76430));
    Span4Mux_v I__17606 (
            .O(N__76507),
            .I(N__76430));
    Span4Mux_h I__17605 (
            .O(N__76504),
            .I(N__76430));
    Span4Mux_v I__17604 (
            .O(N__76501),
            .I(N__76430));
    LocalMux I__17603 (
            .O(N__76496),
            .I(N__76430));
    LocalMux I__17602 (
            .O(N__76493),
            .I(N__76423));
    Span4Mux_v I__17601 (
            .O(N__76490),
            .I(N__76423));
    LocalMux I__17600 (
            .O(N__76487),
            .I(N__76423));
    LocalMux I__17599 (
            .O(N__76484),
            .I(N__76414));
    LocalMux I__17598 (
            .O(N__76473),
            .I(N__76414));
    LocalMux I__17597 (
            .O(N__76466),
            .I(N__76414));
    Sp12to4 I__17596 (
            .O(N__76461),
            .I(N__76414));
    LocalMux I__17595 (
            .O(N__76458),
            .I(pid_front_N_331));
    Odrv4 I__17594 (
            .O(N__76455),
            .I(pid_front_N_331));
    Odrv4 I__17593 (
            .O(N__76450),
            .I(pid_front_N_331));
    Odrv4 I__17592 (
            .O(N__76447),
            .I(pid_front_N_331));
    LocalMux I__17591 (
            .O(N__76444),
            .I(pid_front_N_331));
    LocalMux I__17590 (
            .O(N__76441),
            .I(pid_front_N_331));
    Odrv4 I__17589 (
            .O(N__76430),
            .I(pid_front_N_331));
    Odrv4 I__17588 (
            .O(N__76423),
            .I(pid_front_N_331));
    Odrv12 I__17587 (
            .O(N__76414),
            .I(pid_front_N_331));
    CascadeMux I__17586 (
            .O(N__76395),
            .I(\pid_front.m3_2_03_cascade_ ));
    InMux I__17585 (
            .O(N__76392),
            .I(N__76386));
    InMux I__17584 (
            .O(N__76391),
            .I(N__76386));
    LocalMux I__17583 (
            .O(N__76386),
            .I(\pid_front.error_i_reg_9_rn_rn_2_15 ));
    CascadeMux I__17582 (
            .O(N__76383),
            .I(N__76379));
    InMux I__17581 (
            .O(N__76382),
            .I(N__76376));
    InMux I__17580 (
            .O(N__76379),
            .I(N__76373));
    LocalMux I__17579 (
            .O(N__76376),
            .I(N__76369));
    LocalMux I__17578 (
            .O(N__76373),
            .I(N__76366));
    InMux I__17577 (
            .O(N__76372),
            .I(N__76363));
    Span4Mux_h I__17576 (
            .O(N__76369),
            .I(N__76359));
    Span4Mux_v I__17575 (
            .O(N__76366),
            .I(N__76354));
    LocalMux I__17574 (
            .O(N__76363),
            .I(N__76354));
    InMux I__17573 (
            .O(N__76362),
            .I(N__76351));
    Odrv4 I__17572 (
            .O(N__76359),
            .I(\pid_front.N_15_1 ));
    Odrv4 I__17571 (
            .O(N__76354),
            .I(\pid_front.N_15_1 ));
    LocalMux I__17570 (
            .O(N__76351),
            .I(\pid_front.N_15_1 ));
    InMux I__17569 (
            .O(N__76344),
            .I(N__76341));
    LocalMux I__17568 (
            .O(N__76341),
            .I(N__76338));
    Span4Mux_h I__17567 (
            .O(N__76338),
            .I(N__76334));
    InMux I__17566 (
            .O(N__76337),
            .I(N__76331));
    Odrv4 I__17565 (
            .O(N__76334),
            .I(\pid_front.N_104 ));
    LocalMux I__17564 (
            .O(N__76331),
            .I(\pid_front.N_104 ));
    CascadeMux I__17563 (
            .O(N__76326),
            .I(N__76323));
    InMux I__17562 (
            .O(N__76323),
            .I(N__76315));
    CascadeMux I__17561 (
            .O(N__76322),
            .I(N__76312));
    InMux I__17560 (
            .O(N__76321),
            .I(N__76305));
    InMux I__17559 (
            .O(N__76320),
            .I(N__76305));
    CascadeMux I__17558 (
            .O(N__76319),
            .I(N__76302));
    InMux I__17557 (
            .O(N__76318),
            .I(N__76295));
    LocalMux I__17556 (
            .O(N__76315),
            .I(N__76292));
    InMux I__17555 (
            .O(N__76312),
            .I(N__76287));
    InMux I__17554 (
            .O(N__76311),
            .I(N__76287));
    CascadeMux I__17553 (
            .O(N__76310),
            .I(N__76283));
    LocalMux I__17552 (
            .O(N__76305),
            .I(N__76276));
    InMux I__17551 (
            .O(N__76302),
            .I(N__76273));
    InMux I__17550 (
            .O(N__76301),
            .I(N__76264));
    InMux I__17549 (
            .O(N__76300),
            .I(N__76261));
    InMux I__17548 (
            .O(N__76299),
            .I(N__76258));
    InMux I__17547 (
            .O(N__76298),
            .I(N__76255));
    LocalMux I__17546 (
            .O(N__76295),
            .I(N__76248));
    Span4Mux_v I__17545 (
            .O(N__76292),
            .I(N__76248));
    LocalMux I__17544 (
            .O(N__76287),
            .I(N__76248));
    InMux I__17543 (
            .O(N__76286),
            .I(N__76243));
    InMux I__17542 (
            .O(N__76283),
            .I(N__76243));
    InMux I__17541 (
            .O(N__76282),
            .I(N__76238));
    InMux I__17540 (
            .O(N__76281),
            .I(N__76235));
    InMux I__17539 (
            .O(N__76280),
            .I(N__76230));
    InMux I__17538 (
            .O(N__76279),
            .I(N__76230));
    Span4Mux_v I__17537 (
            .O(N__76276),
            .I(N__76227));
    LocalMux I__17536 (
            .O(N__76273),
            .I(N__76224));
    InMux I__17535 (
            .O(N__76272),
            .I(N__76221));
    InMux I__17534 (
            .O(N__76271),
            .I(N__76218));
    InMux I__17533 (
            .O(N__76270),
            .I(N__76215));
    InMux I__17532 (
            .O(N__76269),
            .I(N__76212));
    CascadeMux I__17531 (
            .O(N__76268),
            .I(N__76209));
    InMux I__17530 (
            .O(N__76267),
            .I(N__76205));
    LocalMux I__17529 (
            .O(N__76264),
            .I(N__76200));
    LocalMux I__17528 (
            .O(N__76261),
            .I(N__76200));
    LocalMux I__17527 (
            .O(N__76258),
            .I(N__76197));
    LocalMux I__17526 (
            .O(N__76255),
            .I(N__76194));
    Span4Mux_h I__17525 (
            .O(N__76248),
            .I(N__76191));
    LocalMux I__17524 (
            .O(N__76243),
            .I(N__76188));
    InMux I__17523 (
            .O(N__76242),
            .I(N__76185));
    InMux I__17522 (
            .O(N__76241),
            .I(N__76182));
    LocalMux I__17521 (
            .O(N__76238),
            .I(N__76171));
    LocalMux I__17520 (
            .O(N__76235),
            .I(N__76171));
    LocalMux I__17519 (
            .O(N__76230),
            .I(N__76171));
    Span4Mux_h I__17518 (
            .O(N__76227),
            .I(N__76171));
    Span4Mux_h I__17517 (
            .O(N__76224),
            .I(N__76171));
    LocalMux I__17516 (
            .O(N__76221),
            .I(N__76162));
    LocalMux I__17515 (
            .O(N__76218),
            .I(N__76162));
    LocalMux I__17514 (
            .O(N__76215),
            .I(N__76162));
    LocalMux I__17513 (
            .O(N__76212),
            .I(N__76162));
    InMux I__17512 (
            .O(N__76209),
            .I(N__76157));
    InMux I__17511 (
            .O(N__76208),
            .I(N__76157));
    LocalMux I__17510 (
            .O(N__76205),
            .I(N__76154));
    Span4Mux_v I__17509 (
            .O(N__76200),
            .I(N__76149));
    Span4Mux_h I__17508 (
            .O(N__76197),
            .I(N__76149));
    Span4Mux_v I__17507 (
            .O(N__76194),
            .I(N__76142));
    Span4Mux_v I__17506 (
            .O(N__76191),
            .I(N__76142));
    Span4Mux_h I__17505 (
            .O(N__76188),
            .I(N__76142));
    LocalMux I__17504 (
            .O(N__76185),
            .I(N__76139));
    LocalMux I__17503 (
            .O(N__76182),
            .I(N__76136));
    Span4Mux_v I__17502 (
            .O(N__76171),
            .I(N__76129));
    Span4Mux_v I__17501 (
            .O(N__76162),
            .I(N__76129));
    LocalMux I__17500 (
            .O(N__76157),
            .I(N__76129));
    Span4Mux_h I__17499 (
            .O(N__76154),
            .I(N__76126));
    Span4Mux_h I__17498 (
            .O(N__76149),
            .I(N__76121));
    Span4Mux_h I__17497 (
            .O(N__76142),
            .I(N__76121));
    Span4Mux_h I__17496 (
            .O(N__76139),
            .I(N__76116));
    Span4Mux_h I__17495 (
            .O(N__76136),
            .I(N__76116));
    Span4Mux_h I__17494 (
            .O(N__76129),
            .I(N__76113));
    Span4Mux_v I__17493 (
            .O(N__76126),
            .I(N__76108));
    Span4Mux_v I__17492 (
            .O(N__76121),
            .I(N__76108));
    Odrv4 I__17491 (
            .O(N__76116),
            .I(xy_ki_3_rep2));
    Odrv4 I__17490 (
            .O(N__76113),
            .I(xy_ki_3_rep2));
    Odrv4 I__17489 (
            .O(N__76108),
            .I(xy_ki_3_rep2));
    CascadeMux I__17488 (
            .O(N__76101),
            .I(\pid_front.N_104_cascade_ ));
    InMux I__17487 (
            .O(N__76098),
            .I(N__76086));
    InMux I__17486 (
            .O(N__76097),
            .I(N__76086));
    InMux I__17485 (
            .O(N__76096),
            .I(N__76086));
    InMux I__17484 (
            .O(N__76095),
            .I(N__76083));
    InMux I__17483 (
            .O(N__76094),
            .I(N__76078));
    InMux I__17482 (
            .O(N__76093),
            .I(N__76078));
    LocalMux I__17481 (
            .O(N__76086),
            .I(N__76075));
    LocalMux I__17480 (
            .O(N__76083),
            .I(\pid_front.N_39_0 ));
    LocalMux I__17479 (
            .O(N__76078),
            .I(\pid_front.N_39_0 ));
    Odrv4 I__17478 (
            .O(N__76075),
            .I(\pid_front.N_39_0 ));
    InMux I__17477 (
            .O(N__76068),
            .I(N__76063));
    InMux I__17476 (
            .O(N__76067),
            .I(N__76055));
    InMux I__17475 (
            .O(N__76066),
            .I(N__76055));
    LocalMux I__17474 (
            .O(N__76063),
            .I(N__76051));
    InMux I__17473 (
            .O(N__76062),
            .I(N__76048));
    InMux I__17472 (
            .O(N__76061),
            .I(N__76043));
    InMux I__17471 (
            .O(N__76060),
            .I(N__76043));
    LocalMux I__17470 (
            .O(N__76055),
            .I(N__76040));
    InMux I__17469 (
            .O(N__76054),
            .I(N__76037));
    Odrv4 I__17468 (
            .O(N__76051),
            .I(\pid_front.N_49_0 ));
    LocalMux I__17467 (
            .O(N__76048),
            .I(\pid_front.N_49_0 ));
    LocalMux I__17466 (
            .O(N__76043),
            .I(\pid_front.N_49_0 ));
    Odrv4 I__17465 (
            .O(N__76040),
            .I(\pid_front.N_49_0 ));
    LocalMux I__17464 (
            .O(N__76037),
            .I(\pid_front.N_49_0 ));
    CascadeMux I__17463 (
            .O(N__76026),
            .I(\pid_front.error_i_reg_esr_RNO_2Z0Z_23_cascade_ ));
    InMux I__17462 (
            .O(N__76023),
            .I(N__76020));
    LocalMux I__17461 (
            .O(N__76020),
            .I(\pid_front.error_i_reg_esr_RNO_3Z0Z_23 ));
    InMux I__17460 (
            .O(N__76017),
            .I(N__76014));
    LocalMux I__17459 (
            .O(N__76014),
            .I(\pid_front.error_i_reg_esr_RNO_1_0_23 ));
    CascadeMux I__17458 (
            .O(N__76011),
            .I(N__76006));
    InMux I__17457 (
            .O(N__76010),
            .I(N__76002));
    InMux I__17456 (
            .O(N__76009),
            .I(N__75999));
    InMux I__17455 (
            .O(N__76006),
            .I(N__75990));
    InMux I__17454 (
            .O(N__76005),
            .I(N__75990));
    LocalMux I__17453 (
            .O(N__76002),
            .I(N__75985));
    LocalMux I__17452 (
            .O(N__75999),
            .I(N__75985));
    CascadeMux I__17451 (
            .O(N__75998),
            .I(N__75981));
    InMux I__17450 (
            .O(N__75997),
            .I(N__75974));
    InMux I__17449 (
            .O(N__75996),
            .I(N__75974));
    InMux I__17448 (
            .O(N__75995),
            .I(N__75974));
    LocalMux I__17447 (
            .O(N__75990),
            .I(N__75969));
    Span4Mux_v I__17446 (
            .O(N__75985),
            .I(N__75969));
    InMux I__17445 (
            .O(N__75984),
            .I(N__75965));
    InMux I__17444 (
            .O(N__75981),
            .I(N__75959));
    LocalMux I__17443 (
            .O(N__75974),
            .I(N__75956));
    Span4Mux_v I__17442 (
            .O(N__75969),
            .I(N__75953));
    InMux I__17441 (
            .O(N__75968),
            .I(N__75950));
    LocalMux I__17440 (
            .O(N__75965),
            .I(N__75947));
    InMux I__17439 (
            .O(N__75964),
            .I(N__75944));
    InMux I__17438 (
            .O(N__75963),
            .I(N__75939));
    InMux I__17437 (
            .O(N__75962),
            .I(N__75939));
    LocalMux I__17436 (
            .O(N__75959),
            .I(N__75936));
    Span4Mux_h I__17435 (
            .O(N__75956),
            .I(N__75933));
    Span4Mux_h I__17434 (
            .O(N__75953),
            .I(N__75930));
    LocalMux I__17433 (
            .O(N__75950),
            .I(N__75925));
    Span4Mux_h I__17432 (
            .O(N__75947),
            .I(N__75925));
    LocalMux I__17431 (
            .O(N__75944),
            .I(N__75916));
    LocalMux I__17430 (
            .O(N__75939),
            .I(N__75916));
    Span4Mux_v I__17429 (
            .O(N__75936),
            .I(N__75916));
    Span4Mux_v I__17428 (
            .O(N__75933),
            .I(N__75916));
    Odrv4 I__17427 (
            .O(N__75930),
            .I(xy_ki_0_rep1));
    Odrv4 I__17426 (
            .O(N__75925),
            .I(xy_ki_0_rep1));
    Odrv4 I__17425 (
            .O(N__75916),
            .I(xy_ki_0_rep1));
    InMux I__17424 (
            .O(N__75909),
            .I(N__75905));
    CascadeMux I__17423 (
            .O(N__75908),
            .I(N__75901));
    LocalMux I__17422 (
            .O(N__75905),
            .I(N__75897));
    InMux I__17421 (
            .O(N__75904),
            .I(N__75893));
    InMux I__17420 (
            .O(N__75901),
            .I(N__75887));
    InMux I__17419 (
            .O(N__75900),
            .I(N__75887));
    Span4Mux_s3_h I__17418 (
            .O(N__75897),
            .I(N__75884));
    CascadeMux I__17417 (
            .O(N__75896),
            .I(N__75880));
    LocalMux I__17416 (
            .O(N__75893),
            .I(N__75876));
    InMux I__17415 (
            .O(N__75892),
            .I(N__75873));
    LocalMux I__17414 (
            .O(N__75887),
            .I(N__75870));
    Span4Mux_v I__17413 (
            .O(N__75884),
            .I(N__75867));
    InMux I__17412 (
            .O(N__75883),
            .I(N__75864));
    InMux I__17411 (
            .O(N__75880),
            .I(N__75859));
    InMux I__17410 (
            .O(N__75879),
            .I(N__75859));
    Span4Mux_h I__17409 (
            .O(N__75876),
            .I(N__75856));
    LocalMux I__17408 (
            .O(N__75873),
            .I(N__75853));
    Span4Mux_h I__17407 (
            .O(N__75870),
            .I(N__75850));
    Span4Mux_h I__17406 (
            .O(N__75867),
            .I(N__75843));
    LocalMux I__17405 (
            .O(N__75864),
            .I(N__75843));
    LocalMux I__17404 (
            .O(N__75859),
            .I(N__75843));
    Span4Mux_v I__17403 (
            .O(N__75856),
            .I(N__75840));
    Odrv12 I__17402 (
            .O(N__75853),
            .I(\pid_side.error_6 ));
    Odrv4 I__17401 (
            .O(N__75850),
            .I(\pid_side.error_6 ));
    Odrv4 I__17400 (
            .O(N__75843),
            .I(\pid_side.error_6 ));
    Odrv4 I__17399 (
            .O(N__75840),
            .I(\pid_side.error_6 ));
    InMux I__17398 (
            .O(N__75831),
            .I(N__75825));
    InMux I__17397 (
            .O(N__75830),
            .I(N__75818));
    InMux I__17396 (
            .O(N__75829),
            .I(N__75813));
    InMux I__17395 (
            .O(N__75828),
            .I(N__75813));
    LocalMux I__17394 (
            .O(N__75825),
            .I(N__75808));
    InMux I__17393 (
            .O(N__75824),
            .I(N__75805));
    InMux I__17392 (
            .O(N__75823),
            .I(N__75802));
    InMux I__17391 (
            .O(N__75822),
            .I(N__75797));
    InMux I__17390 (
            .O(N__75821),
            .I(N__75797));
    LocalMux I__17389 (
            .O(N__75818),
            .I(N__75794));
    LocalMux I__17388 (
            .O(N__75813),
            .I(N__75791));
    InMux I__17387 (
            .O(N__75812),
            .I(N__75786));
    InMux I__17386 (
            .O(N__75811),
            .I(N__75786));
    Span12Mux_s7_h I__17385 (
            .O(N__75808),
            .I(N__75783));
    LocalMux I__17384 (
            .O(N__75805),
            .I(N__75780));
    LocalMux I__17383 (
            .O(N__75802),
            .I(N__75775));
    LocalMux I__17382 (
            .O(N__75797),
            .I(N__75775));
    Span4Mux_v I__17381 (
            .O(N__75794),
            .I(N__75768));
    Span4Mux_v I__17380 (
            .O(N__75791),
            .I(N__75768));
    LocalMux I__17379 (
            .O(N__75786),
            .I(N__75768));
    Odrv12 I__17378 (
            .O(N__75783),
            .I(\pid_side.error_7 ));
    Odrv12 I__17377 (
            .O(N__75780),
            .I(\pid_side.error_7 ));
    Odrv4 I__17376 (
            .O(N__75775),
            .I(\pid_side.error_7 ));
    Odrv4 I__17375 (
            .O(N__75768),
            .I(\pid_side.error_7 ));
    InMux I__17374 (
            .O(N__75759),
            .I(N__75756));
    LocalMux I__17373 (
            .O(N__75756),
            .I(\pid_side.g0_7_1 ));
    InMux I__17372 (
            .O(N__75753),
            .I(N__75745));
    CascadeMux I__17371 (
            .O(N__75752),
            .I(N__75735));
    CascadeMux I__17370 (
            .O(N__75751),
            .I(N__75729));
    CascadeMux I__17369 (
            .O(N__75750),
            .I(N__75726));
    InMux I__17368 (
            .O(N__75749),
            .I(N__75722));
    InMux I__17367 (
            .O(N__75748),
            .I(N__75719));
    LocalMux I__17366 (
            .O(N__75745),
            .I(N__75714));
    InMux I__17365 (
            .O(N__75744),
            .I(N__75709));
    InMux I__17364 (
            .O(N__75743),
            .I(N__75709));
    InMux I__17363 (
            .O(N__75742),
            .I(N__75706));
    CascadeMux I__17362 (
            .O(N__75741),
            .I(N__75698));
    InMux I__17361 (
            .O(N__75740),
            .I(N__75694));
    CascadeMux I__17360 (
            .O(N__75739),
            .I(N__75691));
    InMux I__17359 (
            .O(N__75738),
            .I(N__75687));
    InMux I__17358 (
            .O(N__75735),
            .I(N__75682));
    InMux I__17357 (
            .O(N__75734),
            .I(N__75682));
    InMux I__17356 (
            .O(N__75733),
            .I(N__75677));
    InMux I__17355 (
            .O(N__75732),
            .I(N__75677));
    InMux I__17354 (
            .O(N__75729),
            .I(N__75670));
    InMux I__17353 (
            .O(N__75726),
            .I(N__75670));
    InMux I__17352 (
            .O(N__75725),
            .I(N__75670));
    LocalMux I__17351 (
            .O(N__75722),
            .I(N__75664));
    LocalMux I__17350 (
            .O(N__75719),
            .I(N__75664));
    InMux I__17349 (
            .O(N__75718),
            .I(N__75659));
    InMux I__17348 (
            .O(N__75717),
            .I(N__75659));
    Span4Mux_v I__17347 (
            .O(N__75714),
            .I(N__75656));
    LocalMux I__17346 (
            .O(N__75709),
            .I(N__75653));
    LocalMux I__17345 (
            .O(N__75706),
            .I(N__75650));
    InMux I__17344 (
            .O(N__75705),
            .I(N__75645));
    InMux I__17343 (
            .O(N__75704),
            .I(N__75645));
    InMux I__17342 (
            .O(N__75703),
            .I(N__75642));
    InMux I__17341 (
            .O(N__75702),
            .I(N__75639));
    InMux I__17340 (
            .O(N__75701),
            .I(N__75636));
    InMux I__17339 (
            .O(N__75698),
            .I(N__75631));
    InMux I__17338 (
            .O(N__75697),
            .I(N__75631));
    LocalMux I__17337 (
            .O(N__75694),
            .I(N__75628));
    InMux I__17336 (
            .O(N__75691),
            .I(N__75623));
    InMux I__17335 (
            .O(N__75690),
            .I(N__75623));
    LocalMux I__17334 (
            .O(N__75687),
            .I(N__75620));
    LocalMux I__17333 (
            .O(N__75682),
            .I(N__75613));
    LocalMux I__17332 (
            .O(N__75677),
            .I(N__75613));
    LocalMux I__17331 (
            .O(N__75670),
            .I(N__75613));
    InMux I__17330 (
            .O(N__75669),
            .I(N__75610));
    Span4Mux_v I__17329 (
            .O(N__75664),
            .I(N__75607));
    LocalMux I__17328 (
            .O(N__75659),
            .I(N__75604));
    Span4Mux_v I__17327 (
            .O(N__75656),
            .I(N__75597));
    Span4Mux_v I__17326 (
            .O(N__75653),
            .I(N__75597));
    Span4Mux_h I__17325 (
            .O(N__75650),
            .I(N__75597));
    LocalMux I__17324 (
            .O(N__75645),
            .I(N__75594));
    LocalMux I__17323 (
            .O(N__75642),
            .I(N__75585));
    LocalMux I__17322 (
            .O(N__75639),
            .I(N__75585));
    LocalMux I__17321 (
            .O(N__75636),
            .I(N__75585));
    LocalMux I__17320 (
            .O(N__75631),
            .I(N__75585));
    Span4Mux_v I__17319 (
            .O(N__75628),
            .I(N__75580));
    LocalMux I__17318 (
            .O(N__75623),
            .I(N__75580));
    Sp12to4 I__17317 (
            .O(N__75620),
            .I(N__75573));
    Sp12to4 I__17316 (
            .O(N__75613),
            .I(N__75573));
    LocalMux I__17315 (
            .O(N__75610),
            .I(N__75573));
    Span4Mux_h I__17314 (
            .O(N__75607),
            .I(N__75568));
    Span4Mux_v I__17313 (
            .O(N__75604),
            .I(N__75568));
    Span4Mux_h I__17312 (
            .O(N__75597),
            .I(N__75565));
    Span4Mux_v I__17311 (
            .O(N__75594),
            .I(N__75558));
    Span4Mux_v I__17310 (
            .O(N__75585),
            .I(N__75558));
    Span4Mux_h I__17309 (
            .O(N__75580),
            .I(N__75558));
    Span12Mux_v I__17308 (
            .O(N__75573),
            .I(N__75555));
    Odrv4 I__17307 (
            .O(N__75568),
            .I(xy_ki_3));
    Odrv4 I__17306 (
            .O(N__75565),
            .I(xy_ki_3));
    Odrv4 I__17305 (
            .O(N__75558),
            .I(xy_ki_3));
    Odrv12 I__17304 (
            .O(N__75555),
            .I(xy_ki_3));
    InMux I__17303 (
            .O(N__75546),
            .I(N__75543));
    LocalMux I__17302 (
            .O(N__75543),
            .I(N__75540));
    Odrv4 I__17301 (
            .O(N__75540),
            .I(\pid_side.N_117 ));
    CascadeMux I__17300 (
            .O(N__75537),
            .I(N__75529));
    CascadeMux I__17299 (
            .O(N__75536),
            .I(N__75525));
    CascadeMux I__17298 (
            .O(N__75535),
            .I(N__75522));
    CascadeMux I__17297 (
            .O(N__75534),
            .I(N__75519));
    CascadeMux I__17296 (
            .O(N__75533),
            .I(N__75515));
    InMux I__17295 (
            .O(N__75532),
            .I(N__75512));
    InMux I__17294 (
            .O(N__75529),
            .I(N__75509));
    CascadeMux I__17293 (
            .O(N__75528),
            .I(N__75505));
    InMux I__17292 (
            .O(N__75525),
            .I(N__75500));
    InMux I__17291 (
            .O(N__75522),
            .I(N__75500));
    InMux I__17290 (
            .O(N__75519),
            .I(N__75495));
    InMux I__17289 (
            .O(N__75518),
            .I(N__75495));
    InMux I__17288 (
            .O(N__75515),
            .I(N__75492));
    LocalMux I__17287 (
            .O(N__75512),
            .I(N__75489));
    LocalMux I__17286 (
            .O(N__75509),
            .I(N__75485));
    InMux I__17285 (
            .O(N__75508),
            .I(N__75482));
    InMux I__17284 (
            .O(N__75505),
            .I(N__75478));
    LocalMux I__17283 (
            .O(N__75500),
            .I(N__75465));
    LocalMux I__17282 (
            .O(N__75495),
            .I(N__75465));
    LocalMux I__17281 (
            .O(N__75492),
            .I(N__75465));
    Span4Mux_h I__17280 (
            .O(N__75489),
            .I(N__75465));
    InMux I__17279 (
            .O(N__75488),
            .I(N__75462));
    Span4Mux_h I__17278 (
            .O(N__75485),
            .I(N__75459));
    LocalMux I__17277 (
            .O(N__75482),
            .I(N__75456));
    CascadeMux I__17276 (
            .O(N__75481),
            .I(N__75453));
    LocalMux I__17275 (
            .O(N__75478),
            .I(N__75450));
    InMux I__17274 (
            .O(N__75477),
            .I(N__75445));
    InMux I__17273 (
            .O(N__75476),
            .I(N__75445));
    InMux I__17272 (
            .O(N__75475),
            .I(N__75442));
    InMux I__17271 (
            .O(N__75474),
            .I(N__75439));
    Span4Mux_v I__17270 (
            .O(N__75465),
            .I(N__75434));
    LocalMux I__17269 (
            .O(N__75462),
            .I(N__75434));
    Span4Mux_v I__17268 (
            .O(N__75459),
            .I(N__75429));
    Span4Mux_v I__17267 (
            .O(N__75456),
            .I(N__75429));
    InMux I__17266 (
            .O(N__75453),
            .I(N__75426));
    Span4Mux_v I__17265 (
            .O(N__75450),
            .I(N__75423));
    LocalMux I__17264 (
            .O(N__75445),
            .I(N__75420));
    LocalMux I__17263 (
            .O(N__75442),
            .I(N__75417));
    LocalMux I__17262 (
            .O(N__75439),
            .I(N__75410));
    Span4Mux_v I__17261 (
            .O(N__75434),
            .I(N__75410));
    Span4Mux_h I__17260 (
            .O(N__75429),
            .I(N__75410));
    LocalMux I__17259 (
            .O(N__75426),
            .I(N__75403));
    Span4Mux_h I__17258 (
            .O(N__75423),
            .I(N__75403));
    Span4Mux_v I__17257 (
            .O(N__75420),
            .I(N__75403));
    Span4Mux_h I__17256 (
            .O(N__75417),
            .I(N__75400));
    Span4Mux_h I__17255 (
            .O(N__75410),
            .I(N__75397));
    Odrv4 I__17254 (
            .O(N__75403),
            .I(pid_side_N_166));
    Odrv4 I__17253 (
            .O(N__75400),
            .I(pid_side_N_166));
    Odrv4 I__17252 (
            .O(N__75397),
            .I(pid_side_N_166));
    CascadeMux I__17251 (
            .O(N__75390),
            .I(N__75387));
    InMux I__17250 (
            .O(N__75387),
            .I(N__75384));
    LocalMux I__17249 (
            .O(N__75384),
            .I(N__75381));
    Span4Mux_h I__17248 (
            .O(N__75381),
            .I(N__75378));
    Span4Mux_v I__17247 (
            .O(N__75378),
            .I(N__75375));
    Odrv4 I__17246 (
            .O(N__75375),
            .I(\pid_side.error_i_regZ0Z_5 ));
    CEMux I__17245 (
            .O(N__75372),
            .I(N__75369));
    LocalMux I__17244 (
            .O(N__75369),
            .I(N__75363));
    CEMux I__17243 (
            .O(N__75368),
            .I(N__75360));
    CEMux I__17242 (
            .O(N__75367),
            .I(N__75357));
    CEMux I__17241 (
            .O(N__75366),
            .I(N__75353));
    Span4Mux_h I__17240 (
            .O(N__75363),
            .I(N__75348));
    LocalMux I__17239 (
            .O(N__75360),
            .I(N__75348));
    LocalMux I__17238 (
            .O(N__75357),
            .I(N__75345));
    CEMux I__17237 (
            .O(N__75356),
            .I(N__75341));
    LocalMux I__17236 (
            .O(N__75353),
            .I(N__75338));
    Span4Mux_v I__17235 (
            .O(N__75348),
            .I(N__75333));
    Span4Mux_v I__17234 (
            .O(N__75345),
            .I(N__75333));
    CEMux I__17233 (
            .O(N__75344),
            .I(N__75326));
    LocalMux I__17232 (
            .O(N__75341),
            .I(N__75323));
    Span4Mux_h I__17231 (
            .O(N__75338),
            .I(N__75318));
    Span4Mux_h I__17230 (
            .O(N__75333),
            .I(N__75318));
    CEMux I__17229 (
            .O(N__75332),
            .I(N__75315));
    CEMux I__17228 (
            .O(N__75331),
            .I(N__75312));
    CEMux I__17227 (
            .O(N__75330),
            .I(N__75309));
    CEMux I__17226 (
            .O(N__75329),
            .I(N__75306));
    LocalMux I__17225 (
            .O(N__75326),
            .I(N__75302));
    Span4Mux_v I__17224 (
            .O(N__75323),
            .I(N__75294));
    Span4Mux_h I__17223 (
            .O(N__75318),
            .I(N__75294));
    LocalMux I__17222 (
            .O(N__75315),
            .I(N__75294));
    LocalMux I__17221 (
            .O(N__75312),
            .I(N__75291));
    LocalMux I__17220 (
            .O(N__75309),
            .I(N__75284));
    LocalMux I__17219 (
            .O(N__75306),
            .I(N__75284));
    CEMux I__17218 (
            .O(N__75305),
            .I(N__75281));
    Span4Mux_h I__17217 (
            .O(N__75302),
            .I(N__75278));
    CEMux I__17216 (
            .O(N__75301),
            .I(N__75275));
    Span4Mux_h I__17215 (
            .O(N__75294),
            .I(N__75272));
    Span4Mux_v I__17214 (
            .O(N__75291),
            .I(N__75269));
    CEMux I__17213 (
            .O(N__75290),
            .I(N__75266));
    CEMux I__17212 (
            .O(N__75289),
            .I(N__75263));
    Span4Mux_v I__17211 (
            .O(N__75284),
            .I(N__75260));
    LocalMux I__17210 (
            .O(N__75281),
            .I(N__75255));
    Span4Mux_v I__17209 (
            .O(N__75278),
            .I(N__75255));
    LocalMux I__17208 (
            .O(N__75275),
            .I(N__75250));
    Span4Mux_v I__17207 (
            .O(N__75272),
            .I(N__75250));
    Span4Mux_v I__17206 (
            .O(N__75269),
            .I(N__75247));
    LocalMux I__17205 (
            .O(N__75266),
            .I(N__75240));
    LocalMux I__17204 (
            .O(N__75263),
            .I(N__75240));
    Span4Mux_h I__17203 (
            .O(N__75260),
            .I(N__75240));
    Sp12to4 I__17202 (
            .O(N__75255),
            .I(N__75237));
    Span4Mux_v I__17201 (
            .O(N__75250),
            .I(N__75234));
    Odrv4 I__17200 (
            .O(N__75247),
            .I(\pid_side.state_ns_0_0 ));
    Odrv4 I__17199 (
            .O(N__75240),
            .I(\pid_side.state_ns_0_0 ));
    Odrv12 I__17198 (
            .O(N__75237),
            .I(\pid_side.state_ns_0_0 ));
    Odrv4 I__17197 (
            .O(N__75234),
            .I(\pid_side.state_ns_0_0 ));
    CascadeMux I__17196 (
            .O(N__75225),
            .I(\pid_side.g0_6_1_cascade_ ));
    InMux I__17195 (
            .O(N__75222),
            .I(N__75219));
    LocalMux I__17194 (
            .O(N__75219),
            .I(\pid_side.N_12_1_1 ));
    CascadeMux I__17193 (
            .O(N__75216),
            .I(\pid_side.N_12_1_1_cascade_ ));
    InMux I__17192 (
            .O(N__75213),
            .I(N__75210));
    LocalMux I__17191 (
            .O(N__75210),
            .I(\pid_side.N_89_0_1 ));
    InMux I__17190 (
            .O(N__75207),
            .I(N__75204));
    LocalMux I__17189 (
            .O(N__75204),
            .I(\pid_side.N_116_0 ));
    InMux I__17188 (
            .O(N__75201),
            .I(N__75198));
    LocalMux I__17187 (
            .O(N__75198),
            .I(N__75194));
    InMux I__17186 (
            .O(N__75197),
            .I(N__75189));
    Span4Mux_s3_h I__17185 (
            .O(N__75194),
            .I(N__75186));
    InMux I__17184 (
            .O(N__75193),
            .I(N__75181));
    InMux I__17183 (
            .O(N__75192),
            .I(N__75178));
    LocalMux I__17182 (
            .O(N__75189),
            .I(N__75175));
    Span4Mux_v I__17181 (
            .O(N__75186),
            .I(N__75172));
    InMux I__17180 (
            .O(N__75185),
            .I(N__75167));
    InMux I__17179 (
            .O(N__75184),
            .I(N__75167));
    LocalMux I__17178 (
            .O(N__75181),
            .I(N__75164));
    LocalMux I__17177 (
            .O(N__75178),
            .I(N__75161));
    Span4Mux_s3_h I__17176 (
            .O(N__75175),
            .I(N__75158));
    Span4Mux_h I__17175 (
            .O(N__75172),
            .I(N__75153));
    LocalMux I__17174 (
            .O(N__75167),
            .I(N__75153));
    Span4Mux_h I__17173 (
            .O(N__75164),
            .I(N__75150));
    Span4Mux_v I__17172 (
            .O(N__75161),
            .I(N__75147));
    Odrv4 I__17171 (
            .O(N__75158),
            .I(\pid_side.error_3 ));
    Odrv4 I__17170 (
            .O(N__75153),
            .I(\pid_side.error_3 ));
    Odrv4 I__17169 (
            .O(N__75150),
            .I(\pid_side.error_3 ));
    Odrv4 I__17168 (
            .O(N__75147),
            .I(\pid_side.error_3 ));
    InMux I__17167 (
            .O(N__75138),
            .I(N__75135));
    LocalMux I__17166 (
            .O(N__75135),
            .I(N__75131));
    InMux I__17165 (
            .O(N__75134),
            .I(N__75125));
    Span4Mux_s3_h I__17164 (
            .O(N__75131),
            .I(N__75122));
    CascadeMux I__17163 (
            .O(N__75130),
            .I(N__75119));
    InMux I__17162 (
            .O(N__75129),
            .I(N__75113));
    InMux I__17161 (
            .O(N__75128),
            .I(N__75113));
    LocalMux I__17160 (
            .O(N__75125),
            .I(N__75110));
    Span4Mux_v I__17159 (
            .O(N__75122),
            .I(N__75107));
    InMux I__17158 (
            .O(N__75119),
            .I(N__75102));
    InMux I__17157 (
            .O(N__75118),
            .I(N__75102));
    LocalMux I__17156 (
            .O(N__75113),
            .I(N__75099));
    Span4Mux_s3_h I__17155 (
            .O(N__75110),
            .I(N__75096));
    Span4Mux_h I__17154 (
            .O(N__75107),
            .I(N__75091));
    LocalMux I__17153 (
            .O(N__75102),
            .I(N__75091));
    Span4Mux_v I__17152 (
            .O(N__75099),
            .I(N__75088));
    Odrv4 I__17151 (
            .O(N__75096),
            .I(\pid_side.error_2 ));
    Odrv4 I__17150 (
            .O(N__75091),
            .I(\pid_side.error_2 ));
    Odrv4 I__17149 (
            .O(N__75088),
            .I(\pid_side.error_2 ));
    InMux I__17148 (
            .O(N__75081),
            .I(N__75078));
    LocalMux I__17147 (
            .O(N__75078),
            .I(N__75075));
    Span4Mux_s3_h I__17146 (
            .O(N__75075),
            .I(N__75070));
    InMux I__17145 (
            .O(N__75074),
            .I(N__75065));
    InMux I__17144 (
            .O(N__75073),
            .I(N__75062));
    Span4Mux_v I__17143 (
            .O(N__75070),
            .I(N__75059));
    InMux I__17142 (
            .O(N__75069),
            .I(N__75054));
    InMux I__17141 (
            .O(N__75068),
            .I(N__75054));
    LocalMux I__17140 (
            .O(N__75065),
            .I(N__75051));
    LocalMux I__17139 (
            .O(N__75062),
            .I(N__75047));
    Span4Mux_h I__17138 (
            .O(N__75059),
            .I(N__75042));
    LocalMux I__17137 (
            .O(N__75054),
            .I(N__75042));
    Span4Mux_h I__17136 (
            .O(N__75051),
            .I(N__75039));
    InMux I__17135 (
            .O(N__75050),
            .I(N__75036));
    Odrv12 I__17134 (
            .O(N__75047),
            .I(\pid_side.error_5 ));
    Odrv4 I__17133 (
            .O(N__75042),
            .I(\pid_side.error_5 ));
    Odrv4 I__17132 (
            .O(N__75039),
            .I(\pid_side.error_5 ));
    LocalMux I__17131 (
            .O(N__75036),
            .I(\pid_side.error_5 ));
    InMux I__17130 (
            .O(N__75027),
            .I(N__75024));
    LocalMux I__17129 (
            .O(N__75024),
            .I(N__75020));
    InMux I__17128 (
            .O(N__75023),
            .I(N__75017));
    Span4Mux_s2_h I__17127 (
            .O(N__75020),
            .I(N__75011));
    LocalMux I__17126 (
            .O(N__75017),
            .I(N__75008));
    InMux I__17125 (
            .O(N__75016),
            .I(N__75004));
    InMux I__17124 (
            .O(N__75015),
            .I(N__75001));
    InMux I__17123 (
            .O(N__75014),
            .I(N__74998));
    Span4Mux_h I__17122 (
            .O(N__75011),
            .I(N__74995));
    Span4Mux_h I__17121 (
            .O(N__75008),
            .I(N__74992));
    InMux I__17120 (
            .O(N__75007),
            .I(N__74989));
    LocalMux I__17119 (
            .O(N__75004),
            .I(N__74986));
    LocalMux I__17118 (
            .O(N__75001),
            .I(N__74981));
    LocalMux I__17117 (
            .O(N__74998),
            .I(N__74981));
    Span4Mux_v I__17116 (
            .O(N__74995),
            .I(N__74978));
    Odrv4 I__17115 (
            .O(N__74992),
            .I(\pid_side.error_4 ));
    LocalMux I__17114 (
            .O(N__74989),
            .I(\pid_side.error_4 ));
    Odrv12 I__17113 (
            .O(N__74986),
            .I(\pid_side.error_4 ));
    Odrv4 I__17112 (
            .O(N__74981),
            .I(\pid_side.error_4 ));
    Odrv4 I__17111 (
            .O(N__74978),
            .I(\pid_side.error_4 ));
    CascadeMux I__17110 (
            .O(N__74967),
            .I(\pid_side.g0_10_1_cascade_ ));
    InMux I__17109 (
            .O(N__74964),
            .I(N__74961));
    LocalMux I__17108 (
            .O(N__74961),
            .I(\pid_side.N_12_1_0 ));
    InMux I__17107 (
            .O(N__74958),
            .I(N__74955));
    LocalMux I__17106 (
            .O(N__74955),
            .I(N__74952));
    Odrv12 I__17105 (
            .O(N__74952),
            .I(drone_H_disp_side_15));
    CascadeMux I__17104 (
            .O(N__74949),
            .I(N__74945));
    InMux I__17103 (
            .O(N__74948),
            .I(N__74940));
    InMux I__17102 (
            .O(N__74945),
            .I(N__74940));
    LocalMux I__17101 (
            .O(N__74940),
            .I(N__74937));
    Odrv12 I__17100 (
            .O(N__74937),
            .I(drone_H_disp_side_14));
    InMux I__17099 (
            .O(N__74934),
            .I(\pid_side.error_cry_10 ));
    InMux I__17098 (
            .O(N__74931),
            .I(N__74918));
    InMux I__17097 (
            .O(N__74930),
            .I(N__74915));
    InMux I__17096 (
            .O(N__74929),
            .I(N__74912));
    InMux I__17095 (
            .O(N__74928),
            .I(N__74907));
    InMux I__17094 (
            .O(N__74927),
            .I(N__74907));
    InMux I__17093 (
            .O(N__74926),
            .I(N__74901));
    InMux I__17092 (
            .O(N__74925),
            .I(N__74896));
    InMux I__17091 (
            .O(N__74924),
            .I(N__74896));
    InMux I__17090 (
            .O(N__74923),
            .I(N__74889));
    InMux I__17089 (
            .O(N__74922),
            .I(N__74889));
    InMux I__17088 (
            .O(N__74921),
            .I(N__74889));
    LocalMux I__17087 (
            .O(N__74918),
            .I(N__74886));
    LocalMux I__17086 (
            .O(N__74915),
            .I(N__74880));
    LocalMux I__17085 (
            .O(N__74912),
            .I(N__74875));
    LocalMux I__17084 (
            .O(N__74907),
            .I(N__74875));
    InMux I__17083 (
            .O(N__74906),
            .I(N__74872));
    InMux I__17082 (
            .O(N__74905),
            .I(N__74869));
    InMux I__17081 (
            .O(N__74904),
            .I(N__74865));
    LocalMux I__17080 (
            .O(N__74901),
            .I(N__74858));
    LocalMux I__17079 (
            .O(N__74896),
            .I(N__74858));
    LocalMux I__17078 (
            .O(N__74889),
            .I(N__74858));
    Span4Mux_s3_h I__17077 (
            .O(N__74886),
            .I(N__74855));
    InMux I__17076 (
            .O(N__74885),
            .I(N__74848));
    InMux I__17075 (
            .O(N__74884),
            .I(N__74848));
    InMux I__17074 (
            .O(N__74883),
            .I(N__74848));
    Span4Mux_s2_h I__17073 (
            .O(N__74880),
            .I(N__74845));
    Span4Mux_h I__17072 (
            .O(N__74875),
            .I(N__74838));
    LocalMux I__17071 (
            .O(N__74872),
            .I(N__74835));
    LocalMux I__17070 (
            .O(N__74869),
            .I(N__74832));
    InMux I__17069 (
            .O(N__74868),
            .I(N__74829));
    LocalMux I__17068 (
            .O(N__74865),
            .I(N__74826));
    Span4Mux_v I__17067 (
            .O(N__74858),
            .I(N__74823));
    Span4Mux_v I__17066 (
            .O(N__74855),
            .I(N__74820));
    LocalMux I__17065 (
            .O(N__74848),
            .I(N__74817));
    Span4Mux_h I__17064 (
            .O(N__74845),
            .I(N__74814));
    InMux I__17063 (
            .O(N__74844),
            .I(N__74811));
    InMux I__17062 (
            .O(N__74843),
            .I(N__74804));
    InMux I__17061 (
            .O(N__74842),
            .I(N__74804));
    InMux I__17060 (
            .O(N__74841),
            .I(N__74804));
    Span4Mux_v I__17059 (
            .O(N__74838),
            .I(N__74795));
    Span4Mux_v I__17058 (
            .O(N__74835),
            .I(N__74795));
    Span4Mux_h I__17057 (
            .O(N__74832),
            .I(N__74795));
    LocalMux I__17056 (
            .O(N__74829),
            .I(N__74795));
    Span4Mux_h I__17055 (
            .O(N__74826),
            .I(N__74792));
    Span4Mux_h I__17054 (
            .O(N__74823),
            .I(N__74785));
    Span4Mux_h I__17053 (
            .O(N__74820),
            .I(N__74785));
    Span4Mux_h I__17052 (
            .O(N__74817),
            .I(N__74785));
    Odrv4 I__17051 (
            .O(N__74814),
            .I(\pid_side.error_15 ));
    LocalMux I__17050 (
            .O(N__74811),
            .I(\pid_side.error_15 ));
    LocalMux I__17049 (
            .O(N__74804),
            .I(\pid_side.error_15 ));
    Odrv4 I__17048 (
            .O(N__74795),
            .I(\pid_side.error_15 ));
    Odrv4 I__17047 (
            .O(N__74792),
            .I(\pid_side.error_15 ));
    Odrv4 I__17046 (
            .O(N__74785),
            .I(\pid_side.error_15 ));
    InMux I__17045 (
            .O(N__74772),
            .I(N__74769));
    LocalMux I__17044 (
            .O(N__74769),
            .I(N__74764));
    InMux I__17043 (
            .O(N__74768),
            .I(N__74761));
    InMux I__17042 (
            .O(N__74767),
            .I(N__74758));
    Span4Mux_v I__17041 (
            .O(N__74764),
            .I(N__74751));
    LocalMux I__17040 (
            .O(N__74761),
            .I(N__74751));
    LocalMux I__17039 (
            .O(N__74758),
            .I(N__74747));
    InMux I__17038 (
            .O(N__74757),
            .I(N__74742));
    InMux I__17037 (
            .O(N__74756),
            .I(N__74742));
    Span4Mux_v I__17036 (
            .O(N__74751),
            .I(N__74739));
    InMux I__17035 (
            .O(N__74750),
            .I(N__74736));
    Span4Mux_h I__17034 (
            .O(N__74747),
            .I(N__74729));
    LocalMux I__17033 (
            .O(N__74742),
            .I(N__74729));
    Span4Mux_h I__17032 (
            .O(N__74739),
            .I(N__74726));
    LocalMux I__17031 (
            .O(N__74736),
            .I(N__74723));
    InMux I__17030 (
            .O(N__74735),
            .I(N__74720));
    InMux I__17029 (
            .O(N__74734),
            .I(N__74717));
    Span4Mux_v I__17028 (
            .O(N__74729),
            .I(N__74714));
    Odrv4 I__17027 (
            .O(N__74726),
            .I(\pid_side.error_8 ));
    Odrv4 I__17026 (
            .O(N__74723),
            .I(\pid_side.error_8 ));
    LocalMux I__17025 (
            .O(N__74720),
            .I(\pid_side.error_8 ));
    LocalMux I__17024 (
            .O(N__74717),
            .I(\pid_side.error_8 ));
    Odrv4 I__17023 (
            .O(N__74714),
            .I(\pid_side.error_8 ));
    CascadeMux I__17022 (
            .O(N__74703),
            .I(\pid_side.N_48_1_0_cascade_ ));
    InMux I__17021 (
            .O(N__74700),
            .I(N__74694));
    InMux I__17020 (
            .O(N__74699),
            .I(N__74694));
    LocalMux I__17019 (
            .O(N__74694),
            .I(\pid_side.N_51_1_0 ));
    InMux I__17018 (
            .O(N__74691),
            .I(N__74688));
    LocalMux I__17017 (
            .O(N__74688),
            .I(\pid_side.N_48_1_0 ));
    CascadeMux I__17016 (
            .O(N__74685),
            .I(\pid_side.error_i_reg_esr_RNO_9Z0Z_21_cascade_ ));
    InMux I__17015 (
            .O(N__74682),
            .I(N__74679));
    LocalMux I__17014 (
            .O(N__74679),
            .I(\pid_side.error_i_reg_esr_RNO_10Z0Z_21 ));
    InMux I__17013 (
            .O(N__74676),
            .I(N__74673));
    LocalMux I__17012 (
            .O(N__74673),
            .I(N__74670));
    Span4Mux_v I__17011 (
            .O(N__74670),
            .I(N__74667));
    Odrv4 I__17010 (
            .O(N__74667),
            .I(\pid_side.N_116_0_0 ));
    InMux I__17009 (
            .O(N__74664),
            .I(N__74661));
    LocalMux I__17008 (
            .O(N__74661),
            .I(\pid_side.N_51_1 ));
    InMux I__17007 (
            .O(N__74658),
            .I(N__74652));
    InMux I__17006 (
            .O(N__74657),
            .I(N__74649));
    InMux I__17005 (
            .O(N__74656),
            .I(N__74646));
    InMux I__17004 (
            .O(N__74655),
            .I(N__74643));
    LocalMux I__17003 (
            .O(N__74652),
            .I(N__74637));
    LocalMux I__17002 (
            .O(N__74649),
            .I(N__74637));
    LocalMux I__17001 (
            .O(N__74646),
            .I(N__74634));
    LocalMux I__17000 (
            .O(N__74643),
            .I(N__74631));
    CascadeMux I__16999 (
            .O(N__74642),
            .I(N__74625));
    Span12Mux_v I__16998 (
            .O(N__74637),
            .I(N__74621));
    Span4Mux_v I__16997 (
            .O(N__74634),
            .I(N__74616));
    Span4Mux_h I__16996 (
            .O(N__74631),
            .I(N__74616));
    InMux I__16995 (
            .O(N__74630),
            .I(N__74613));
    InMux I__16994 (
            .O(N__74629),
            .I(N__74608));
    InMux I__16993 (
            .O(N__74628),
            .I(N__74608));
    InMux I__16992 (
            .O(N__74625),
            .I(N__74603));
    InMux I__16991 (
            .O(N__74624),
            .I(N__74603));
    Odrv12 I__16990 (
            .O(N__74621),
            .I(\pid_side.error_9 ));
    Odrv4 I__16989 (
            .O(N__74616),
            .I(\pid_side.error_9 ));
    LocalMux I__16988 (
            .O(N__74613),
            .I(\pid_side.error_9 ));
    LocalMux I__16987 (
            .O(N__74608),
            .I(\pid_side.error_9 ));
    LocalMux I__16986 (
            .O(N__74603),
            .I(\pid_side.error_9 ));
    InMux I__16985 (
            .O(N__74592),
            .I(N__74587));
    InMux I__16984 (
            .O(N__74591),
            .I(N__74584));
    InMux I__16983 (
            .O(N__74590),
            .I(N__74579));
    LocalMux I__16982 (
            .O(N__74587),
            .I(N__74576));
    LocalMux I__16981 (
            .O(N__74584),
            .I(N__74571));
    InMux I__16980 (
            .O(N__74583),
            .I(N__74566));
    InMux I__16979 (
            .O(N__74582),
            .I(N__74566));
    LocalMux I__16978 (
            .O(N__74579),
            .I(N__74561));
    Span4Mux_v I__16977 (
            .O(N__74576),
            .I(N__74561));
    CascadeMux I__16976 (
            .O(N__74575),
            .I(N__74558));
    InMux I__16975 (
            .O(N__74574),
            .I(N__74554));
    Span4Mux_h I__16974 (
            .O(N__74571),
            .I(N__74549));
    LocalMux I__16973 (
            .O(N__74566),
            .I(N__74549));
    Span4Mux_v I__16972 (
            .O(N__74561),
            .I(N__74544));
    InMux I__16971 (
            .O(N__74558),
            .I(N__74541));
    InMux I__16970 (
            .O(N__74557),
            .I(N__74538));
    LocalMux I__16969 (
            .O(N__74554),
            .I(N__74533));
    Span4Mux_v I__16968 (
            .O(N__74549),
            .I(N__74533));
    InMux I__16967 (
            .O(N__74548),
            .I(N__74528));
    InMux I__16966 (
            .O(N__74547),
            .I(N__74528));
    Span4Mux_h I__16965 (
            .O(N__74544),
            .I(N__74525));
    LocalMux I__16964 (
            .O(N__74541),
            .I(\pid_side.error_10 ));
    LocalMux I__16963 (
            .O(N__74538),
            .I(\pid_side.error_10 ));
    Odrv4 I__16962 (
            .O(N__74533),
            .I(\pid_side.error_10 ));
    LocalMux I__16961 (
            .O(N__74528),
            .I(\pid_side.error_10 ));
    Odrv4 I__16960 (
            .O(N__74525),
            .I(\pid_side.error_10 ));
    CascadeMux I__16959 (
            .O(N__74514),
            .I(N__74510));
    InMux I__16958 (
            .O(N__74513),
            .I(N__74506));
    InMux I__16957 (
            .O(N__74510),
            .I(N__74503));
    InMux I__16956 (
            .O(N__74509),
            .I(N__74499));
    LocalMux I__16955 (
            .O(N__74506),
            .I(N__74496));
    LocalMux I__16954 (
            .O(N__74503),
            .I(N__74493));
    InMux I__16953 (
            .O(N__74502),
            .I(N__74490));
    LocalMux I__16952 (
            .O(N__74499),
            .I(N__74486));
    Span4Mux_s2_h I__16951 (
            .O(N__74496),
            .I(N__74483));
    Span4Mux_h I__16950 (
            .O(N__74493),
            .I(N__74476));
    LocalMux I__16949 (
            .O(N__74490),
            .I(N__74473));
    InMux I__16948 (
            .O(N__74489),
            .I(N__74470));
    Span4Mux_s2_h I__16947 (
            .O(N__74486),
            .I(N__74467));
    Span4Mux_v I__16946 (
            .O(N__74483),
            .I(N__74464));
    InMux I__16945 (
            .O(N__74482),
            .I(N__74461));
    InMux I__16944 (
            .O(N__74481),
            .I(N__74458));
    InMux I__16943 (
            .O(N__74480),
            .I(N__74455));
    InMux I__16942 (
            .O(N__74479),
            .I(N__74452));
    Span4Mux_v I__16941 (
            .O(N__74476),
            .I(N__74445));
    Span4Mux_h I__16940 (
            .O(N__74473),
            .I(N__74445));
    LocalMux I__16939 (
            .O(N__74470),
            .I(N__74445));
    Span4Mux_h I__16938 (
            .O(N__74467),
            .I(N__74442));
    Span4Mux_h I__16937 (
            .O(N__74464),
            .I(N__74439));
    LocalMux I__16936 (
            .O(N__74461),
            .I(\pid_side.error_13 ));
    LocalMux I__16935 (
            .O(N__74458),
            .I(\pid_side.error_13 ));
    LocalMux I__16934 (
            .O(N__74455),
            .I(\pid_side.error_13 ));
    LocalMux I__16933 (
            .O(N__74452),
            .I(\pid_side.error_13 ));
    Odrv4 I__16932 (
            .O(N__74445),
            .I(\pid_side.error_13 ));
    Odrv4 I__16931 (
            .O(N__74442),
            .I(\pid_side.error_13 ));
    Odrv4 I__16930 (
            .O(N__74439),
            .I(\pid_side.error_13 ));
    CascadeMux I__16929 (
            .O(N__74424),
            .I(\pid_side.G_5_0_m4_1_cascade_ ));
    InMux I__16928 (
            .O(N__74421),
            .I(N__74413));
    InMux I__16927 (
            .O(N__74420),
            .I(N__74413));
    CascadeMux I__16926 (
            .O(N__74419),
            .I(N__74410));
    InMux I__16925 (
            .O(N__74418),
            .I(N__74405));
    LocalMux I__16924 (
            .O(N__74413),
            .I(N__74399));
    InMux I__16923 (
            .O(N__74410),
            .I(N__74394));
    InMux I__16922 (
            .O(N__74409),
            .I(N__74394));
    InMux I__16921 (
            .O(N__74408),
            .I(N__74391));
    LocalMux I__16920 (
            .O(N__74405),
            .I(N__74388));
    InMux I__16919 (
            .O(N__74404),
            .I(N__74384));
    InMux I__16918 (
            .O(N__74403),
            .I(N__74376));
    InMux I__16917 (
            .O(N__74402),
            .I(N__74376));
    Span4Mux_v I__16916 (
            .O(N__74399),
            .I(N__74371));
    LocalMux I__16915 (
            .O(N__74394),
            .I(N__74371));
    LocalMux I__16914 (
            .O(N__74391),
            .I(N__74368));
    Span4Mux_s2_h I__16913 (
            .O(N__74388),
            .I(N__74365));
    InMux I__16912 (
            .O(N__74387),
            .I(N__74362));
    LocalMux I__16911 (
            .O(N__74384),
            .I(N__74359));
    InMux I__16910 (
            .O(N__74383),
            .I(N__74356));
    InMux I__16909 (
            .O(N__74382),
            .I(N__74351));
    InMux I__16908 (
            .O(N__74381),
            .I(N__74351));
    LocalMux I__16907 (
            .O(N__74376),
            .I(N__74348));
    Span4Mux_h I__16906 (
            .O(N__74371),
            .I(N__74345));
    Span12Mux_s7_h I__16905 (
            .O(N__74368),
            .I(N__74342));
    Span4Mux_h I__16904 (
            .O(N__74365),
            .I(N__74339));
    LocalMux I__16903 (
            .O(N__74362),
            .I(\pid_side.error_14 ));
    Odrv4 I__16902 (
            .O(N__74359),
            .I(\pid_side.error_14 ));
    LocalMux I__16901 (
            .O(N__74356),
            .I(\pid_side.error_14 ));
    LocalMux I__16900 (
            .O(N__74351),
            .I(\pid_side.error_14 ));
    Odrv12 I__16899 (
            .O(N__74348),
            .I(\pid_side.error_14 ));
    Odrv4 I__16898 (
            .O(N__74345),
            .I(\pid_side.error_14 ));
    Odrv12 I__16897 (
            .O(N__74342),
            .I(\pid_side.error_14 ));
    Odrv4 I__16896 (
            .O(N__74339),
            .I(\pid_side.error_14 ));
    InMux I__16895 (
            .O(N__74322),
            .I(N__74319));
    LocalMux I__16894 (
            .O(N__74319),
            .I(N__74316));
    Span4Mux_h I__16893 (
            .O(N__74316),
            .I(N__74313));
    Odrv4 I__16892 (
            .O(N__74313),
            .I(\pid_side.N_7 ));
    InMux I__16891 (
            .O(N__74310),
            .I(N__74307));
    LocalMux I__16890 (
            .O(N__74307),
            .I(side_command_3));
    CascadeMux I__16889 (
            .O(N__74304),
            .I(N__74301));
    InMux I__16888 (
            .O(N__74301),
            .I(N__74298));
    LocalMux I__16887 (
            .O(N__74298),
            .I(N__74295));
    Odrv12 I__16886 (
            .O(N__74295),
            .I(drone_H_disp_side_i_7));
    InMux I__16885 (
            .O(N__74292),
            .I(\pid_side.error_cry_2_0 ));
    InMux I__16884 (
            .O(N__74289),
            .I(N__74286));
    LocalMux I__16883 (
            .O(N__74286),
            .I(N__74283));
    Span4Mux_h I__16882 (
            .O(N__74283),
            .I(N__74280));
    Span4Mux_h I__16881 (
            .O(N__74280),
            .I(N__74277));
    Odrv4 I__16880 (
            .O(N__74277),
            .I(drone_H_disp_side_i_8));
    CascadeMux I__16879 (
            .O(N__74274),
            .I(N__74271));
    InMux I__16878 (
            .O(N__74271),
            .I(N__74268));
    LocalMux I__16877 (
            .O(N__74268),
            .I(N__74265));
    Odrv4 I__16876 (
            .O(N__74265),
            .I(side_command_4));
    InMux I__16875 (
            .O(N__74262),
            .I(bfn_18_18_0_));
    InMux I__16874 (
            .O(N__74259),
            .I(N__74256));
    LocalMux I__16873 (
            .O(N__74256),
            .I(N__74253));
    Span4Mux_h I__16872 (
            .O(N__74253),
            .I(N__74250));
    Span4Mux_h I__16871 (
            .O(N__74250),
            .I(N__74247));
    Odrv4 I__16870 (
            .O(N__74247),
            .I(drone_H_disp_side_i_9));
    CascadeMux I__16869 (
            .O(N__74244),
            .I(N__74241));
    InMux I__16868 (
            .O(N__74241),
            .I(N__74238));
    LocalMux I__16867 (
            .O(N__74238),
            .I(N__74235));
    Odrv12 I__16866 (
            .O(N__74235),
            .I(side_command_5));
    InMux I__16865 (
            .O(N__74232),
            .I(\pid_side.error_cry_4 ));
    InMux I__16864 (
            .O(N__74229),
            .I(N__74226));
    LocalMux I__16863 (
            .O(N__74226),
            .I(N__74223));
    Span4Mux_h I__16862 (
            .O(N__74223),
            .I(N__74220));
    Span4Mux_h I__16861 (
            .O(N__74220),
            .I(N__74217));
    Odrv4 I__16860 (
            .O(N__74217),
            .I(drone_H_disp_side_i_10));
    CascadeMux I__16859 (
            .O(N__74214),
            .I(N__74211));
    InMux I__16858 (
            .O(N__74211),
            .I(N__74208));
    LocalMux I__16857 (
            .O(N__74208),
            .I(N__74205));
    Odrv4 I__16856 (
            .O(N__74205),
            .I(side_command_6));
    InMux I__16855 (
            .O(N__74202),
            .I(\pid_side.error_cry_5 ));
    InMux I__16854 (
            .O(N__74199),
            .I(N__74196));
    LocalMux I__16853 (
            .O(N__74196),
            .I(\pid_side.error_axbZ0Z_7 ));
    InMux I__16852 (
            .O(N__74193),
            .I(N__74190));
    LocalMux I__16851 (
            .O(N__74190),
            .I(N__74185));
    InMux I__16850 (
            .O(N__74189),
            .I(N__74182));
    InMux I__16849 (
            .O(N__74188),
            .I(N__74178));
    Span4Mux_v I__16848 (
            .O(N__74185),
            .I(N__74173));
    LocalMux I__16847 (
            .O(N__74182),
            .I(N__74170));
    InMux I__16846 (
            .O(N__74181),
            .I(N__74167));
    LocalMux I__16845 (
            .O(N__74178),
            .I(N__74161));
    InMux I__16844 (
            .O(N__74177),
            .I(N__74156));
    InMux I__16843 (
            .O(N__74176),
            .I(N__74156));
    Span4Mux_v I__16842 (
            .O(N__74173),
            .I(N__74153));
    Span4Mux_s3_h I__16841 (
            .O(N__74170),
            .I(N__74149));
    LocalMux I__16840 (
            .O(N__74167),
            .I(N__74146));
    InMux I__16839 (
            .O(N__74166),
            .I(N__74139));
    InMux I__16838 (
            .O(N__74165),
            .I(N__74139));
    InMux I__16837 (
            .O(N__74164),
            .I(N__74139));
    Span4Mux_h I__16836 (
            .O(N__74161),
            .I(N__74134));
    LocalMux I__16835 (
            .O(N__74156),
            .I(N__74134));
    Span4Mux_h I__16834 (
            .O(N__74153),
            .I(N__74131));
    InMux I__16833 (
            .O(N__74152),
            .I(N__74128));
    Span4Mux_h I__16832 (
            .O(N__74149),
            .I(N__74123));
    Span4Mux_h I__16831 (
            .O(N__74146),
            .I(N__74123));
    LocalMux I__16830 (
            .O(N__74139),
            .I(N__74118));
    Span4Mux_v I__16829 (
            .O(N__74134),
            .I(N__74118));
    Odrv4 I__16828 (
            .O(N__74131),
            .I(\pid_side.error_11 ));
    LocalMux I__16827 (
            .O(N__74128),
            .I(\pid_side.error_11 ));
    Odrv4 I__16826 (
            .O(N__74123),
            .I(\pid_side.error_11 ));
    Odrv4 I__16825 (
            .O(N__74118),
            .I(\pid_side.error_11 ));
    InMux I__16824 (
            .O(N__74109),
            .I(\pid_side.error_cry_6 ));
    InMux I__16823 (
            .O(N__74106),
            .I(N__74103));
    LocalMux I__16822 (
            .O(N__74103),
            .I(\pid_side.error_axb_8_l_ofxZ0 ));
    CascadeMux I__16821 (
            .O(N__74100),
            .I(N__74097));
    InMux I__16820 (
            .O(N__74097),
            .I(N__74094));
    LocalMux I__16819 (
            .O(N__74094),
            .I(N__74089));
    InMux I__16818 (
            .O(N__74093),
            .I(N__74084));
    InMux I__16817 (
            .O(N__74092),
            .I(N__74084));
    Span4Mux_h I__16816 (
            .O(N__74089),
            .I(N__74079));
    LocalMux I__16815 (
            .O(N__74084),
            .I(N__74079));
    Span4Mux_h I__16814 (
            .O(N__74079),
            .I(N__74076));
    Odrv4 I__16813 (
            .O(N__74076),
            .I(drone_H_disp_side_12));
    InMux I__16812 (
            .O(N__74073),
            .I(N__74068));
    InMux I__16811 (
            .O(N__74072),
            .I(N__74064));
    InMux I__16810 (
            .O(N__74071),
            .I(N__74060));
    LocalMux I__16809 (
            .O(N__74068),
            .I(N__74057));
    InMux I__16808 (
            .O(N__74067),
            .I(N__74053));
    LocalMux I__16807 (
            .O(N__74064),
            .I(N__74050));
    InMux I__16806 (
            .O(N__74063),
            .I(N__74045));
    LocalMux I__16805 (
            .O(N__74060),
            .I(N__74042));
    Span4Mux_s2_h I__16804 (
            .O(N__74057),
            .I(N__74039));
    InMux I__16803 (
            .O(N__74056),
            .I(N__74035));
    LocalMux I__16802 (
            .O(N__74053),
            .I(N__74030));
    Span4Mux_h I__16801 (
            .O(N__74050),
            .I(N__74030));
    InMux I__16800 (
            .O(N__74049),
            .I(N__74025));
    InMux I__16799 (
            .O(N__74048),
            .I(N__74025));
    LocalMux I__16798 (
            .O(N__74045),
            .I(N__74022));
    Span4Mux_s2_h I__16797 (
            .O(N__74042),
            .I(N__74019));
    Span4Mux_v I__16796 (
            .O(N__74039),
            .I(N__74016));
    InMux I__16795 (
            .O(N__74038),
            .I(N__74013));
    LocalMux I__16794 (
            .O(N__74035),
            .I(N__74006));
    Span4Mux_v I__16793 (
            .O(N__74030),
            .I(N__74006));
    LocalMux I__16792 (
            .O(N__74025),
            .I(N__74006));
    Span4Mux_h I__16791 (
            .O(N__74022),
            .I(N__74001));
    Span4Mux_h I__16790 (
            .O(N__74019),
            .I(N__74001));
    Span4Mux_h I__16789 (
            .O(N__74016),
            .I(N__73998));
    LocalMux I__16788 (
            .O(N__74013),
            .I(\pid_side.error_12 ));
    Odrv4 I__16787 (
            .O(N__74006),
            .I(\pid_side.error_12 ));
    Odrv4 I__16786 (
            .O(N__74001),
            .I(\pid_side.error_12 ));
    Odrv4 I__16785 (
            .O(N__73998),
            .I(\pid_side.error_12 ));
    InMux I__16784 (
            .O(N__73989),
            .I(\pid_side.error_cry_7 ));
    InMux I__16783 (
            .O(N__73986),
            .I(N__73983));
    LocalMux I__16782 (
            .O(N__73983),
            .I(drone_H_disp_side_i_12));
    CascadeMux I__16781 (
            .O(N__73980),
            .I(N__73977));
    InMux I__16780 (
            .O(N__73977),
            .I(N__73974));
    LocalMux I__16779 (
            .O(N__73974),
            .I(N__73970));
    InMux I__16778 (
            .O(N__73973),
            .I(N__73967));
    Span4Mux_h I__16777 (
            .O(N__73970),
            .I(N__73962));
    LocalMux I__16776 (
            .O(N__73967),
            .I(N__73962));
    Span4Mux_h I__16775 (
            .O(N__73962),
            .I(N__73959));
    Odrv4 I__16774 (
            .O(N__73959),
            .I(drone_H_disp_side_13));
    InMux I__16773 (
            .O(N__73956),
            .I(\pid_side.error_cry_8 ));
    InMux I__16772 (
            .O(N__73953),
            .I(N__73950));
    LocalMux I__16771 (
            .O(N__73950),
            .I(N__73947));
    Odrv4 I__16770 (
            .O(N__73947),
            .I(drone_H_disp_side_i_13));
    InMux I__16769 (
            .O(N__73944),
            .I(\pid_side.error_cry_9 ));
    InMux I__16768 (
            .O(N__73941),
            .I(N__73935));
    InMux I__16767 (
            .O(N__73940),
            .I(N__73935));
    LocalMux I__16766 (
            .O(N__73935),
            .I(N__73932));
    Odrv4 I__16765 (
            .O(N__73932),
            .I(side_command_7));
    CEMux I__16764 (
            .O(N__73929),
            .I(N__73926));
    LocalMux I__16763 (
            .O(N__73926),
            .I(N__73923));
    Span4Mux_h I__16762 (
            .O(N__73923),
            .I(N__73920));
    Sp12to4 I__16761 (
            .O(N__73920),
            .I(N__73917));
    Span12Mux_v I__16760 (
            .O(N__73917),
            .I(N__73914));
    Odrv12 I__16759 (
            .O(N__73914),
            .I(\Commands_frame_decoder.source_CH2data_1_sqmuxa_0 ));
    InMux I__16758 (
            .O(N__73911),
            .I(N__73908));
    LocalMux I__16757 (
            .O(N__73908),
            .I(N__73905));
    Odrv12 I__16756 (
            .O(N__73905),
            .I(dron_frame_decoder_1_source_H_disp_side_fast_0));
    InMux I__16755 (
            .O(N__73902),
            .I(N__73899));
    LocalMux I__16754 (
            .O(N__73899),
            .I(\pid_side.error_axb_0 ));
    InMux I__16753 (
            .O(N__73896),
            .I(N__73893));
    LocalMux I__16752 (
            .O(N__73893),
            .I(N__73890));
    Span4Mux_h I__16751 (
            .O(N__73890),
            .I(N__73887));
    Span4Mux_h I__16750 (
            .O(N__73887),
            .I(N__73884));
    Odrv4 I__16749 (
            .O(N__73884),
            .I(\pid_side.error_axbZ0Z_1 ));
    InMux I__16748 (
            .O(N__73881),
            .I(N__73878));
    LocalMux I__16747 (
            .O(N__73878),
            .I(N__73874));
    InMux I__16746 (
            .O(N__73877),
            .I(N__73869));
    Span4Mux_v I__16745 (
            .O(N__73874),
            .I(N__73864));
    InMux I__16744 (
            .O(N__73873),
            .I(N__73861));
    InMux I__16743 (
            .O(N__73872),
            .I(N__73858));
    LocalMux I__16742 (
            .O(N__73869),
            .I(N__73855));
    InMux I__16741 (
            .O(N__73868),
            .I(N__73850));
    InMux I__16740 (
            .O(N__73867),
            .I(N__73850));
    Span4Mux_v I__16739 (
            .O(N__73864),
            .I(N__73847));
    LocalMux I__16738 (
            .O(N__73861),
            .I(N__73844));
    LocalMux I__16737 (
            .O(N__73858),
            .I(N__73839));
    Span4Mux_v I__16736 (
            .O(N__73855),
            .I(N__73839));
    LocalMux I__16735 (
            .O(N__73850),
            .I(N__73836));
    Span4Mux_h I__16734 (
            .O(N__73847),
            .I(N__73833));
    Span4Mux_s3_h I__16733 (
            .O(N__73844),
            .I(N__73830));
    Span4Mux_h I__16732 (
            .O(N__73839),
            .I(N__73825));
    Span4Mux_h I__16731 (
            .O(N__73836),
            .I(N__73825));
    Odrv4 I__16730 (
            .O(N__73833),
            .I(\pid_side.error_1 ));
    Odrv4 I__16729 (
            .O(N__73830),
            .I(\pid_side.error_1 ));
    Odrv4 I__16728 (
            .O(N__73825),
            .I(\pid_side.error_1 ));
    InMux I__16727 (
            .O(N__73818),
            .I(\pid_side.error_cry_0 ));
    InMux I__16726 (
            .O(N__73815),
            .I(N__73812));
    LocalMux I__16725 (
            .O(N__73812),
            .I(N__73809));
    Odrv12 I__16724 (
            .O(N__73809),
            .I(\pid_side.error_axbZ0Z_2 ));
    InMux I__16723 (
            .O(N__73806),
            .I(\pid_side.error_cry_1 ));
    InMux I__16722 (
            .O(N__73803),
            .I(N__73800));
    LocalMux I__16721 (
            .O(N__73800),
            .I(N__73797));
    Odrv12 I__16720 (
            .O(N__73797),
            .I(\pid_side.error_axbZ0Z_3 ));
    InMux I__16719 (
            .O(N__73794),
            .I(\pid_side.error_cry_2 ));
    InMux I__16718 (
            .O(N__73791),
            .I(N__73788));
    LocalMux I__16717 (
            .O(N__73788),
            .I(N__73785));
    Odrv12 I__16716 (
            .O(N__73785),
            .I(drone_H_disp_side_i_4));
    CascadeMux I__16715 (
            .O(N__73782),
            .I(N__73779));
    InMux I__16714 (
            .O(N__73779),
            .I(N__73776));
    LocalMux I__16713 (
            .O(N__73776),
            .I(side_command_0));
    InMux I__16712 (
            .O(N__73773),
            .I(\pid_side.error_cry_3 ));
    InMux I__16711 (
            .O(N__73770),
            .I(N__73767));
    LocalMux I__16710 (
            .O(N__73767),
            .I(N__73764));
    Odrv12 I__16709 (
            .O(N__73764),
            .I(drone_H_disp_side_i_5));
    CascadeMux I__16708 (
            .O(N__73761),
            .I(N__73758));
    InMux I__16707 (
            .O(N__73758),
            .I(N__73755));
    LocalMux I__16706 (
            .O(N__73755),
            .I(side_command_1));
    InMux I__16705 (
            .O(N__73752),
            .I(\pid_side.error_cry_0_0 ));
    InMux I__16704 (
            .O(N__73749),
            .I(N__73746));
    LocalMux I__16703 (
            .O(N__73746),
            .I(side_command_2));
    CascadeMux I__16702 (
            .O(N__73743),
            .I(N__73740));
    InMux I__16701 (
            .O(N__73740),
            .I(N__73737));
    LocalMux I__16700 (
            .O(N__73737),
            .I(N__73734));
    Odrv12 I__16699 (
            .O(N__73734),
            .I(drone_H_disp_side_i_6));
    InMux I__16698 (
            .O(N__73731),
            .I(\pid_side.error_cry_1_0 ));
    CascadeMux I__16697 (
            .O(N__73728),
            .I(\pid_side.un1_pid_prereg_0_9_cascade_ ));
    CascadeMux I__16696 (
            .O(N__73725),
            .I(N__73722));
    InMux I__16695 (
            .O(N__73722),
            .I(N__73718));
    InMux I__16694 (
            .O(N__73721),
            .I(N__73715));
    LocalMux I__16693 (
            .O(N__73718),
            .I(\pid_side.un1_pid_prereg_0_8 ));
    LocalMux I__16692 (
            .O(N__73715),
            .I(\pid_side.un1_pid_prereg_0_8 ));
    CascadeMux I__16691 (
            .O(N__73710),
            .I(N__73707));
    InMux I__16690 (
            .O(N__73707),
            .I(N__73704));
    LocalMux I__16689 (
            .O(N__73704),
            .I(N__73701));
    Span4Mux_h I__16688 (
            .O(N__73701),
            .I(N__73698));
    Odrv4 I__16687 (
            .O(N__73698),
            .I(\pid_side.error_d_reg_prev_esr_RNIIOAQ4Z0Z_18 ));
    InMux I__16686 (
            .O(N__73695),
            .I(N__73692));
    LocalMux I__16685 (
            .O(N__73692),
            .I(N__73688));
    InMux I__16684 (
            .O(N__73691),
            .I(N__73685));
    Span4Mux_h I__16683 (
            .O(N__73688),
            .I(N__73682));
    LocalMux I__16682 (
            .O(N__73685),
            .I(N__73679));
    Odrv4 I__16681 (
            .O(N__73682),
            .I(\pid_side.un1_pid_prereg_0 ));
    Odrv4 I__16680 (
            .O(N__73679),
            .I(\pid_side.un1_pid_prereg_0 ));
    CascadeMux I__16679 (
            .O(N__73674),
            .I(N__73671));
    InMux I__16678 (
            .O(N__73671),
            .I(N__73668));
    LocalMux I__16677 (
            .O(N__73668),
            .I(N__73665));
    Span4Mux_v I__16676 (
            .O(N__73665),
            .I(N__73662));
    Span4Mux_h I__16675 (
            .O(N__73662),
            .I(N__73659));
    Odrv4 I__16674 (
            .O(N__73659),
            .I(\pid_side.error_d_reg_prev_esr_RNIQ8P41Z0Z_0 ));
    InMux I__16673 (
            .O(N__73656),
            .I(N__73652));
    InMux I__16672 (
            .O(N__73655),
            .I(N__73647));
    LocalMux I__16671 (
            .O(N__73652),
            .I(N__73643));
    InMux I__16670 (
            .O(N__73651),
            .I(N__73640));
    InMux I__16669 (
            .O(N__73650),
            .I(N__73635));
    LocalMux I__16668 (
            .O(N__73647),
            .I(N__73632));
    InMux I__16667 (
            .O(N__73646),
            .I(N__73629));
    Span4Mux_h I__16666 (
            .O(N__73643),
            .I(N__73623));
    LocalMux I__16665 (
            .O(N__73640),
            .I(N__73620));
    InMux I__16664 (
            .O(N__73639),
            .I(N__73617));
    InMux I__16663 (
            .O(N__73638),
            .I(N__73614));
    LocalMux I__16662 (
            .O(N__73635),
            .I(N__73611));
    Span4Mux_v I__16661 (
            .O(N__73632),
            .I(N__73606));
    LocalMux I__16660 (
            .O(N__73629),
            .I(N__73606));
    InMux I__16659 (
            .O(N__73628),
            .I(N__73602));
    InMux I__16658 (
            .O(N__73627),
            .I(N__73599));
    InMux I__16657 (
            .O(N__73626),
            .I(N__73596));
    Span4Mux_h I__16656 (
            .O(N__73623),
            .I(N__73591));
    Span4Mux_v I__16655 (
            .O(N__73620),
            .I(N__73591));
    LocalMux I__16654 (
            .O(N__73617),
            .I(N__73585));
    LocalMux I__16653 (
            .O(N__73614),
            .I(N__73585));
    Span4Mux_v I__16652 (
            .O(N__73611),
            .I(N__73580));
    Span4Mux_v I__16651 (
            .O(N__73606),
            .I(N__73580));
    InMux I__16650 (
            .O(N__73605),
            .I(N__73576));
    LocalMux I__16649 (
            .O(N__73602),
            .I(N__73573));
    LocalMux I__16648 (
            .O(N__73599),
            .I(N__73570));
    LocalMux I__16647 (
            .O(N__73596),
            .I(N__73567));
    Span4Mux_h I__16646 (
            .O(N__73591),
            .I(N__73564));
    CascadeMux I__16645 (
            .O(N__73590),
            .I(N__73560));
    Span4Mux_v I__16644 (
            .O(N__73585),
            .I(N__73555));
    Span4Mux_h I__16643 (
            .O(N__73580),
            .I(N__73555));
    InMux I__16642 (
            .O(N__73579),
            .I(N__73552));
    LocalMux I__16641 (
            .O(N__73576),
            .I(N__73547));
    Span4Mux_v I__16640 (
            .O(N__73573),
            .I(N__73547));
    Span4Mux_v I__16639 (
            .O(N__73570),
            .I(N__73540));
    Span4Mux_v I__16638 (
            .O(N__73567),
            .I(N__73540));
    Span4Mux_h I__16637 (
            .O(N__73564),
            .I(N__73540));
    InMux I__16636 (
            .O(N__73563),
            .I(N__73537));
    InMux I__16635 (
            .O(N__73560),
            .I(N__73534));
    Span4Mux_h I__16634 (
            .O(N__73555),
            .I(N__73529));
    LocalMux I__16633 (
            .O(N__73552),
            .I(N__73529));
    Span4Mux_v I__16632 (
            .O(N__73547),
            .I(N__73522));
    Span4Mux_v I__16631 (
            .O(N__73540),
            .I(N__73522));
    LocalMux I__16630 (
            .O(N__73537),
            .I(N__73522));
    LocalMux I__16629 (
            .O(N__73534),
            .I(uart_pc_data_6));
    Odrv4 I__16628 (
            .O(N__73529),
            .I(uart_pc_data_6));
    Odrv4 I__16627 (
            .O(N__73522),
            .I(uart_pc_data_6));
    InMux I__16626 (
            .O(N__73515),
            .I(N__73510));
    InMux I__16625 (
            .O(N__73514),
            .I(N__73505));
    InMux I__16624 (
            .O(N__73513),
            .I(N__73505));
    LocalMux I__16623 (
            .O(N__73510),
            .I(\pid_side.un1_pid_prereg_0_11 ));
    LocalMux I__16622 (
            .O(N__73505),
            .I(\pid_side.un1_pid_prereg_0_11 ));
    InMux I__16621 (
            .O(N__73500),
            .I(N__73494));
    InMux I__16620 (
            .O(N__73499),
            .I(N__73494));
    LocalMux I__16619 (
            .O(N__73494),
            .I(\pid_side.un1_pid_prereg_0_10 ));
    CascadeMux I__16618 (
            .O(N__73491),
            .I(\pid_side.un1_pid_prereg_0_12_cascade_ ));
    InMux I__16617 (
            .O(N__73488),
            .I(N__73485));
    LocalMux I__16616 (
            .O(N__73485),
            .I(\pid_side.error_d_reg_prev_esr_RNIV6JN9Z0Z_19 ));
    InMux I__16615 (
            .O(N__73482),
            .I(N__73478));
    InMux I__16614 (
            .O(N__73481),
            .I(N__73475));
    LocalMux I__16613 (
            .O(N__73478),
            .I(\pid_side.un1_pid_prereg_0_2 ));
    LocalMux I__16612 (
            .O(N__73475),
            .I(\pid_side.un1_pid_prereg_0_2 ));
    CascadeMux I__16611 (
            .O(N__73470),
            .I(N__73467));
    InMux I__16610 (
            .O(N__73467),
            .I(N__73462));
    InMux I__16609 (
            .O(N__73466),
            .I(N__73459));
    InMux I__16608 (
            .O(N__73465),
            .I(N__73456));
    LocalMux I__16607 (
            .O(N__73462),
            .I(\pid_side.un1_pid_prereg_0_3 ));
    LocalMux I__16606 (
            .O(N__73459),
            .I(\pid_side.un1_pid_prereg_0_3 ));
    LocalMux I__16605 (
            .O(N__73456),
            .I(\pid_side.un1_pid_prereg_0_3 ));
    CascadeMux I__16604 (
            .O(N__73449),
            .I(N__73446));
    InMux I__16603 (
            .O(N__73446),
            .I(N__73443));
    LocalMux I__16602 (
            .O(N__73443),
            .I(\pid_side.error_d_reg_prev_esr_RNI620Q4Z0Z_15 ));
    InMux I__16601 (
            .O(N__73440),
            .I(N__73437));
    LocalMux I__16600 (
            .O(N__73437),
            .I(N__73434));
    Span4Mux_h I__16599 (
            .O(N__73434),
            .I(N__73431));
    Sp12to4 I__16598 (
            .O(N__73431),
            .I(N__73427));
    InMux I__16597 (
            .O(N__73430),
            .I(N__73424));
    Odrv12 I__16596 (
            .O(N__73427),
            .I(\pid_side.un1_pid_prereg_0_12 ));
    LocalMux I__16595 (
            .O(N__73424),
            .I(\pid_side.un1_pid_prereg_0_12 ));
    InMux I__16594 (
            .O(N__73419),
            .I(N__73416));
    LocalMux I__16593 (
            .O(N__73416),
            .I(N__73413));
    Span4Mux_v I__16592 (
            .O(N__73413),
            .I(N__73408));
    InMux I__16591 (
            .O(N__73412),
            .I(N__73403));
    InMux I__16590 (
            .O(N__73411),
            .I(N__73403));
    Odrv4 I__16589 (
            .O(N__73408),
            .I(\pid_side.un1_pid_prereg_0_13 ));
    LocalMux I__16588 (
            .O(N__73403),
            .I(\pid_side.un1_pid_prereg_0_13 ));
    InMux I__16587 (
            .O(N__73398),
            .I(N__73395));
    LocalMux I__16586 (
            .O(N__73395),
            .I(N__73392));
    Odrv4 I__16585 (
            .O(N__73392),
            .I(\pid_side.error_d_reg_prev_esr_RNI578S4Z0Z_20 ));
    InMux I__16584 (
            .O(N__73389),
            .I(N__73386));
    LocalMux I__16583 (
            .O(N__73386),
            .I(N__73382));
    InMux I__16582 (
            .O(N__73385),
            .I(N__73379));
    Odrv4 I__16581 (
            .O(N__73382),
            .I(\pid_side.un1_pid_prereg_0_1 ));
    LocalMux I__16580 (
            .O(N__73379),
            .I(\pid_side.un1_pid_prereg_0_1 ));
    InMux I__16579 (
            .O(N__73374),
            .I(N__73367));
    InMux I__16578 (
            .O(N__73373),
            .I(N__73367));
    InMux I__16577 (
            .O(N__73372),
            .I(N__73364));
    LocalMux I__16576 (
            .O(N__73367),
            .I(\pid_side.un1_pid_prereg_0_0 ));
    LocalMux I__16575 (
            .O(N__73364),
            .I(\pid_side.un1_pid_prereg_0_0 ));
    CascadeMux I__16574 (
            .O(N__73359),
            .I(N__73356));
    InMux I__16573 (
            .O(N__73356),
            .I(N__73353));
    LocalMux I__16572 (
            .O(N__73353),
            .I(\pid_side.error_d_reg_prev_esr_RNI1OK5FZ0Z_12 ));
    InMux I__16571 (
            .O(N__73350),
            .I(N__73346));
    InMux I__16570 (
            .O(N__73349),
            .I(N__73343));
    LocalMux I__16569 (
            .O(N__73346),
            .I(N__73339));
    LocalMux I__16568 (
            .O(N__73343),
            .I(N__73336));
    InMux I__16567 (
            .O(N__73342),
            .I(N__73333));
    Odrv12 I__16566 (
            .O(N__73339),
            .I(\pid_side.error_i_reg_esr_RNI2MSRZ0Z_19 ));
    Odrv4 I__16565 (
            .O(N__73336),
            .I(\pid_side.error_i_reg_esr_RNI2MSRZ0Z_19 ));
    LocalMux I__16564 (
            .O(N__73333),
            .I(\pid_side.error_i_reg_esr_RNI2MSRZ0Z_19 ));
    InMux I__16563 (
            .O(N__73326),
            .I(N__73322));
    InMux I__16562 (
            .O(N__73325),
            .I(N__73319));
    LocalMux I__16561 (
            .O(N__73322),
            .I(\pid_side.un1_pid_prereg_0_7 ));
    LocalMux I__16560 (
            .O(N__73319),
            .I(\pid_side.un1_pid_prereg_0_7 ));
    InMux I__16559 (
            .O(N__73314),
            .I(N__73310));
    InMux I__16558 (
            .O(N__73313),
            .I(N__73307));
    LocalMux I__16557 (
            .O(N__73310),
            .I(\pid_side.un1_pid_prereg_0_6 ));
    LocalMux I__16556 (
            .O(N__73307),
            .I(\pid_side.un1_pid_prereg_0_6 ));
    CascadeMux I__16555 (
            .O(N__73302),
            .I(\pid_side.un1_pid_prereg_0_8_cascade_ ));
    InMux I__16554 (
            .O(N__73299),
            .I(N__73296));
    LocalMux I__16553 (
            .O(N__73296),
            .I(N__73293));
    Odrv4 I__16552 (
            .O(N__73293),
            .I(\pid_side.error_d_reg_prev_esr_RNIOVFK9Z0Z_17 ));
    InMux I__16551 (
            .O(N__73290),
            .I(N__73286));
    InMux I__16550 (
            .O(N__73289),
            .I(N__73282));
    LocalMux I__16549 (
            .O(N__73286),
            .I(N__73279));
    InMux I__16548 (
            .O(N__73285),
            .I(N__73276));
    LocalMux I__16547 (
            .O(N__73282),
            .I(N__73273));
    Span4Mux_v I__16546 (
            .O(N__73279),
            .I(N__73270));
    LocalMux I__16545 (
            .O(N__73276),
            .I(N__73267));
    Span4Mux_h I__16544 (
            .O(N__73273),
            .I(N__73264));
    Odrv4 I__16543 (
            .O(N__73270),
            .I(\pid_side.error_i_reg_esr_RNIRGURZ0Z_20 ));
    Odrv4 I__16542 (
            .O(N__73267),
            .I(\pid_side.error_i_reg_esr_RNIRGURZ0Z_20 ));
    Odrv4 I__16541 (
            .O(N__73264),
            .I(\pid_side.error_i_reg_esr_RNIRGURZ0Z_20 ));
    InMux I__16540 (
            .O(N__73257),
            .I(N__73254));
    LocalMux I__16539 (
            .O(N__73254),
            .I(N__73250));
    InMux I__16538 (
            .O(N__73253),
            .I(N__73247));
    Odrv4 I__16537 (
            .O(N__73250),
            .I(\pid_side.un1_pid_prereg_0_9 ));
    LocalMux I__16536 (
            .O(N__73247),
            .I(\pid_side.un1_pid_prereg_0_9 ));
    CascadeMux I__16535 (
            .O(N__73242),
            .I(\pid_side.un1_pid_prereg_0_21_cascade_ ));
    InMux I__16534 (
            .O(N__73239),
            .I(N__73236));
    LocalMux I__16533 (
            .O(N__73236),
            .I(N__73233));
    Span4Mux_v I__16532 (
            .O(N__73233),
            .I(N__73230));
    Sp12to4 I__16531 (
            .O(N__73230),
            .I(N__73226));
    InMux I__16530 (
            .O(N__73229),
            .I(N__73223));
    Odrv12 I__16529 (
            .O(N__73226),
            .I(\pid_side.un1_pid_prereg_0_20 ));
    LocalMux I__16528 (
            .O(N__73223),
            .I(\pid_side.un1_pid_prereg_0_20 ));
    InMux I__16527 (
            .O(N__73218),
            .I(N__73215));
    LocalMux I__16526 (
            .O(N__73215),
            .I(\pid_side.error_d_reg_prev_esr_RNISK5B3Z0Z_22 ));
    CascadeMux I__16525 (
            .O(N__73212),
            .I(N__73201));
    CascadeMux I__16524 (
            .O(N__73211),
            .I(N__73198));
    CascadeMux I__16523 (
            .O(N__73210),
            .I(N__73195));
    CascadeMux I__16522 (
            .O(N__73209),
            .I(N__73191));
    CascadeMux I__16521 (
            .O(N__73208),
            .I(N__73187));
    CascadeMux I__16520 (
            .O(N__73207),
            .I(N__73183));
    CascadeMux I__16519 (
            .O(N__73206),
            .I(N__73179));
    CascadeMux I__16518 (
            .O(N__73205),
            .I(N__73176));
    InMux I__16517 (
            .O(N__73204),
            .I(N__73167));
    InMux I__16516 (
            .O(N__73201),
            .I(N__73167));
    InMux I__16515 (
            .O(N__73198),
            .I(N__73167));
    InMux I__16514 (
            .O(N__73195),
            .I(N__73167));
    InMux I__16513 (
            .O(N__73194),
            .I(N__73162));
    InMux I__16512 (
            .O(N__73191),
            .I(N__73162));
    InMux I__16511 (
            .O(N__73190),
            .I(N__73157));
    InMux I__16510 (
            .O(N__73187),
            .I(N__73157));
    InMux I__16509 (
            .O(N__73186),
            .I(N__73154));
    InMux I__16508 (
            .O(N__73183),
            .I(N__73149));
    InMux I__16507 (
            .O(N__73182),
            .I(N__73149));
    InMux I__16506 (
            .O(N__73179),
            .I(N__73144));
    InMux I__16505 (
            .O(N__73176),
            .I(N__73144));
    LocalMux I__16504 (
            .O(N__73167),
            .I(N__73141));
    LocalMux I__16503 (
            .O(N__73162),
            .I(N__73136));
    LocalMux I__16502 (
            .O(N__73157),
            .I(N__73136));
    LocalMux I__16501 (
            .O(N__73154),
            .I(N__73131));
    LocalMux I__16500 (
            .O(N__73149),
            .I(N__73131));
    LocalMux I__16499 (
            .O(N__73144),
            .I(N__73128));
    Span4Mux_v I__16498 (
            .O(N__73141),
            .I(N__73125));
    Span4Mux_v I__16497 (
            .O(N__73136),
            .I(N__73120));
    Span4Mux_h I__16496 (
            .O(N__73131),
            .I(N__73120));
    Odrv4 I__16495 (
            .O(N__73128),
            .I(\pid_side.error_d_reg_prevZ0Z_22 ));
    Odrv4 I__16494 (
            .O(N__73125),
            .I(\pid_side.error_d_reg_prevZ0Z_22 ));
    Odrv4 I__16493 (
            .O(N__73120),
            .I(\pid_side.error_d_reg_prevZ0Z_22 ));
    InMux I__16492 (
            .O(N__73113),
            .I(N__73107));
    InMux I__16491 (
            .O(N__73112),
            .I(N__73107));
    LocalMux I__16490 (
            .O(N__73107),
            .I(\pid_side.error_d_reg_prevZ0Z_21 ));
    InMux I__16489 (
            .O(N__73104),
            .I(N__73100));
    InMux I__16488 (
            .O(N__73103),
            .I(N__73097));
    LocalMux I__16487 (
            .O(N__73100),
            .I(N__73094));
    LocalMux I__16486 (
            .O(N__73097),
            .I(N__73091));
    Span4Mux_h I__16485 (
            .O(N__73094),
            .I(N__73088));
    Span4Mux_h I__16484 (
            .O(N__73091),
            .I(N__73085));
    Odrv4 I__16483 (
            .O(N__73088),
            .I(\pid_side.error_d_reg_prev_esr_RNIVNLOZ0Z_21 ));
    Odrv4 I__16482 (
            .O(N__73085),
            .I(\pid_side.error_d_reg_prev_esr_RNIVNLOZ0Z_21 ));
    InMux I__16481 (
            .O(N__73080),
            .I(N__73077));
    LocalMux I__16480 (
            .O(N__73077),
            .I(\pid_side.error_d_reg_prev_esr_RNICOLL9Z0Z_18 ));
    CascadeMux I__16479 (
            .O(N__73074),
            .I(\pid_side.un1_pid_prereg_0_10_cascade_ ));
    CascadeMux I__16478 (
            .O(N__73071),
            .I(N__73068));
    InMux I__16477 (
            .O(N__73068),
            .I(N__73065));
    LocalMux I__16476 (
            .O(N__73065),
            .I(N__73062));
    Odrv4 I__16475 (
            .O(N__73062),
            .I(\pid_side.error_d_reg_prev_esr_RNIQVAR4Z0Z_19 ));
    InMux I__16474 (
            .O(N__73059),
            .I(N__73055));
    InMux I__16473 (
            .O(N__73058),
            .I(N__73052));
    LocalMux I__16472 (
            .O(N__73055),
            .I(N__73049));
    LocalMux I__16471 (
            .O(N__73052),
            .I(\pid_side.error_d_reg_prev_esr_RNIVNLO_0Z0Z_21 ));
    Odrv4 I__16470 (
            .O(N__73049),
            .I(\pid_side.error_d_reg_prev_esr_RNIVNLO_0Z0Z_21 ));
    InMux I__16469 (
            .O(N__73044),
            .I(N__73040));
    InMux I__16468 (
            .O(N__73043),
            .I(N__73037));
    LocalMux I__16467 (
            .O(N__73040),
            .I(N__73034));
    LocalMux I__16466 (
            .O(N__73037),
            .I(N__73031));
    Span4Mux_v I__16465 (
            .O(N__73034),
            .I(N__73027));
    Span4Mux_h I__16464 (
            .O(N__73031),
            .I(N__73024));
    InMux I__16463 (
            .O(N__73030),
            .I(N__73021));
    Odrv4 I__16462 (
            .O(N__73027),
            .I(\pid_side.error_i_reg_esr_RNIK2OSZ0Z_21 ));
    Odrv4 I__16461 (
            .O(N__73024),
            .I(\pid_side.error_i_reg_esr_RNIK2OSZ0Z_21 ));
    LocalMux I__16460 (
            .O(N__73021),
            .I(\pid_side.error_i_reg_esr_RNIK2OSZ0Z_21 ));
    InMux I__16459 (
            .O(N__73014),
            .I(N__73008));
    InMux I__16458 (
            .O(N__73013),
            .I(N__73008));
    LocalMux I__16457 (
            .O(N__73008),
            .I(N__73005));
    Odrv12 I__16456 (
            .O(N__73005),
            .I(\pid_side.N_2380_i ));
    CascadeMux I__16455 (
            .O(N__73002),
            .I(N__72998));
    CascadeMux I__16454 (
            .O(N__73001),
            .I(N__72995));
    InMux I__16453 (
            .O(N__72998),
            .I(N__72992));
    InMux I__16452 (
            .O(N__72995),
            .I(N__72989));
    LocalMux I__16451 (
            .O(N__72992),
            .I(N__72984));
    LocalMux I__16450 (
            .O(N__72989),
            .I(N__72984));
    Span4Mux_h I__16449 (
            .O(N__72984),
            .I(N__72981));
    Odrv4 I__16448 (
            .O(N__72981),
            .I(\pid_side.error_p_reg_esr_RNIIAPH3Z0Z_8 ));
    InMux I__16447 (
            .O(N__72978),
            .I(N__72975));
    LocalMux I__16446 (
            .O(N__72975),
            .I(\pid_side.error_p_reg_esr_RNIKGHS6Z0Z_10 ));
    CascadeMux I__16445 (
            .O(N__72972),
            .I(\pid_side.N_2386_i_cascade_ ));
    InMux I__16444 (
            .O(N__72969),
            .I(N__72966));
    LocalMux I__16443 (
            .O(N__72966),
            .I(\pid_side.error_p_reg_esr_RNIRE1B1Z0Z_10 ));
    InMux I__16442 (
            .O(N__72963),
            .I(N__72959));
    InMux I__16441 (
            .O(N__72962),
            .I(N__72956));
    LocalMux I__16440 (
            .O(N__72959),
            .I(\pid_side.error_d_reg_prev_esr_RNITU3P4_0Z0Z_10 ));
    LocalMux I__16439 (
            .O(N__72956),
            .I(\pid_side.error_d_reg_prev_esr_RNITU3P4_0Z0Z_10 ));
    InMux I__16438 (
            .O(N__72951),
            .I(N__72945));
    InMux I__16437 (
            .O(N__72950),
            .I(N__72945));
    LocalMux I__16436 (
            .O(N__72945),
            .I(N__72942));
    Span4Mux_h I__16435 (
            .O(N__72942),
            .I(N__72939));
    Odrv4 I__16434 (
            .O(N__72939),
            .I(\pid_side.error_p_reg_esr_RNI1VTC1Z0Z_9 ));
    CascadeMux I__16433 (
            .O(N__72936),
            .I(\pid_side.error_p_reg_esr_RNIRE1B1Z0Z_10_cascade_ ));
    InMux I__16432 (
            .O(N__72933),
            .I(N__72928));
    InMux I__16431 (
            .O(N__72932),
            .I(N__72923));
    InMux I__16430 (
            .O(N__72931),
            .I(N__72923));
    LocalMux I__16429 (
            .O(N__72928),
            .I(N__72920));
    LocalMux I__16428 (
            .O(N__72923),
            .I(N__72917));
    Span4Mux_v I__16427 (
            .O(N__72920),
            .I(N__72912));
    Span4Mux_v I__16426 (
            .O(N__72917),
            .I(N__72912));
    Odrv4 I__16425 (
            .O(N__72912),
            .I(\pid_side.error_i_reg_esr_RNI6OOIZ0Z_10 ));
    CascadeMux I__16424 (
            .O(N__72909),
            .I(N__72906));
    InMux I__16423 (
            .O(N__72906),
            .I(N__72903));
    LocalMux I__16422 (
            .O(N__72903),
            .I(\pid_side.error_p_reg_esr_RNIV4S38Z0Z_10 ));
    InMux I__16421 (
            .O(N__72900),
            .I(N__72896));
    InMux I__16420 (
            .O(N__72899),
            .I(N__72893));
    LocalMux I__16419 (
            .O(N__72896),
            .I(N__72889));
    LocalMux I__16418 (
            .O(N__72893),
            .I(N__72886));
    InMux I__16417 (
            .O(N__72892),
            .I(N__72883));
    Span4Mux_h I__16416 (
            .O(N__72889),
            .I(N__72880));
    Span4Mux_v I__16415 (
            .O(N__72886),
            .I(N__72877));
    LocalMux I__16414 (
            .O(N__72883),
            .I(\pid_side.error_i_reg_esr_RNISESSZ0Z_25 ));
    Odrv4 I__16413 (
            .O(N__72880),
            .I(\pid_side.error_i_reg_esr_RNISESSZ0Z_25 ));
    Odrv4 I__16412 (
            .O(N__72877),
            .I(\pid_side.error_i_reg_esr_RNISESSZ0Z_25 ));
    InMux I__16411 (
            .O(N__72870),
            .I(N__72867));
    LocalMux I__16410 (
            .O(N__72867),
            .I(N__72863));
    InMux I__16409 (
            .O(N__72866),
            .I(N__72860));
    Odrv4 I__16408 (
            .O(N__72863),
            .I(\pid_side.un1_pid_prereg_0_18 ));
    LocalMux I__16407 (
            .O(N__72860),
            .I(\pid_side.un1_pid_prereg_0_18 ));
    InMux I__16406 (
            .O(N__72855),
            .I(N__72852));
    LocalMux I__16405 (
            .O(N__72852),
            .I(N__72849));
    Span4Mux_v I__16404 (
            .O(N__72849),
            .I(N__72845));
    InMux I__16403 (
            .O(N__72848),
            .I(N__72842));
    Odrv4 I__16402 (
            .O(N__72845),
            .I(\pid_side.un1_pid_prereg_0_19 ));
    LocalMux I__16401 (
            .O(N__72842),
            .I(\pid_side.un1_pid_prereg_0_19 ));
    CascadeMux I__16400 (
            .O(N__72837),
            .I(\pid_side.un1_pid_prereg_0_20_cascade_ ));
    InMux I__16399 (
            .O(N__72834),
            .I(N__72831));
    LocalMux I__16398 (
            .O(N__72831),
            .I(\pid_side.error_d_reg_prev_esr_RNIK39M6Z0Z_22 ));
    InMux I__16397 (
            .O(N__72828),
            .I(N__72823));
    InMux I__16396 (
            .O(N__72827),
            .I(N__72820));
    InMux I__16395 (
            .O(N__72826),
            .I(N__72817));
    LocalMux I__16394 (
            .O(N__72823),
            .I(N__72814));
    LocalMux I__16393 (
            .O(N__72820),
            .I(N__72811));
    LocalMux I__16392 (
            .O(N__72817),
            .I(N__72808));
    Span4Mux_v I__16391 (
            .O(N__72814),
            .I(N__72805));
    Span4Mux_h I__16390 (
            .O(N__72811),
            .I(N__72802));
    Odrv12 I__16389 (
            .O(N__72808),
            .I(\pid_side.error_i_reg_esr_RNIUHTSZ0Z_26 ));
    Odrv4 I__16388 (
            .O(N__72805),
            .I(\pid_side.error_i_reg_esr_RNIUHTSZ0Z_26 ));
    Odrv4 I__16387 (
            .O(N__72802),
            .I(\pid_side.error_i_reg_esr_RNIUHTSZ0Z_26 ));
    InMux I__16386 (
            .O(N__72795),
            .I(N__72792));
    LocalMux I__16385 (
            .O(N__72792),
            .I(N__72789));
    Span4Mux_v I__16384 (
            .O(N__72789),
            .I(N__72785));
    InMux I__16383 (
            .O(N__72788),
            .I(N__72782));
    Odrv4 I__16382 (
            .O(N__72785),
            .I(\pid_side.un1_pid_prereg_0_21 ));
    LocalMux I__16381 (
            .O(N__72782),
            .I(\pid_side.un1_pid_prereg_0_21 ));
    InMux I__16380 (
            .O(N__72777),
            .I(N__72774));
    LocalMux I__16379 (
            .O(N__72774),
            .I(N__72771));
    Odrv4 I__16378 (
            .O(N__72771),
            .I(\pid_side.pid_preregZ0Z_17 ));
    InMux I__16377 (
            .O(N__72768),
            .I(N__72765));
    LocalMux I__16376 (
            .O(N__72765),
            .I(N__72762));
    Odrv4 I__16375 (
            .O(N__72762),
            .I(\pid_side.pid_preregZ0Z_18 ));
    CascadeMux I__16374 (
            .O(N__72759),
            .I(N__72756));
    InMux I__16373 (
            .O(N__72756),
            .I(N__72753));
    LocalMux I__16372 (
            .O(N__72753),
            .I(N__72750));
    Span4Mux_v I__16371 (
            .O(N__72750),
            .I(N__72747));
    Odrv4 I__16370 (
            .O(N__72747),
            .I(\pid_side.pid_preregZ0Z_19 ));
    InMux I__16369 (
            .O(N__72744),
            .I(N__72741));
    LocalMux I__16368 (
            .O(N__72741),
            .I(N__72738));
    Odrv4 I__16367 (
            .O(N__72738),
            .I(\pid_side.pid_preregZ0Z_16 ));
    InMux I__16366 (
            .O(N__72735),
            .I(N__72732));
    LocalMux I__16365 (
            .O(N__72732),
            .I(N__72729));
    Span4Mux_h I__16364 (
            .O(N__72729),
            .I(N__72726));
    Odrv4 I__16363 (
            .O(N__72726),
            .I(\pid_side.un11lto30_i_a2_3_and ));
    CascadeMux I__16362 (
            .O(N__72723),
            .I(N__72720));
    InMux I__16361 (
            .O(N__72720),
            .I(N__72716));
    InMux I__16360 (
            .O(N__72719),
            .I(N__72713));
    LocalMux I__16359 (
            .O(N__72716),
            .I(N__72710));
    LocalMux I__16358 (
            .O(N__72713),
            .I(N__72707));
    Span4Mux_h I__16357 (
            .O(N__72710),
            .I(N__72704));
    Odrv4 I__16356 (
            .O(N__72707),
            .I(\pid_side.pid_preregZ0Z_15 ));
    Odrv4 I__16355 (
            .O(N__72704),
            .I(\pid_side.pid_preregZ0Z_15 ));
    CascadeMux I__16354 (
            .O(N__72699),
            .I(\pid_side.un11lto30_i_a2_3_and_cascade_ ));
    InMux I__16353 (
            .O(N__72696),
            .I(N__72693));
    LocalMux I__16352 (
            .O(N__72693),
            .I(N__72689));
    InMux I__16351 (
            .O(N__72692),
            .I(N__72686));
    Span4Mux_h I__16350 (
            .O(N__72689),
            .I(N__72680));
    LocalMux I__16349 (
            .O(N__72686),
            .I(N__72680));
    InMux I__16348 (
            .O(N__72685),
            .I(N__72677));
    Span4Mux_h I__16347 (
            .O(N__72680),
            .I(N__72674));
    LocalMux I__16346 (
            .O(N__72677),
            .I(\pid_side.pid_preregZ0Z_14 ));
    Odrv4 I__16345 (
            .O(N__72674),
            .I(\pid_side.pid_preregZ0Z_14 ));
    InMux I__16344 (
            .O(N__72669),
            .I(N__72666));
    LocalMux I__16343 (
            .O(N__72666),
            .I(N__72663));
    Span4Mux_h I__16342 (
            .O(N__72663),
            .I(N__72660));
    Odrv4 I__16341 (
            .O(N__72660),
            .I(\pid_side.source_pid_1_sqmuxa_1_0_a2_0_0 ));
    CascadeMux I__16340 (
            .O(N__72657),
            .I(N__72651));
    CascadeMux I__16339 (
            .O(N__72656),
            .I(N__72648));
    CascadeMux I__16338 (
            .O(N__72655),
            .I(N__72645));
    InMux I__16337 (
            .O(N__72654),
            .I(N__72638));
    InMux I__16336 (
            .O(N__72651),
            .I(N__72624));
    InMux I__16335 (
            .O(N__72648),
            .I(N__72624));
    InMux I__16334 (
            .O(N__72645),
            .I(N__72624));
    InMux I__16333 (
            .O(N__72644),
            .I(N__72624));
    InMux I__16332 (
            .O(N__72643),
            .I(N__72624));
    InMux I__16331 (
            .O(N__72642),
            .I(N__72624));
    CascadeMux I__16330 (
            .O(N__72641),
            .I(N__72621));
    LocalMux I__16329 (
            .O(N__72638),
            .I(N__72615));
    CascadeMux I__16328 (
            .O(N__72637),
            .I(N__72610));
    LocalMux I__16327 (
            .O(N__72624),
            .I(N__72607));
    InMux I__16326 (
            .O(N__72621),
            .I(N__72604));
    InMux I__16325 (
            .O(N__72620),
            .I(N__72601));
    InMux I__16324 (
            .O(N__72619),
            .I(N__72596));
    InMux I__16323 (
            .O(N__72618),
            .I(N__72596));
    Span4Mux_v I__16322 (
            .O(N__72615),
            .I(N__72593));
    InMux I__16321 (
            .O(N__72614),
            .I(N__72588));
    InMux I__16320 (
            .O(N__72613),
            .I(N__72588));
    InMux I__16319 (
            .O(N__72610),
            .I(N__72584));
    Span4Mux_h I__16318 (
            .O(N__72607),
            .I(N__72581));
    LocalMux I__16317 (
            .O(N__72604),
            .I(N__72570));
    LocalMux I__16316 (
            .O(N__72601),
            .I(N__72570));
    LocalMux I__16315 (
            .O(N__72596),
            .I(N__72570));
    Span4Mux_h I__16314 (
            .O(N__72593),
            .I(N__72570));
    LocalMux I__16313 (
            .O(N__72588),
            .I(N__72570));
    InMux I__16312 (
            .O(N__72587),
            .I(N__72567));
    LocalMux I__16311 (
            .O(N__72584),
            .I(N__72562));
    Span4Mux_h I__16310 (
            .O(N__72581),
            .I(N__72562));
    Span4Mux_v I__16309 (
            .O(N__72570),
            .I(N__72559));
    LocalMux I__16308 (
            .O(N__72567),
            .I(\pid_side.stateZ0Z_1 ));
    Odrv4 I__16307 (
            .O(N__72562),
            .I(\pid_side.stateZ0Z_1 ));
    Odrv4 I__16306 (
            .O(N__72559),
            .I(\pid_side.stateZ0Z_1 ));
    InMux I__16305 (
            .O(N__72552),
            .I(N__72549));
    LocalMux I__16304 (
            .O(N__72549),
            .I(N__72545));
    CascadeMux I__16303 (
            .O(N__72548),
            .I(N__72541));
    Span4Mux_v I__16302 (
            .O(N__72545),
            .I(N__72538));
    InMux I__16301 (
            .O(N__72544),
            .I(N__72533));
    InMux I__16300 (
            .O(N__72541),
            .I(N__72533));
    Span4Mux_v I__16299 (
            .O(N__72538),
            .I(N__72530));
    LocalMux I__16298 (
            .O(N__72533),
            .I(N__72527));
    Odrv4 I__16297 (
            .O(N__72530),
            .I(\pid_side.error_i_acumm_preregZ0Z_28 ));
    Odrv12 I__16296 (
            .O(N__72527),
            .I(\pid_side.error_i_acumm_preregZ0Z_28 ));
    InMux I__16295 (
            .O(N__72522),
            .I(N__72510));
    InMux I__16294 (
            .O(N__72521),
            .I(N__72510));
    InMux I__16293 (
            .O(N__72520),
            .I(N__72510));
    InMux I__16292 (
            .O(N__72519),
            .I(N__72510));
    LocalMux I__16291 (
            .O(N__72510),
            .I(N__72507));
    Span4Mux_v I__16290 (
            .O(N__72507),
            .I(N__72504));
    Span4Mux_v I__16289 (
            .O(N__72504),
            .I(N__72501));
    Odrv4 I__16288 (
            .O(N__72501),
            .I(\pid_side.error_i_acumm_3_sqmuxa ));
    CascadeMux I__16287 (
            .O(N__72498),
            .I(N__72495));
    InMux I__16286 (
            .O(N__72495),
            .I(N__72492));
    LocalMux I__16285 (
            .O(N__72492),
            .I(\pid_side.error_p_reg_esr_RNI5RKP3Z0Z_5 ));
    CascadeMux I__16284 (
            .O(N__72489),
            .I(N__72486));
    InMux I__16283 (
            .O(N__72486),
            .I(N__72482));
    CascadeMux I__16282 (
            .O(N__72485),
            .I(N__72478));
    LocalMux I__16281 (
            .O(N__72482),
            .I(N__72475));
    InMux I__16280 (
            .O(N__72481),
            .I(N__72472));
    InMux I__16279 (
            .O(N__72478),
            .I(N__72469));
    Span4Mux_v I__16278 (
            .O(N__72475),
            .I(N__72466));
    LocalMux I__16277 (
            .O(N__72472),
            .I(N__72463));
    LocalMux I__16276 (
            .O(N__72469),
            .I(N__72460));
    Odrv4 I__16275 (
            .O(N__72466),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_0_c_RNITGKN ));
    Odrv4 I__16274 (
            .O(N__72463),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_0_c_RNITGKN ));
    Odrv4 I__16273 (
            .O(N__72460),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_0_c_RNITGKN ));
    InMux I__16272 (
            .O(N__72453),
            .I(N__72450));
    LocalMux I__16271 (
            .O(N__72450),
            .I(\pid_side.error_d_reg_prev_esr_RNIM6H42Z0Z_0 ));
    InMux I__16270 (
            .O(N__72447),
            .I(N__72444));
    LocalMux I__16269 (
            .O(N__72444),
            .I(N__72441));
    Odrv4 I__16268 (
            .O(N__72441),
            .I(\pid_front.error_i_reg_9_sn_17 ));
    CascadeMux I__16267 (
            .O(N__72438),
            .I(\pid_front.error_i_reg_9_rn_1_17_cascade_ ));
    InMux I__16266 (
            .O(N__72435),
            .I(N__72432));
    LocalMux I__16265 (
            .O(N__72432),
            .I(N__72429));
    Span4Mux_h I__16264 (
            .O(N__72429),
            .I(N__72426));
    Odrv4 I__16263 (
            .O(N__72426),
            .I(\pid_front.error_i_regZ0Z_17 ));
    CEMux I__16262 (
            .O(N__72423),
            .I(N__72419));
    CEMux I__16261 (
            .O(N__72422),
            .I(N__72409));
    LocalMux I__16260 (
            .O(N__72419),
            .I(N__72403));
    CEMux I__16259 (
            .O(N__72418),
            .I(N__72400));
    CEMux I__16258 (
            .O(N__72417),
            .I(N__72397));
    CEMux I__16257 (
            .O(N__72416),
            .I(N__72394));
    CEMux I__16256 (
            .O(N__72415),
            .I(N__72391));
    CEMux I__16255 (
            .O(N__72414),
            .I(N__72387));
    CEMux I__16254 (
            .O(N__72413),
            .I(N__72384));
    CEMux I__16253 (
            .O(N__72412),
            .I(N__72381));
    LocalMux I__16252 (
            .O(N__72409),
            .I(N__72378));
    CEMux I__16251 (
            .O(N__72408),
            .I(N__72375));
    CEMux I__16250 (
            .O(N__72407),
            .I(N__72372));
    CEMux I__16249 (
            .O(N__72406),
            .I(N__72369));
    Span4Mux_h I__16248 (
            .O(N__72403),
            .I(N__72360));
    LocalMux I__16247 (
            .O(N__72400),
            .I(N__72360));
    LocalMux I__16246 (
            .O(N__72397),
            .I(N__72360));
    LocalMux I__16245 (
            .O(N__72394),
            .I(N__72360));
    LocalMux I__16244 (
            .O(N__72391),
            .I(N__72357));
    CEMux I__16243 (
            .O(N__72390),
            .I(N__72354));
    LocalMux I__16242 (
            .O(N__72387),
            .I(N__72350));
    LocalMux I__16241 (
            .O(N__72384),
            .I(N__72347));
    LocalMux I__16240 (
            .O(N__72381),
            .I(N__72342));
    Span4Mux_h I__16239 (
            .O(N__72378),
            .I(N__72342));
    LocalMux I__16238 (
            .O(N__72375),
            .I(N__72339));
    LocalMux I__16237 (
            .O(N__72372),
            .I(N__72336));
    LocalMux I__16236 (
            .O(N__72369),
            .I(N__72331));
    Span4Mux_v I__16235 (
            .O(N__72360),
            .I(N__72331));
    Span4Mux_v I__16234 (
            .O(N__72357),
            .I(N__72326));
    LocalMux I__16233 (
            .O(N__72354),
            .I(N__72326));
    CEMux I__16232 (
            .O(N__72353),
            .I(N__72323));
    Span4Mux_h I__16231 (
            .O(N__72350),
            .I(N__72320));
    Span4Mux_h I__16230 (
            .O(N__72347),
            .I(N__72317));
    Span4Mux_h I__16229 (
            .O(N__72342),
            .I(N__72314));
    Span4Mux_v I__16228 (
            .O(N__72339),
            .I(N__72311));
    Span4Mux_h I__16227 (
            .O(N__72336),
            .I(N__72308));
    Span4Mux_h I__16226 (
            .O(N__72331),
            .I(N__72303));
    Span4Mux_h I__16225 (
            .O(N__72326),
            .I(N__72303));
    LocalMux I__16224 (
            .O(N__72323),
            .I(N__72300));
    Span4Mux_h I__16223 (
            .O(N__72320),
            .I(N__72297));
    Span4Mux_h I__16222 (
            .O(N__72317),
            .I(N__72292));
    Span4Mux_h I__16221 (
            .O(N__72314),
            .I(N__72292));
    Span4Mux_h I__16220 (
            .O(N__72311),
            .I(N__72289));
    Span4Mux_h I__16219 (
            .O(N__72308),
            .I(N__72284));
    Span4Mux_h I__16218 (
            .O(N__72303),
            .I(N__72284));
    Odrv12 I__16217 (
            .O(N__72300),
            .I(\pid_front.state_ns_0_0 ));
    Odrv4 I__16216 (
            .O(N__72297),
            .I(\pid_front.state_ns_0_0 ));
    Odrv4 I__16215 (
            .O(N__72292),
            .I(\pid_front.state_ns_0_0 ));
    Odrv4 I__16214 (
            .O(N__72289),
            .I(\pid_front.state_ns_0_0 ));
    Odrv4 I__16213 (
            .O(N__72284),
            .I(\pid_front.state_ns_0_0 ));
    InMux I__16212 (
            .O(N__72273),
            .I(N__72270));
    LocalMux I__16211 (
            .O(N__72270),
            .I(\pid_front.error_i_reg_esr_RNO_4_0_17 ));
    InMux I__16210 (
            .O(N__72267),
            .I(N__72264));
    LocalMux I__16209 (
            .O(N__72264),
            .I(N__72259));
    InMux I__16208 (
            .O(N__72263),
            .I(N__72254));
    InMux I__16207 (
            .O(N__72262),
            .I(N__72254));
    Span4Mux_v I__16206 (
            .O(N__72259),
            .I(N__72251));
    LocalMux I__16205 (
            .O(N__72254),
            .I(N__72248));
    Span4Mux_h I__16204 (
            .O(N__72251),
            .I(N__72245));
    Span4Mux_h I__16203 (
            .O(N__72248),
            .I(N__72242));
    Odrv4 I__16202 (
            .O(N__72245),
            .I(\pid_front.N_51_1 ));
    Odrv4 I__16201 (
            .O(N__72242),
            .I(\pid_front.N_51_1 ));
    InMux I__16200 (
            .O(N__72237),
            .I(N__72233));
    InMux I__16199 (
            .O(N__72236),
            .I(N__72230));
    LocalMux I__16198 (
            .O(N__72233),
            .I(N__72227));
    LocalMux I__16197 (
            .O(N__72230),
            .I(N__72224));
    Span4Mux_h I__16196 (
            .O(N__72227),
            .I(N__72218));
    Span4Mux_h I__16195 (
            .O(N__72224),
            .I(N__72218));
    InMux I__16194 (
            .O(N__72223),
            .I(N__72215));
    Odrv4 I__16193 (
            .O(N__72218),
            .I(\pid_front.N_48_1 ));
    LocalMux I__16192 (
            .O(N__72215),
            .I(\pid_front.N_48_1 ));
    InMux I__16191 (
            .O(N__72210),
            .I(N__72207));
    LocalMux I__16190 (
            .O(N__72207),
            .I(N__72204));
    Span4Mux_v I__16189 (
            .O(N__72204),
            .I(N__72200));
    InMux I__16188 (
            .O(N__72203),
            .I(N__72197));
    Odrv4 I__16187 (
            .O(N__72200),
            .I(\pid_front.N_47_1 ));
    LocalMux I__16186 (
            .O(N__72197),
            .I(\pid_front.N_47_1 ));
    CascadeMux I__16185 (
            .O(N__72192),
            .I(\pid_front.m89_0_ns_1_cascade_ ));
    InMux I__16184 (
            .O(N__72189),
            .I(N__72186));
    LocalMux I__16183 (
            .O(N__72186),
            .I(N__72182));
    InMux I__16182 (
            .O(N__72185),
            .I(N__72179));
    Span4Mux_v I__16181 (
            .O(N__72182),
            .I(N__72174));
    LocalMux I__16180 (
            .O(N__72179),
            .I(N__72174));
    Span4Mux_h I__16179 (
            .O(N__72174),
            .I(N__72171));
    Odrv4 I__16178 (
            .O(N__72171),
            .I(\pid_front.N_45_1 ));
    InMux I__16177 (
            .O(N__72168),
            .I(N__72161));
    InMux I__16176 (
            .O(N__72167),
            .I(N__72161));
    InMux I__16175 (
            .O(N__72166),
            .I(N__72158));
    LocalMux I__16174 (
            .O(N__72161),
            .I(\pid_front.N_90_0 ));
    LocalMux I__16173 (
            .O(N__72158),
            .I(\pid_front.N_90_0 ));
    InMux I__16172 (
            .O(N__72153),
            .I(N__72149));
    InMux I__16171 (
            .O(N__72152),
            .I(N__72146));
    LocalMux I__16170 (
            .O(N__72149),
            .I(N__72143));
    LocalMux I__16169 (
            .O(N__72146),
            .I(N__72140));
    Span4Mux_v I__16168 (
            .O(N__72143),
            .I(N__72137));
    Span4Mux_v I__16167 (
            .O(N__72140),
            .I(N__72134));
    Span4Mux_h I__16166 (
            .O(N__72137),
            .I(N__72127));
    Span4Mux_h I__16165 (
            .O(N__72134),
            .I(N__72124));
    InMux I__16164 (
            .O(N__72133),
            .I(N__72121));
    InMux I__16163 (
            .O(N__72132),
            .I(N__72117));
    InMux I__16162 (
            .O(N__72131),
            .I(N__72112));
    InMux I__16161 (
            .O(N__72130),
            .I(N__72112));
    Span4Mux_h I__16160 (
            .O(N__72127),
            .I(N__72107));
    Span4Mux_h I__16159 (
            .O(N__72124),
            .I(N__72102));
    LocalMux I__16158 (
            .O(N__72121),
            .I(N__72102));
    InMux I__16157 (
            .O(N__72120),
            .I(N__72099));
    LocalMux I__16156 (
            .O(N__72117),
            .I(N__72094));
    LocalMux I__16155 (
            .O(N__72112),
            .I(N__72094));
    InMux I__16154 (
            .O(N__72111),
            .I(N__72088));
    InMux I__16153 (
            .O(N__72110),
            .I(N__72088));
    Span4Mux_h I__16152 (
            .O(N__72107),
            .I(N__72083));
    Span4Mux_h I__16151 (
            .O(N__72102),
            .I(N__72083));
    LocalMux I__16150 (
            .O(N__72099),
            .I(N__72078));
    Span4Mux_h I__16149 (
            .O(N__72094),
            .I(N__72078));
    InMux I__16148 (
            .O(N__72093),
            .I(N__72075));
    LocalMux I__16147 (
            .O(N__72088),
            .I(N__72072));
    Odrv4 I__16146 (
            .O(N__72083),
            .I(\pid_front.error_14 ));
    Odrv4 I__16145 (
            .O(N__72078),
            .I(\pid_front.error_14 ));
    LocalMux I__16144 (
            .O(N__72075),
            .I(\pid_front.error_14 ));
    Odrv12 I__16143 (
            .O(N__72072),
            .I(\pid_front.error_14 ));
    CascadeMux I__16142 (
            .O(N__72063),
            .I(N__72058));
    CascadeMux I__16141 (
            .O(N__72062),
            .I(N__72054));
    CascadeMux I__16140 (
            .O(N__72061),
            .I(N__72047));
    InMux I__16139 (
            .O(N__72058),
            .I(N__72041));
    CascadeMux I__16138 (
            .O(N__72057),
            .I(N__72033));
    InMux I__16137 (
            .O(N__72054),
            .I(N__72027));
    InMux I__16136 (
            .O(N__72053),
            .I(N__72027));
    InMux I__16135 (
            .O(N__72052),
            .I(N__72022));
    InMux I__16134 (
            .O(N__72051),
            .I(N__72022));
    InMux I__16133 (
            .O(N__72050),
            .I(N__72017));
    InMux I__16132 (
            .O(N__72047),
            .I(N__72017));
    InMux I__16131 (
            .O(N__72046),
            .I(N__72012));
    InMux I__16130 (
            .O(N__72045),
            .I(N__72012));
    InMux I__16129 (
            .O(N__72044),
            .I(N__72009));
    LocalMux I__16128 (
            .O(N__72041),
            .I(N__72005));
    InMux I__16127 (
            .O(N__72040),
            .I(N__72002));
    InMux I__16126 (
            .O(N__72039),
            .I(N__71997));
    InMux I__16125 (
            .O(N__72038),
            .I(N__71997));
    InMux I__16124 (
            .O(N__72037),
            .I(N__71992));
    InMux I__16123 (
            .O(N__72036),
            .I(N__71992));
    InMux I__16122 (
            .O(N__72033),
            .I(N__71989));
    CascadeMux I__16121 (
            .O(N__72032),
            .I(N__71984));
    LocalMux I__16120 (
            .O(N__72027),
            .I(N__71981));
    LocalMux I__16119 (
            .O(N__72022),
            .I(N__71978));
    LocalMux I__16118 (
            .O(N__72017),
            .I(N__71975));
    LocalMux I__16117 (
            .O(N__72012),
            .I(N__71971));
    LocalMux I__16116 (
            .O(N__72009),
            .I(N__71963));
    InMux I__16115 (
            .O(N__72008),
            .I(N__71960));
    Span4Mux_h I__16114 (
            .O(N__72005),
            .I(N__71953));
    LocalMux I__16113 (
            .O(N__72002),
            .I(N__71953));
    LocalMux I__16112 (
            .O(N__71997),
            .I(N__71953));
    LocalMux I__16111 (
            .O(N__71992),
            .I(N__71950));
    LocalMux I__16110 (
            .O(N__71989),
            .I(N__71947));
    InMux I__16109 (
            .O(N__71988),
            .I(N__71944));
    InMux I__16108 (
            .O(N__71987),
            .I(N__71939));
    InMux I__16107 (
            .O(N__71984),
            .I(N__71939));
    Span4Mux_v I__16106 (
            .O(N__71981),
            .I(N__71936));
    Span4Mux_v I__16105 (
            .O(N__71978),
            .I(N__71931));
    Span4Mux_h I__16104 (
            .O(N__71975),
            .I(N__71931));
    InMux I__16103 (
            .O(N__71974),
            .I(N__71928));
    Span4Mux_h I__16102 (
            .O(N__71971),
            .I(N__71925));
    InMux I__16101 (
            .O(N__71970),
            .I(N__71922));
    InMux I__16100 (
            .O(N__71969),
            .I(N__71917));
    InMux I__16099 (
            .O(N__71968),
            .I(N__71917));
    InMux I__16098 (
            .O(N__71967),
            .I(N__71912));
    InMux I__16097 (
            .O(N__71966),
            .I(N__71912));
    Span4Mux_h I__16096 (
            .O(N__71963),
            .I(N__71903));
    LocalMux I__16095 (
            .O(N__71960),
            .I(N__71903));
    Span4Mux_v I__16094 (
            .O(N__71953),
            .I(N__71903));
    Span4Mux_h I__16093 (
            .O(N__71950),
            .I(N__71903));
    Span4Mux_h I__16092 (
            .O(N__71947),
            .I(N__71896));
    LocalMux I__16091 (
            .O(N__71944),
            .I(N__71896));
    LocalMux I__16090 (
            .O(N__71939),
            .I(N__71896));
    Span4Mux_h I__16089 (
            .O(N__71936),
            .I(N__71891));
    Span4Mux_v I__16088 (
            .O(N__71931),
            .I(N__71891));
    LocalMux I__16087 (
            .O(N__71928),
            .I(xy_ki_1));
    Odrv4 I__16086 (
            .O(N__71925),
            .I(xy_ki_1));
    LocalMux I__16085 (
            .O(N__71922),
            .I(xy_ki_1));
    LocalMux I__16084 (
            .O(N__71917),
            .I(xy_ki_1));
    LocalMux I__16083 (
            .O(N__71912),
            .I(xy_ki_1));
    Odrv4 I__16082 (
            .O(N__71903),
            .I(xy_ki_1));
    Odrv4 I__16081 (
            .O(N__71896),
            .I(xy_ki_1));
    Odrv4 I__16080 (
            .O(N__71891),
            .I(xy_ki_1));
    InMux I__16079 (
            .O(N__71874),
            .I(N__71871));
    LocalMux I__16078 (
            .O(N__71871),
            .I(\pid_front.error_i_reg_esr_RNO_5_0_17 ));
    InMux I__16077 (
            .O(N__71868),
            .I(N__71865));
    LocalMux I__16076 (
            .O(N__71865),
            .I(N__71862));
    Span4Mux_h I__16075 (
            .O(N__71862),
            .I(N__71859));
    Span4Mux_v I__16074 (
            .O(N__71859),
            .I(N__71856));
    Span4Mux_h I__16073 (
            .O(N__71856),
            .I(N__71853));
    Odrv4 I__16072 (
            .O(N__71853),
            .I(\pid_alt.state_RNIFCSD1Z0Z_0 ));
    IoInMux I__16071 (
            .O(N__71850),
            .I(N__71847));
    LocalMux I__16070 (
            .O(N__71847),
            .I(N__71844));
    Span4Mux_s3_v I__16069 (
            .O(N__71844),
            .I(N__71841));
    Odrv4 I__16068 (
            .O(N__71841),
            .I(\pid_alt.N_939_0 ));
    InMux I__16067 (
            .O(N__71838),
            .I(N__71834));
    InMux I__16066 (
            .O(N__71837),
            .I(N__71830));
    LocalMux I__16065 (
            .O(N__71834),
            .I(N__71827));
    InMux I__16064 (
            .O(N__71833),
            .I(N__71824));
    LocalMux I__16063 (
            .O(N__71830),
            .I(N__71821));
    Span4Mux_h I__16062 (
            .O(N__71827),
            .I(N__71818));
    LocalMux I__16061 (
            .O(N__71824),
            .I(N__71815));
    Span4Mux_h I__16060 (
            .O(N__71821),
            .I(N__71810));
    Span4Mux_v I__16059 (
            .O(N__71818),
            .I(N__71810));
    Odrv4 I__16058 (
            .O(N__71815),
            .I(\pid_side.pid_preregZ0Z_10 ));
    Odrv4 I__16057 (
            .O(N__71810),
            .I(\pid_side.pid_preregZ0Z_10 ));
    InMux I__16056 (
            .O(N__71805),
            .I(N__71801));
    CascadeMux I__16055 (
            .O(N__71804),
            .I(N__71798));
    LocalMux I__16054 (
            .O(N__71801),
            .I(N__71794));
    InMux I__16053 (
            .O(N__71798),
            .I(N__71791));
    InMux I__16052 (
            .O(N__71797),
            .I(N__71788));
    Span4Mux_v I__16051 (
            .O(N__71794),
            .I(N__71783));
    LocalMux I__16050 (
            .O(N__71791),
            .I(N__71783));
    LocalMux I__16049 (
            .O(N__71788),
            .I(N__71780));
    Span4Mux_h I__16048 (
            .O(N__71783),
            .I(N__71777));
    Odrv4 I__16047 (
            .O(N__71780),
            .I(\pid_side.pid_preregZ0Z_7 ));
    Odrv4 I__16046 (
            .O(N__71777),
            .I(\pid_side.pid_preregZ0Z_7 ));
    CascadeMux I__16045 (
            .O(N__71772),
            .I(N__71768));
    InMux I__16044 (
            .O(N__71771),
            .I(N__71764));
    InMux I__16043 (
            .O(N__71768),
            .I(N__71761));
    CascadeMux I__16042 (
            .O(N__71767),
            .I(N__71758));
    LocalMux I__16041 (
            .O(N__71764),
            .I(N__71755));
    LocalMux I__16040 (
            .O(N__71761),
            .I(N__71752));
    InMux I__16039 (
            .O(N__71758),
            .I(N__71749));
    Span4Mux_v I__16038 (
            .O(N__71755),
            .I(N__71744));
    Span4Mux_v I__16037 (
            .O(N__71752),
            .I(N__71744));
    LocalMux I__16036 (
            .O(N__71749),
            .I(N__71741));
    Span4Mux_h I__16035 (
            .O(N__71744),
            .I(N__71738));
    Odrv4 I__16034 (
            .O(N__71741),
            .I(\pid_side.pid_preregZ0Z_11 ));
    Odrv4 I__16033 (
            .O(N__71738),
            .I(\pid_side.pid_preregZ0Z_11 ));
    InMux I__16032 (
            .O(N__71733),
            .I(N__71727));
    InMux I__16031 (
            .O(N__71732),
            .I(N__71727));
    LocalMux I__16030 (
            .O(N__71727),
            .I(N__71723));
    InMux I__16029 (
            .O(N__71726),
            .I(N__71720));
    Span4Mux_h I__16028 (
            .O(N__71723),
            .I(N__71717));
    LocalMux I__16027 (
            .O(N__71720),
            .I(\pid_side.pid_preregZ0Z_6 ));
    Odrv4 I__16026 (
            .O(N__71717),
            .I(\pid_side.pid_preregZ0Z_6 ));
    InMux I__16025 (
            .O(N__71712),
            .I(N__71705));
    InMux I__16024 (
            .O(N__71711),
            .I(N__71702));
    InMux I__16023 (
            .O(N__71710),
            .I(N__71694));
    InMux I__16022 (
            .O(N__71709),
            .I(N__71694));
    InMux I__16021 (
            .O(N__71708),
            .I(N__71694));
    LocalMux I__16020 (
            .O(N__71705),
            .I(N__71689));
    LocalMux I__16019 (
            .O(N__71702),
            .I(N__71689));
    InMux I__16018 (
            .O(N__71701),
            .I(N__71686));
    LocalMux I__16017 (
            .O(N__71694),
            .I(N__71683));
    Span4Mux_h I__16016 (
            .O(N__71689),
            .I(N__71678));
    LocalMux I__16015 (
            .O(N__71686),
            .I(N__71678));
    Span4Mux_h I__16014 (
            .O(N__71683),
            .I(N__71675));
    Odrv4 I__16013 (
            .O(N__71678),
            .I(\pid_side.pid_preregZ0Z_13 ));
    Odrv4 I__16012 (
            .O(N__71675),
            .I(\pid_side.pid_preregZ0Z_13 ));
    InMux I__16011 (
            .O(N__71670),
            .I(N__71666));
    InMux I__16010 (
            .O(N__71669),
            .I(N__71663));
    LocalMux I__16009 (
            .O(N__71666),
            .I(N__71659));
    LocalMux I__16008 (
            .O(N__71663),
            .I(N__71656));
    InMux I__16007 (
            .O(N__71662),
            .I(N__71653));
    Span4Mux_h I__16006 (
            .O(N__71659),
            .I(N__71650));
    Span4Mux_v I__16005 (
            .O(N__71656),
            .I(N__71647));
    LocalMux I__16004 (
            .O(N__71653),
            .I(N__71644));
    Span4Mux_v I__16003 (
            .O(N__71650),
            .I(N__71641));
    Odrv4 I__16002 (
            .O(N__71647),
            .I(\pid_side.pid_preregZ0Z_9 ));
    Odrv4 I__16001 (
            .O(N__71644),
            .I(\pid_side.pid_preregZ0Z_9 ));
    Odrv4 I__16000 (
            .O(N__71641),
            .I(\pid_side.pid_preregZ0Z_9 ));
    CascadeMux I__15999 (
            .O(N__71634),
            .I(\pid_side.source_pid_1_sqmuxa_1_0_a2_1_4_cascade_ ));
    InMux I__15998 (
            .O(N__71631),
            .I(N__71627));
    InMux I__15997 (
            .O(N__71630),
            .I(N__71624));
    LocalMux I__15996 (
            .O(N__71627),
            .I(N__71620));
    LocalMux I__15995 (
            .O(N__71624),
            .I(N__71617));
    InMux I__15994 (
            .O(N__71623),
            .I(N__71614));
    Span4Mux_h I__15993 (
            .O(N__71620),
            .I(N__71611));
    Span4Mux_h I__15992 (
            .O(N__71617),
            .I(N__71608));
    LocalMux I__15991 (
            .O(N__71614),
            .I(N__71605));
    Span4Mux_v I__15990 (
            .O(N__71611),
            .I(N__71602));
    Odrv4 I__15989 (
            .O(N__71608),
            .I(\pid_side.pid_preregZ0Z_8 ));
    Odrv4 I__15988 (
            .O(N__71605),
            .I(\pid_side.pid_preregZ0Z_8 ));
    Odrv4 I__15987 (
            .O(N__71602),
            .I(\pid_side.pid_preregZ0Z_8 ));
    InMux I__15986 (
            .O(N__71595),
            .I(N__71592));
    LocalMux I__15985 (
            .O(N__71592),
            .I(N__71587));
    InMux I__15984 (
            .O(N__71591),
            .I(N__71584));
    InMux I__15983 (
            .O(N__71590),
            .I(N__71581));
    Span4Mux_h I__15982 (
            .O(N__71587),
            .I(N__71578));
    LocalMux I__15981 (
            .O(N__71584),
            .I(N__71573));
    LocalMux I__15980 (
            .O(N__71581),
            .I(N__71573));
    Span4Mux_h I__15979 (
            .O(N__71578),
            .I(N__71570));
    Span4Mux_v I__15978 (
            .O(N__71573),
            .I(N__71567));
    Odrv4 I__15977 (
            .O(N__71570),
            .I(\pid_side.N_99 ));
    Odrv4 I__15976 (
            .O(N__71567),
            .I(\pid_side.N_99 ));
    CascadeMux I__15975 (
            .O(N__71562),
            .I(N__71553));
    InMux I__15974 (
            .O(N__71561),
            .I(N__71537));
    InMux I__15973 (
            .O(N__71560),
            .I(N__71537));
    InMux I__15972 (
            .O(N__71559),
            .I(N__71537));
    InMux I__15971 (
            .O(N__71558),
            .I(N__71532));
    InMux I__15970 (
            .O(N__71557),
            .I(N__71532));
    InMux I__15969 (
            .O(N__71556),
            .I(N__71527));
    InMux I__15968 (
            .O(N__71553),
            .I(N__71520));
    InMux I__15967 (
            .O(N__71552),
            .I(N__71520));
    CascadeMux I__15966 (
            .O(N__71551),
            .I(N__71513));
    CascadeMux I__15965 (
            .O(N__71550),
            .I(N__71510));
    InMux I__15964 (
            .O(N__71549),
            .I(N__71506));
    InMux I__15963 (
            .O(N__71548),
            .I(N__71503));
    InMux I__15962 (
            .O(N__71547),
            .I(N__71498));
    InMux I__15961 (
            .O(N__71546),
            .I(N__71495));
    InMux I__15960 (
            .O(N__71545),
            .I(N__71490));
    InMux I__15959 (
            .O(N__71544),
            .I(N__71490));
    LocalMux I__15958 (
            .O(N__71537),
            .I(N__71485));
    LocalMux I__15957 (
            .O(N__71532),
            .I(N__71485));
    CascadeMux I__15956 (
            .O(N__71531),
            .I(N__71482));
    InMux I__15955 (
            .O(N__71530),
            .I(N__71477));
    LocalMux I__15954 (
            .O(N__71527),
            .I(N__71474));
    InMux I__15953 (
            .O(N__71526),
            .I(N__71469));
    InMux I__15952 (
            .O(N__71525),
            .I(N__71469));
    LocalMux I__15951 (
            .O(N__71520),
            .I(N__71466));
    InMux I__15950 (
            .O(N__71519),
            .I(N__71461));
    InMux I__15949 (
            .O(N__71518),
            .I(N__71461));
    InMux I__15948 (
            .O(N__71517),
            .I(N__71455));
    InMux I__15947 (
            .O(N__71516),
            .I(N__71455));
    InMux I__15946 (
            .O(N__71513),
            .I(N__71450));
    InMux I__15945 (
            .O(N__71510),
            .I(N__71450));
    InMux I__15944 (
            .O(N__71509),
            .I(N__71447));
    LocalMux I__15943 (
            .O(N__71506),
            .I(N__71444));
    LocalMux I__15942 (
            .O(N__71503),
            .I(N__71441));
    InMux I__15941 (
            .O(N__71502),
            .I(N__71438));
    InMux I__15940 (
            .O(N__71501),
            .I(N__71435));
    LocalMux I__15939 (
            .O(N__71498),
            .I(N__71428));
    LocalMux I__15938 (
            .O(N__71495),
            .I(N__71428));
    LocalMux I__15937 (
            .O(N__71490),
            .I(N__71428));
    Span4Mux_v I__15936 (
            .O(N__71485),
            .I(N__71425));
    InMux I__15935 (
            .O(N__71482),
            .I(N__71418));
    InMux I__15934 (
            .O(N__71481),
            .I(N__71418));
    InMux I__15933 (
            .O(N__71480),
            .I(N__71418));
    LocalMux I__15932 (
            .O(N__71477),
            .I(N__71415));
    Span4Mux_h I__15931 (
            .O(N__71474),
            .I(N__71412));
    LocalMux I__15930 (
            .O(N__71469),
            .I(N__71407));
    Span4Mux_h I__15929 (
            .O(N__71466),
            .I(N__71407));
    LocalMux I__15928 (
            .O(N__71461),
            .I(N__71404));
    InMux I__15927 (
            .O(N__71460),
            .I(N__71401));
    LocalMux I__15926 (
            .O(N__71455),
            .I(N__71396));
    LocalMux I__15925 (
            .O(N__71450),
            .I(N__71396));
    LocalMux I__15924 (
            .O(N__71447),
            .I(N__71393));
    Span4Mux_h I__15923 (
            .O(N__71444),
            .I(N__71390));
    Span4Mux_h I__15922 (
            .O(N__71441),
            .I(N__71387));
    LocalMux I__15921 (
            .O(N__71438),
            .I(N__71380));
    LocalMux I__15920 (
            .O(N__71435),
            .I(N__71380));
    Span4Mux_v I__15919 (
            .O(N__71428),
            .I(N__71380));
    Span4Mux_h I__15918 (
            .O(N__71425),
            .I(N__71375));
    LocalMux I__15917 (
            .O(N__71418),
            .I(N__71375));
    Span4Mux_v I__15916 (
            .O(N__71415),
            .I(N__71368));
    Span4Mux_v I__15915 (
            .O(N__71412),
            .I(N__71368));
    Span4Mux_v I__15914 (
            .O(N__71407),
            .I(N__71368));
    Span4Mux_v I__15913 (
            .O(N__71404),
            .I(N__71363));
    LocalMux I__15912 (
            .O(N__71401),
            .I(N__71363));
    Span4Mux_v I__15911 (
            .O(N__71396),
            .I(N__71358));
    Span4Mux_h I__15910 (
            .O(N__71393),
            .I(N__71358));
    Span4Mux_h I__15909 (
            .O(N__71390),
            .I(N__71355));
    Span4Mux_v I__15908 (
            .O(N__71387),
            .I(N__71350));
    Span4Mux_v I__15907 (
            .O(N__71380),
            .I(N__71350));
    Span4Mux_h I__15906 (
            .O(N__71375),
            .I(N__71345));
    Span4Mux_h I__15905 (
            .O(N__71368),
            .I(N__71345));
    Span4Mux_h I__15904 (
            .O(N__71363),
            .I(N__71340));
    Span4Mux_h I__15903 (
            .O(N__71358),
            .I(N__71340));
    Odrv4 I__15902 (
            .O(N__71355),
            .I(xy_ki_2));
    Odrv4 I__15901 (
            .O(N__71350),
            .I(xy_ki_2));
    Odrv4 I__15900 (
            .O(N__71345),
            .I(xy_ki_2));
    Odrv4 I__15899 (
            .O(N__71340),
            .I(xy_ki_2));
    CascadeMux I__15898 (
            .O(N__71331),
            .I(\pid_front.error_i_reg_esr_RNO_0_0_23_cascade_ ));
    InMux I__15897 (
            .O(N__71328),
            .I(N__71325));
    LocalMux I__15896 (
            .O(N__71325),
            .I(N__71322));
    Span4Mux_h I__15895 (
            .O(N__71322),
            .I(N__71319));
    Odrv4 I__15894 (
            .O(N__71319),
            .I(\pid_front.error_i_regZ0Z_23 ));
    CascadeMux I__15893 (
            .O(N__71316),
            .I(\pid_front.error_cry_9_c_RNICELJ1Z0Z_0_cascade_ ));
    InMux I__15892 (
            .O(N__71313),
            .I(N__71310));
    LocalMux I__15891 (
            .O(N__71310),
            .I(\pid_front.error_cry_9_c_RNICELJZ0Z1 ));
    InMux I__15890 (
            .O(N__71307),
            .I(N__71301));
    InMux I__15889 (
            .O(N__71306),
            .I(N__71298));
    InMux I__15888 (
            .O(N__71305),
            .I(N__71293));
    InMux I__15887 (
            .O(N__71304),
            .I(N__71293));
    LocalMux I__15886 (
            .O(N__71301),
            .I(\pid_front.N_46_1 ));
    LocalMux I__15885 (
            .O(N__71298),
            .I(\pid_front.N_46_1 ));
    LocalMux I__15884 (
            .O(N__71293),
            .I(\pid_front.N_46_1 ));
    InMux I__15883 (
            .O(N__71286),
            .I(N__71283));
    LocalMux I__15882 (
            .O(N__71283),
            .I(N__71278));
    InMux I__15881 (
            .O(N__71282),
            .I(N__71275));
    InMux I__15880 (
            .O(N__71281),
            .I(N__71272));
    Span4Mux_v I__15879 (
            .O(N__71278),
            .I(N__71266));
    LocalMux I__15878 (
            .O(N__71275),
            .I(N__71266));
    LocalMux I__15877 (
            .O(N__71272),
            .I(N__71262));
    InMux I__15876 (
            .O(N__71271),
            .I(N__71259));
    Span4Mux_v I__15875 (
            .O(N__71266),
            .I(N__71256));
    InMux I__15874 (
            .O(N__71265),
            .I(N__71253));
    Span4Mux_v I__15873 (
            .O(N__71262),
            .I(N__71246));
    LocalMux I__15872 (
            .O(N__71259),
            .I(N__71246));
    Span4Mux_v I__15871 (
            .O(N__71256),
            .I(N__71246));
    LocalMux I__15870 (
            .O(N__71253),
            .I(N__71243));
    Odrv4 I__15869 (
            .O(N__71246),
            .I(pid_front_error_i_reg_9_sn_19));
    Odrv4 I__15868 (
            .O(N__71243),
            .I(pid_front_error_i_reg_9_sn_19));
    CascadeMux I__15867 (
            .O(N__71238),
            .I(\pid_front.N_46_1_cascade_ ));
    InMux I__15866 (
            .O(N__71235),
            .I(N__71232));
    LocalMux I__15865 (
            .O(N__71232),
            .I(\pid_front.error_i_reg_esr_RNO_1Z0Z_19 ));
    InMux I__15864 (
            .O(N__71229),
            .I(N__71226));
    LocalMux I__15863 (
            .O(N__71226),
            .I(N__71223));
    Odrv12 I__15862 (
            .O(N__71223),
            .I(\pid_front.O_5 ));
    InMux I__15861 (
            .O(N__71220),
            .I(N__71211));
    InMux I__15860 (
            .O(N__71219),
            .I(N__71211));
    InMux I__15859 (
            .O(N__71218),
            .I(N__71211));
    LocalMux I__15858 (
            .O(N__71211),
            .I(N__71208));
    Span4Mux_v I__15857 (
            .O(N__71208),
            .I(N__71205));
    Span4Mux_h I__15856 (
            .O(N__71205),
            .I(N__71202));
    Odrv4 I__15855 (
            .O(N__71202),
            .I(\pid_front.error_d_regZ0Z_3 ));
    InMux I__15854 (
            .O(N__71199),
            .I(N__71195));
    InMux I__15853 (
            .O(N__71198),
            .I(N__71192));
    LocalMux I__15852 (
            .O(N__71195),
            .I(N__71189));
    LocalMux I__15851 (
            .O(N__71192),
            .I(N__71185));
    Span4Mux_v I__15850 (
            .O(N__71189),
            .I(N__71180));
    InMux I__15849 (
            .O(N__71188),
            .I(N__71176));
    Span4Mux_v I__15848 (
            .O(N__71185),
            .I(N__71171));
    InMux I__15847 (
            .O(N__71184),
            .I(N__71162));
    InMux I__15846 (
            .O(N__71183),
            .I(N__71162));
    Span4Mux_h I__15845 (
            .O(N__71180),
            .I(N__71159));
    InMux I__15844 (
            .O(N__71179),
            .I(N__71156));
    LocalMux I__15843 (
            .O(N__71176),
            .I(N__71153));
    InMux I__15842 (
            .O(N__71175),
            .I(N__71148));
    InMux I__15841 (
            .O(N__71174),
            .I(N__71148));
    Span4Mux_h I__15840 (
            .O(N__71171),
            .I(N__71145));
    InMux I__15839 (
            .O(N__71170),
            .I(N__71140));
    InMux I__15838 (
            .O(N__71169),
            .I(N__71140));
    InMux I__15837 (
            .O(N__71168),
            .I(N__71137));
    InMux I__15836 (
            .O(N__71167),
            .I(N__71134));
    LocalMux I__15835 (
            .O(N__71162),
            .I(N__71125));
    Span4Mux_h I__15834 (
            .O(N__71159),
            .I(N__71113));
    LocalMux I__15833 (
            .O(N__71156),
            .I(N__71113));
    Span4Mux_v I__15832 (
            .O(N__71153),
            .I(N__71113));
    LocalMux I__15831 (
            .O(N__71148),
            .I(N__71113));
    Span4Mux_h I__15830 (
            .O(N__71145),
            .I(N__71110));
    LocalMux I__15829 (
            .O(N__71140),
            .I(N__71103));
    LocalMux I__15828 (
            .O(N__71137),
            .I(N__71103));
    LocalMux I__15827 (
            .O(N__71134),
            .I(N__71103));
    InMux I__15826 (
            .O(N__71133),
            .I(N__71098));
    InMux I__15825 (
            .O(N__71132),
            .I(N__71098));
    InMux I__15824 (
            .O(N__71131),
            .I(N__71089));
    InMux I__15823 (
            .O(N__71130),
            .I(N__71089));
    InMux I__15822 (
            .O(N__71129),
            .I(N__71089));
    InMux I__15821 (
            .O(N__71128),
            .I(N__71089));
    Span4Mux_h I__15820 (
            .O(N__71125),
            .I(N__71086));
    InMux I__15819 (
            .O(N__71124),
            .I(N__71079));
    InMux I__15818 (
            .O(N__71123),
            .I(N__71079));
    InMux I__15817 (
            .O(N__71122),
            .I(N__71079));
    Span4Mux_h I__15816 (
            .O(N__71113),
            .I(N__71076));
    Span4Mux_h I__15815 (
            .O(N__71110),
            .I(N__71071));
    Span4Mux_h I__15814 (
            .O(N__71103),
            .I(N__71071));
    LocalMux I__15813 (
            .O(N__71098),
            .I(N__71066));
    LocalMux I__15812 (
            .O(N__71089),
            .I(N__71066));
    Odrv4 I__15811 (
            .O(N__71086),
            .I(\pid_front.error_15 ));
    LocalMux I__15810 (
            .O(N__71079),
            .I(\pid_front.error_15 ));
    Odrv4 I__15809 (
            .O(N__71076),
            .I(\pid_front.error_15 ));
    Odrv4 I__15808 (
            .O(N__71071),
            .I(\pid_front.error_15 ));
    Odrv12 I__15807 (
            .O(N__71066),
            .I(\pid_front.error_15 ));
    CascadeMux I__15806 (
            .O(N__71055),
            .I(\pid_front.N_131_cascade_ ));
    InMux I__15805 (
            .O(N__71052),
            .I(N__71049));
    LocalMux I__15804 (
            .O(N__71049),
            .I(N__71046));
    Span4Mux_v I__15803 (
            .O(N__71046),
            .I(N__71043));
    Odrv4 I__15802 (
            .O(N__71043),
            .I(\pid_front.m5_2_03 ));
    CascadeMux I__15801 (
            .O(N__71040),
            .I(pid_side_N_166_mux_cascade_));
    InMux I__15800 (
            .O(N__71037),
            .I(N__71033));
    InMux I__15799 (
            .O(N__71036),
            .I(N__71030));
    LocalMux I__15798 (
            .O(N__71033),
            .I(pid_front_error_i_reg_9_rn_sn_15));
    LocalMux I__15797 (
            .O(N__71030),
            .I(pid_front_error_i_reg_9_rn_sn_15));
    CascadeMux I__15796 (
            .O(N__71025),
            .I(pid_front_error_i_reg_9_rn_sn_15_cascade_));
    InMux I__15795 (
            .O(N__71022),
            .I(N__71017));
    InMux I__15794 (
            .O(N__71021),
            .I(N__71013));
    InMux I__15793 (
            .O(N__71020),
            .I(N__71010));
    LocalMux I__15792 (
            .O(N__71017),
            .I(N__71007));
    InMux I__15791 (
            .O(N__71016),
            .I(N__71004));
    LocalMux I__15790 (
            .O(N__71013),
            .I(N__71001));
    LocalMux I__15789 (
            .O(N__71010),
            .I(N__70998));
    Span4Mux_v I__15788 (
            .O(N__71007),
            .I(N__70995));
    LocalMux I__15787 (
            .O(N__71004),
            .I(N__70992));
    Span4Mux_v I__15786 (
            .O(N__71001),
            .I(N__70989));
    Odrv4 I__15785 (
            .O(N__70998),
            .I(\pid_front.m1_0_03 ));
    Odrv4 I__15784 (
            .O(N__70995),
            .I(\pid_front.m1_0_03 ));
    Odrv12 I__15783 (
            .O(N__70992),
            .I(\pid_front.m1_0_03 ));
    Odrv4 I__15782 (
            .O(N__70989),
            .I(\pid_front.m1_0_03 ));
    CascadeMux I__15781 (
            .O(N__70980),
            .I(N__70974));
    CascadeMux I__15780 (
            .O(N__70979),
            .I(N__70970));
    InMux I__15779 (
            .O(N__70978),
            .I(N__70965));
    CascadeMux I__15778 (
            .O(N__70977),
            .I(N__70961));
    InMux I__15777 (
            .O(N__70974),
            .I(N__70958));
    CascadeMux I__15776 (
            .O(N__70973),
            .I(N__70954));
    InMux I__15775 (
            .O(N__70970),
            .I(N__70951));
    InMux I__15774 (
            .O(N__70969),
            .I(N__70946));
    InMux I__15773 (
            .O(N__70968),
            .I(N__70946));
    LocalMux I__15772 (
            .O(N__70965),
            .I(N__70943));
    InMux I__15771 (
            .O(N__70964),
            .I(N__70940));
    InMux I__15770 (
            .O(N__70961),
            .I(N__70937));
    LocalMux I__15769 (
            .O(N__70958),
            .I(N__70934));
    InMux I__15768 (
            .O(N__70957),
            .I(N__70929));
    InMux I__15767 (
            .O(N__70954),
            .I(N__70929));
    LocalMux I__15766 (
            .O(N__70951),
            .I(N__70923));
    LocalMux I__15765 (
            .O(N__70946),
            .I(N__70923));
    Span4Mux_v I__15764 (
            .O(N__70943),
            .I(N__70920));
    LocalMux I__15763 (
            .O(N__70940),
            .I(N__70915));
    LocalMux I__15762 (
            .O(N__70937),
            .I(N__70915));
    Span4Mux_v I__15761 (
            .O(N__70934),
            .I(N__70910));
    LocalMux I__15760 (
            .O(N__70929),
            .I(N__70910));
    CascadeMux I__15759 (
            .O(N__70928),
            .I(N__70907));
    Span4Mux_h I__15758 (
            .O(N__70923),
            .I(N__70904));
    Span4Mux_h I__15757 (
            .O(N__70920),
            .I(N__70899));
    Span4Mux_v I__15756 (
            .O(N__70915),
            .I(N__70894));
    Span4Mux_v I__15755 (
            .O(N__70910),
            .I(N__70894));
    InMux I__15754 (
            .O(N__70907),
            .I(N__70891));
    Span4Mux_v I__15753 (
            .O(N__70904),
            .I(N__70888));
    InMux I__15752 (
            .O(N__70903),
            .I(N__70885));
    InMux I__15751 (
            .O(N__70902),
            .I(N__70882));
    Odrv4 I__15750 (
            .O(N__70899),
            .I(pid_side_N_166_mux));
    Odrv4 I__15749 (
            .O(N__70894),
            .I(pid_side_N_166_mux));
    LocalMux I__15748 (
            .O(N__70891),
            .I(pid_side_N_166_mux));
    Odrv4 I__15747 (
            .O(N__70888),
            .I(pid_side_N_166_mux));
    LocalMux I__15746 (
            .O(N__70885),
            .I(pid_side_N_166_mux));
    LocalMux I__15745 (
            .O(N__70882),
            .I(pid_side_N_166_mux));
    InMux I__15744 (
            .O(N__70869),
            .I(N__70865));
    InMux I__15743 (
            .O(N__70868),
            .I(N__70862));
    LocalMux I__15742 (
            .O(N__70865),
            .I(N__70859));
    LocalMux I__15741 (
            .O(N__70862),
            .I(N__70854));
    Span4Mux_h I__15740 (
            .O(N__70859),
            .I(N__70851));
    InMux I__15739 (
            .O(N__70858),
            .I(N__70848));
    InMux I__15738 (
            .O(N__70857),
            .I(N__70845));
    Odrv4 I__15737 (
            .O(N__70854),
            .I(\pid_front.N_12_1 ));
    Odrv4 I__15736 (
            .O(N__70851),
            .I(\pid_front.N_12_1 ));
    LocalMux I__15735 (
            .O(N__70848),
            .I(\pid_front.N_12_1 ));
    LocalMux I__15734 (
            .O(N__70845),
            .I(\pid_front.N_12_1 ));
    CascadeMux I__15733 (
            .O(N__70836),
            .I(N__70833));
    InMux I__15732 (
            .O(N__70833),
            .I(N__70830));
    LocalMux I__15731 (
            .O(N__70830),
            .I(N__70827));
    Span4Mux_h I__15730 (
            .O(N__70827),
            .I(N__70824));
    Odrv4 I__15729 (
            .O(N__70824),
            .I(\pid_front.error_i_regZ0Z_1 ));
    InMux I__15728 (
            .O(N__70821),
            .I(N__70818));
    LocalMux I__15727 (
            .O(N__70818),
            .I(\pid_side.m1_2_03 ));
    InMux I__15726 (
            .O(N__70815),
            .I(N__70812));
    LocalMux I__15725 (
            .O(N__70812),
            .I(\pid_side.error_i_reg_9_rn_rn_2_13 ));
    CascadeMux I__15724 (
            .O(N__70809),
            .I(N__70806));
    InMux I__15723 (
            .O(N__70806),
            .I(N__70803));
    LocalMux I__15722 (
            .O(N__70803),
            .I(\pid_front.error_i_reg_esr_RNO_1Z0Z_15 ));
    InMux I__15721 (
            .O(N__70800),
            .I(N__70797));
    LocalMux I__15720 (
            .O(N__70797),
            .I(\pid_front.error_i_reg_esr_RNO_2Z0Z_15 ));
    CascadeMux I__15719 (
            .O(N__70794),
            .I(N__70791));
    InMux I__15718 (
            .O(N__70791),
            .I(N__70788));
    LocalMux I__15717 (
            .O(N__70788),
            .I(N__70785));
    Span4Mux_h I__15716 (
            .O(N__70785),
            .I(N__70782));
    Odrv4 I__15715 (
            .O(N__70782),
            .I(\pid_front.error_i_regZ0Z_15 ));
    InMux I__15714 (
            .O(N__70779),
            .I(N__70776));
    LocalMux I__15713 (
            .O(N__70776),
            .I(\pid_front.N_134 ));
    InMux I__15712 (
            .O(N__70773),
            .I(N__70770));
    LocalMux I__15711 (
            .O(N__70770),
            .I(N__70767));
    Span4Mux_v I__15710 (
            .O(N__70767),
            .I(N__70764));
    Odrv4 I__15709 (
            .O(N__70764),
            .I(\pid_side.N_48_1 ));
    CascadeMux I__15708 (
            .O(N__70761),
            .I(\pid_side.N_48_1_cascade_ ));
    InMux I__15707 (
            .O(N__70758),
            .I(N__70755));
    LocalMux I__15706 (
            .O(N__70755),
            .I(\pid_side.N_89_0 ));
    InMux I__15705 (
            .O(N__70752),
            .I(N__70749));
    LocalMux I__15704 (
            .O(N__70749),
            .I(\pid_side.N_126 ));
    InMux I__15703 (
            .O(N__70746),
            .I(N__70743));
    LocalMux I__15702 (
            .O(N__70743),
            .I(\pid_side.N_88_0 ));
    InMux I__15701 (
            .O(N__70740),
            .I(N__70737));
    LocalMux I__15700 (
            .O(N__70737),
            .I(N__70734));
    Span4Mux_v I__15699 (
            .O(N__70734),
            .I(N__70731));
    Odrv4 I__15698 (
            .O(N__70731),
            .I(\pid_side.error_i_reg_9_sn_13 ));
    CascadeMux I__15697 (
            .O(N__70728),
            .I(\pid_side.N_127_cascade_ ));
    CascadeMux I__15696 (
            .O(N__70725),
            .I(N__70722));
    InMux I__15695 (
            .O(N__70722),
            .I(N__70719));
    LocalMux I__15694 (
            .O(N__70719),
            .I(N__70716));
    Span4Mux_v I__15693 (
            .O(N__70716),
            .I(N__70713));
    Odrv4 I__15692 (
            .O(N__70713),
            .I(\pid_side.error_i_regZ0Z_13 ));
    InMux I__15691 (
            .O(N__70710),
            .I(N__70704));
    InMux I__15690 (
            .O(N__70709),
            .I(N__70704));
    LocalMux I__15689 (
            .O(N__70704),
            .I(N__70700));
    InMux I__15688 (
            .O(N__70703),
            .I(N__70697));
    Span4Mux_v I__15687 (
            .O(N__70700),
            .I(N__70694));
    LocalMux I__15686 (
            .O(N__70697),
            .I(N__70691));
    Span4Mux_h I__15685 (
            .O(N__70694),
            .I(N__70686));
    Span4Mux_h I__15684 (
            .O(N__70691),
            .I(N__70686));
    Span4Mux_h I__15683 (
            .O(N__70686),
            .I(N__70683));
    Odrv4 I__15682 (
            .O(N__70683),
            .I(xy_ki_6));
    CascadeMux I__15681 (
            .O(N__70680),
            .I(N__70677));
    InMux I__15680 (
            .O(N__70677),
            .I(N__70672));
    InMux I__15679 (
            .O(N__70676),
            .I(N__70669));
    InMux I__15678 (
            .O(N__70675),
            .I(N__70666));
    LocalMux I__15677 (
            .O(N__70672),
            .I(N__70663));
    LocalMux I__15676 (
            .O(N__70669),
            .I(N__70660));
    LocalMux I__15675 (
            .O(N__70666),
            .I(N__70657));
    Span4Mux_h I__15674 (
            .O(N__70663),
            .I(N__70652));
    Span4Mux_h I__15673 (
            .O(N__70660),
            .I(N__70652));
    Span4Mux_h I__15672 (
            .O(N__70657),
            .I(N__70649));
    Span4Mux_h I__15671 (
            .O(N__70652),
            .I(N__70646));
    Span4Mux_h I__15670 (
            .O(N__70649),
            .I(N__70643));
    Odrv4 I__15669 (
            .O(N__70646),
            .I(xy_ki_5));
    Odrv4 I__15668 (
            .O(N__70643),
            .I(xy_ki_5));
    CascadeMux I__15667 (
            .O(N__70638),
            .I(N__70635));
    InMux I__15666 (
            .O(N__70635),
            .I(N__70630));
    InMux I__15665 (
            .O(N__70634),
            .I(N__70625));
    InMux I__15664 (
            .O(N__70633),
            .I(N__70625));
    LocalMux I__15663 (
            .O(N__70630),
            .I(N__70622));
    LocalMux I__15662 (
            .O(N__70625),
            .I(N__70619));
    Span4Mux_h I__15661 (
            .O(N__70622),
            .I(N__70616));
    Span4Mux_h I__15660 (
            .O(N__70619),
            .I(N__70613));
    Span4Mux_h I__15659 (
            .O(N__70616),
            .I(N__70610));
    Span4Mux_h I__15658 (
            .O(N__70613),
            .I(N__70607));
    Odrv4 I__15657 (
            .O(N__70610),
            .I(xy_ki_7));
    Odrv4 I__15656 (
            .O(N__70607),
            .I(xy_ki_7));
    InMux I__15655 (
            .O(N__70602),
            .I(N__70596));
    InMux I__15654 (
            .O(N__70601),
            .I(N__70596));
    LocalMux I__15653 (
            .O(N__70596),
            .I(N__70593));
    Span4Mux_h I__15652 (
            .O(N__70593),
            .I(N__70590));
    Sp12to4 I__15651 (
            .O(N__70590),
            .I(N__70587));
    Odrv12 I__15650 (
            .O(N__70587),
            .I(pid_side_m153_e_4));
    InMux I__15649 (
            .O(N__70584),
            .I(N__70581));
    LocalMux I__15648 (
            .O(N__70581),
            .I(N__70576));
    InMux I__15647 (
            .O(N__70580),
            .I(N__70573));
    InMux I__15646 (
            .O(N__70579),
            .I(N__70569));
    Span4Mux_v I__15645 (
            .O(N__70576),
            .I(N__70566));
    LocalMux I__15644 (
            .O(N__70573),
            .I(N__70563));
    InMux I__15643 (
            .O(N__70572),
            .I(N__70560));
    LocalMux I__15642 (
            .O(N__70569),
            .I(N__70557));
    Odrv4 I__15641 (
            .O(N__70566),
            .I(\pid_side.m1_0_03 ));
    Odrv4 I__15640 (
            .O(N__70563),
            .I(\pid_side.m1_0_03 ));
    LocalMux I__15639 (
            .O(N__70560),
            .I(\pid_side.m1_0_03 ));
    Odrv4 I__15638 (
            .O(N__70557),
            .I(\pid_side.m1_0_03 ));
    CascadeMux I__15637 (
            .O(N__70548),
            .I(\pid_side.N_89_0_1_cascade_ ));
    InMux I__15636 (
            .O(N__70545),
            .I(N__70542));
    LocalMux I__15635 (
            .O(N__70542),
            .I(\pid_side.error_i_reg_9_rn_2_13 ));
    InMux I__15634 (
            .O(N__70539),
            .I(N__70536));
    LocalMux I__15633 (
            .O(N__70536),
            .I(N__70532));
    InMux I__15632 (
            .O(N__70535),
            .I(N__70529));
    Span4Mux_h I__15631 (
            .O(N__70532),
            .I(N__70524));
    LocalMux I__15630 (
            .O(N__70529),
            .I(N__70524));
    Span4Mux_h I__15629 (
            .O(N__70524),
            .I(N__70521));
    Span4Mux_h I__15628 (
            .O(N__70521),
            .I(N__70518));
    Odrv4 I__15627 (
            .O(N__70518),
            .I(\pid_front.error_p_reg_esr_RNITCC61Z0Z_18 ));
    InMux I__15626 (
            .O(N__70515),
            .I(N__70512));
    LocalMux I__15625 (
            .O(N__70512),
            .I(N__70509));
    Span4Mux_h I__15624 (
            .O(N__70509),
            .I(N__70505));
    InMux I__15623 (
            .O(N__70508),
            .I(N__70502));
    Span4Mux_h I__15622 (
            .O(N__70505),
            .I(N__70499));
    LocalMux I__15621 (
            .O(N__70502),
            .I(\pid_front.error_d_reg_prevZ0Z_18 ));
    Odrv4 I__15620 (
            .O(N__70499),
            .I(\pid_front.error_d_reg_prevZ0Z_18 ));
    CEMux I__15619 (
            .O(N__70494),
            .I(N__70491));
    LocalMux I__15618 (
            .O(N__70491),
            .I(N__70487));
    CEMux I__15617 (
            .O(N__70490),
            .I(N__70484));
    Span4Mux_h I__15616 (
            .O(N__70487),
            .I(N__70479));
    LocalMux I__15615 (
            .O(N__70484),
            .I(N__70476));
    CEMux I__15614 (
            .O(N__70483),
            .I(N__70473));
    CEMux I__15613 (
            .O(N__70482),
            .I(N__70464));
    Span4Mux_v I__15612 (
            .O(N__70479),
            .I(N__70457));
    Span4Mux_v I__15611 (
            .O(N__70476),
            .I(N__70457));
    LocalMux I__15610 (
            .O(N__70473),
            .I(N__70457));
    CEMux I__15609 (
            .O(N__70472),
            .I(N__70454));
    CEMux I__15608 (
            .O(N__70471),
            .I(N__70450));
    CEMux I__15607 (
            .O(N__70470),
            .I(N__70447));
    CEMux I__15606 (
            .O(N__70469),
            .I(N__70444));
    CEMux I__15605 (
            .O(N__70468),
            .I(N__70441));
    CEMux I__15604 (
            .O(N__70467),
            .I(N__70438));
    LocalMux I__15603 (
            .O(N__70464),
            .I(N__70435));
    Span4Mux_v I__15602 (
            .O(N__70457),
            .I(N__70432));
    LocalMux I__15601 (
            .O(N__70454),
            .I(N__70429));
    CEMux I__15600 (
            .O(N__70453),
            .I(N__70424));
    LocalMux I__15599 (
            .O(N__70450),
            .I(N__70421));
    LocalMux I__15598 (
            .O(N__70447),
            .I(N__70416));
    LocalMux I__15597 (
            .O(N__70444),
            .I(N__70416));
    LocalMux I__15596 (
            .O(N__70441),
            .I(N__70413));
    LocalMux I__15595 (
            .O(N__70438),
            .I(N__70410));
    Span4Mux_h I__15594 (
            .O(N__70435),
            .I(N__70407));
    Span4Mux_h I__15593 (
            .O(N__70432),
            .I(N__70402));
    Span4Mux_v I__15592 (
            .O(N__70429),
            .I(N__70402));
    CEMux I__15591 (
            .O(N__70428),
            .I(N__70399));
    CEMux I__15590 (
            .O(N__70427),
            .I(N__70396));
    LocalMux I__15589 (
            .O(N__70424),
            .I(N__70393));
    Span4Mux_h I__15588 (
            .O(N__70421),
            .I(N__70390));
    Span4Mux_v I__15587 (
            .O(N__70416),
            .I(N__70387));
    Span4Mux_v I__15586 (
            .O(N__70413),
            .I(N__70384));
    Span4Mux_v I__15585 (
            .O(N__70410),
            .I(N__70377));
    Span4Mux_h I__15584 (
            .O(N__70407),
            .I(N__70377));
    Span4Mux_h I__15583 (
            .O(N__70402),
            .I(N__70377));
    LocalMux I__15582 (
            .O(N__70399),
            .I(\pid_front.N_764_0 ));
    LocalMux I__15581 (
            .O(N__70396),
            .I(\pid_front.N_764_0 ));
    Odrv12 I__15580 (
            .O(N__70393),
            .I(\pid_front.N_764_0 ));
    Odrv4 I__15579 (
            .O(N__70390),
            .I(\pid_front.N_764_0 ));
    Odrv4 I__15578 (
            .O(N__70387),
            .I(\pid_front.N_764_0 ));
    Odrv4 I__15577 (
            .O(N__70384),
            .I(\pid_front.N_764_0 ));
    Odrv4 I__15576 (
            .O(N__70377),
            .I(\pid_front.N_764_0 ));
    InMux I__15575 (
            .O(N__70362),
            .I(N__70359));
    LocalMux I__15574 (
            .O(N__70359),
            .I(N__70343));
    SRMux I__15573 (
            .O(N__70358),
            .I(N__70314));
    SRMux I__15572 (
            .O(N__70357),
            .I(N__70314));
    SRMux I__15571 (
            .O(N__70356),
            .I(N__70314));
    SRMux I__15570 (
            .O(N__70355),
            .I(N__70314));
    SRMux I__15569 (
            .O(N__70354),
            .I(N__70314));
    SRMux I__15568 (
            .O(N__70353),
            .I(N__70314));
    SRMux I__15567 (
            .O(N__70352),
            .I(N__70314));
    SRMux I__15566 (
            .O(N__70351),
            .I(N__70314));
    SRMux I__15565 (
            .O(N__70350),
            .I(N__70314));
    SRMux I__15564 (
            .O(N__70349),
            .I(N__70314));
    SRMux I__15563 (
            .O(N__70348),
            .I(N__70314));
    SRMux I__15562 (
            .O(N__70347),
            .I(N__70314));
    SRMux I__15561 (
            .O(N__70346),
            .I(N__70314));
    Glb2LocalMux I__15560 (
            .O(N__70343),
            .I(N__70314));
    GlobalMux I__15559 (
            .O(N__70314),
            .I(N__70311));
    gio2CtrlBuf I__15558 (
            .O(N__70311),
            .I(\pid_front.N_1705_g ));
    InMux I__15557 (
            .O(N__70308),
            .I(N__70302));
    InMux I__15556 (
            .O(N__70307),
            .I(N__70302));
    LocalMux I__15555 (
            .O(N__70302),
            .I(N__70299));
    Odrv12 I__15554 (
            .O(N__70299),
            .I(drone_H_disp_side_11));
    InMux I__15553 (
            .O(N__70296),
            .I(N__70293));
    LocalMux I__15552 (
            .O(N__70293),
            .I(N__70290));
    Span4Mux_v I__15551 (
            .O(N__70290),
            .I(N__70286));
    InMux I__15550 (
            .O(N__70289),
            .I(N__70283));
    Odrv4 I__15549 (
            .O(N__70286),
            .I(\pid_side.N_9_1 ));
    LocalMux I__15548 (
            .O(N__70283),
            .I(\pid_side.N_9_1 ));
    CascadeMux I__15547 (
            .O(N__70278),
            .I(\pid_side.m87_0_ns_1_cascade_ ));
    CascadeMux I__15546 (
            .O(N__70275),
            .I(\pid_side.N_88_0_cascade_ ));
    InMux I__15545 (
            .O(N__70272),
            .I(N__70263));
    InMux I__15544 (
            .O(N__70271),
            .I(N__70263));
    InMux I__15543 (
            .O(N__70270),
            .I(N__70263));
    LocalMux I__15542 (
            .O(N__70263),
            .I(\pid_side.N_90_0 ));
    InMux I__15541 (
            .O(N__70260),
            .I(N__70257));
    LocalMux I__15540 (
            .O(N__70257),
            .I(\pid_side.m21_ns_1 ));
    CascadeMux I__15539 (
            .O(N__70254),
            .I(\pid_side.g0_i_m4_1_cascade_ ));
    InMux I__15538 (
            .O(N__70251),
            .I(N__70248));
    LocalMux I__15537 (
            .O(N__70248),
            .I(N__70245));
    Odrv4 I__15536 (
            .O(N__70245),
            .I(\pid_side.N_8_0 ));
    CascadeMux I__15535 (
            .O(N__70242),
            .I(\pid_side.N_36_0_cascade_ ));
    InMux I__15534 (
            .O(N__70239),
            .I(N__70236));
    LocalMux I__15533 (
            .O(N__70236),
            .I(\pid_side.error_i_reg_esr_RNO_2Z0Z_16 ));
    InMux I__15532 (
            .O(N__70233),
            .I(N__70230));
    LocalMux I__15531 (
            .O(N__70230),
            .I(\pid_side.N_36_0 ));
    CascadeMux I__15530 (
            .O(N__70227),
            .I(\pid_side.N_57_0_cascade_ ));
    CascadeMux I__15529 (
            .O(N__70224),
            .I(\pid_side.N_59_0_cascade_ ));
    InMux I__15528 (
            .O(N__70221),
            .I(N__70218));
    LocalMux I__15527 (
            .O(N__70218),
            .I(\pid_side.N_89_i ));
    CascadeMux I__15526 (
            .O(N__70215),
            .I(N__70212));
    InMux I__15525 (
            .O(N__70212),
            .I(N__70209));
    LocalMux I__15524 (
            .O(N__70209),
            .I(\pid_side.error_i_regZ0Z_24 ));
    InMux I__15523 (
            .O(N__70206),
            .I(N__70203));
    LocalMux I__15522 (
            .O(N__70203),
            .I(N__70199));
    InMux I__15521 (
            .O(N__70202),
            .I(N__70196));
    Span4Mux_h I__15520 (
            .O(N__70199),
            .I(N__70193));
    LocalMux I__15519 (
            .O(N__70196),
            .I(N__70190));
    Span4Mux_h I__15518 (
            .O(N__70193),
            .I(N__70185));
    Span4Mux_v I__15517 (
            .O(N__70190),
            .I(N__70185));
    Span4Mux_v I__15516 (
            .O(N__70185),
            .I(N__70182));
    Sp12to4 I__15515 (
            .O(N__70182),
            .I(N__70179));
    Odrv12 I__15514 (
            .O(N__70179),
            .I(\pid_front.error_p_regZ0Z_18 ));
    InMux I__15513 (
            .O(N__70176),
            .I(N__70173));
    LocalMux I__15512 (
            .O(N__70173),
            .I(N__70170));
    Odrv4 I__15511 (
            .O(N__70170),
            .I(\pid_side.error_d_reg_prev_esr_RNISM2K9Z0Z_15 ));
    CascadeMux I__15510 (
            .O(N__70167),
            .I(\pid_side.un1_pid_prereg_0_5_cascade_ ));
    CascadeMux I__15509 (
            .O(N__70164),
            .I(N__70161));
    InMux I__15508 (
            .O(N__70161),
            .I(N__70158));
    LocalMux I__15507 (
            .O(N__70158),
            .I(N__70155));
    Odrv4 I__15506 (
            .O(N__70155),
            .I(\pid_side.error_d_reg_prev_esr_RNIMK2Q4Z0Z_16 ));
    InMux I__15505 (
            .O(N__70152),
            .I(N__70149));
    LocalMux I__15504 (
            .O(N__70149),
            .I(N__70144));
    InMux I__15503 (
            .O(N__70148),
            .I(N__70139));
    InMux I__15502 (
            .O(N__70147),
            .I(N__70139));
    Odrv12 I__15501 (
            .O(N__70144),
            .I(\pid_side.error_i_reg_esr_RNI0JRRZ0Z_18 ));
    LocalMux I__15500 (
            .O(N__70139),
            .I(\pid_side.error_i_reg_esr_RNI0JRRZ0Z_18 ));
    InMux I__15499 (
            .O(N__70134),
            .I(N__70128));
    InMux I__15498 (
            .O(N__70133),
            .I(N__70128));
    LocalMux I__15497 (
            .O(N__70128),
            .I(\pid_side.un1_pid_prereg_0_5 ));
    CascadeMux I__15496 (
            .O(N__70125),
            .I(\pid_side.un1_pid_prereg_0_6_cascade_ ));
    InMux I__15495 (
            .O(N__70122),
            .I(N__70119));
    LocalMux I__15494 (
            .O(N__70119),
            .I(N__70116));
    Odrv4 I__15493 (
            .O(N__70116),
            .I(\pid_side.error_d_reg_prev_esr_RNISR7K9Z0Z_16 ));
    CascadeMux I__15492 (
            .O(N__70113),
            .I(\pid_side.un1_pid_prereg_0_7_cascade_ ));
    CascadeMux I__15491 (
            .O(N__70110),
            .I(N__70107));
    InMux I__15490 (
            .O(N__70107),
            .I(N__70104));
    LocalMux I__15489 (
            .O(N__70104),
            .I(N__70101));
    Odrv12 I__15488 (
            .O(N__70101),
            .I(\pid_side.error_d_reg_prev_esr_RNI675Q4Z0Z_17 ));
    InMux I__15487 (
            .O(N__70098),
            .I(N__70095));
    LocalMux I__15486 (
            .O(N__70095),
            .I(N__70092));
    Span4Mux_v I__15485 (
            .O(N__70092),
            .I(N__70087));
    InMux I__15484 (
            .O(N__70091),
            .I(N__70084));
    InMux I__15483 (
            .O(N__70090),
            .I(N__70081));
    Odrv4 I__15482 (
            .O(N__70087),
            .I(\pid_side.error_i_reg_esr_RNIUFQRZ0Z_17 ));
    LocalMux I__15481 (
            .O(N__70084),
            .I(\pid_side.error_i_reg_esr_RNIUFQRZ0Z_17 ));
    LocalMux I__15480 (
            .O(N__70081),
            .I(\pid_side.error_i_reg_esr_RNIUFQRZ0Z_17 ));
    InMux I__15479 (
            .O(N__70074),
            .I(N__70065));
    InMux I__15478 (
            .O(N__70073),
            .I(N__70065));
    InMux I__15477 (
            .O(N__70072),
            .I(N__70065));
    LocalMux I__15476 (
            .O(N__70065),
            .I(\pid_side.un1_pid_prereg_0_4 ));
    InMux I__15475 (
            .O(N__70062),
            .I(N__70059));
    LocalMux I__15474 (
            .O(N__70059),
            .I(N__70056));
    Odrv4 I__15473 (
            .O(N__70056),
            .I(\pid_side.error_d_reg_prev_esr_RNI72LM6Z0Z_22 ));
    CascadeMux I__15472 (
            .O(N__70053),
            .I(N__70050));
    InMux I__15471 (
            .O(N__70050),
            .I(N__70047));
    LocalMux I__15470 (
            .O(N__70047),
            .I(N__70044));
    Odrv4 I__15469 (
            .O(N__70044),
            .I(\pid_side.error_d_reg_prev_esr_RNI30AB3Z0Z_22 ));
    InMux I__15468 (
            .O(N__70041),
            .I(N__70038));
    LocalMux I__15467 (
            .O(N__70038),
            .I(N__70035));
    Span4Mux_v I__15466 (
            .O(N__70035),
            .I(N__70032));
    Span4Mux_h I__15465 (
            .O(N__70032),
            .I(N__70029));
    Odrv4 I__15464 (
            .O(N__70029),
            .I(\pid_side.pid_preregZ0Z_29 ));
    InMux I__15463 (
            .O(N__70026),
            .I(\pid_side.un1_pid_prereg_0_cry_28 ));
    InMux I__15462 (
            .O(N__70023),
            .I(N__70020));
    LocalMux I__15461 (
            .O(N__70020),
            .I(N__70017));
    Odrv4 I__15460 (
            .O(N__70017),
            .I(\pid_side.un1_pid_prereg_0_axb_30 ));
    InMux I__15459 (
            .O(N__70014),
            .I(\pid_side.un1_pid_prereg_0_cry_29 ));
    CascadeMux I__15458 (
            .O(N__70011),
            .I(N__70007));
    CascadeMux I__15457 (
            .O(N__70010),
            .I(N__70002));
    InMux I__15456 (
            .O(N__70007),
            .I(N__69985));
    InMux I__15455 (
            .O(N__70006),
            .I(N__69980));
    InMux I__15454 (
            .O(N__70005),
            .I(N__69980));
    InMux I__15453 (
            .O(N__70002),
            .I(N__69973));
    InMux I__15452 (
            .O(N__70001),
            .I(N__69973));
    InMux I__15451 (
            .O(N__70000),
            .I(N__69973));
    InMux I__15450 (
            .O(N__69999),
            .I(N__69956));
    InMux I__15449 (
            .O(N__69998),
            .I(N__69956));
    InMux I__15448 (
            .O(N__69997),
            .I(N__69956));
    InMux I__15447 (
            .O(N__69996),
            .I(N__69956));
    InMux I__15446 (
            .O(N__69995),
            .I(N__69956));
    InMux I__15445 (
            .O(N__69994),
            .I(N__69956));
    InMux I__15444 (
            .O(N__69993),
            .I(N__69956));
    InMux I__15443 (
            .O(N__69992),
            .I(N__69956));
    InMux I__15442 (
            .O(N__69991),
            .I(N__69951));
    InMux I__15441 (
            .O(N__69990),
            .I(N__69951));
    InMux I__15440 (
            .O(N__69989),
            .I(N__69946));
    InMux I__15439 (
            .O(N__69988),
            .I(N__69946));
    LocalMux I__15438 (
            .O(N__69985),
            .I(N__69943));
    LocalMux I__15437 (
            .O(N__69980),
            .I(N__69938));
    LocalMux I__15436 (
            .O(N__69973),
            .I(N__69938));
    LocalMux I__15435 (
            .O(N__69956),
            .I(N__69935));
    LocalMux I__15434 (
            .O(N__69951),
            .I(N__69930));
    LocalMux I__15433 (
            .O(N__69946),
            .I(N__69930));
    Span4Mux_v I__15432 (
            .O(N__69943),
            .I(N__69925));
    Span4Mux_h I__15431 (
            .O(N__69938),
            .I(N__69925));
    Span12Mux_h I__15430 (
            .O(N__69935),
            .I(N__69922));
    Span12Mux_v I__15429 (
            .O(N__69930),
            .I(N__69919));
    Span4Mux_v I__15428 (
            .O(N__69925),
            .I(N__69916));
    Odrv12 I__15427 (
            .O(N__69922),
            .I(\pid_side.pid_preregZ0Z_30 ));
    Odrv12 I__15426 (
            .O(N__69919),
            .I(\pid_side.pid_preregZ0Z_30 ));
    Odrv4 I__15425 (
            .O(N__69916),
            .I(\pid_side.pid_preregZ0Z_30 ));
    InMux I__15424 (
            .O(N__69909),
            .I(N__69905));
    InMux I__15423 (
            .O(N__69908),
            .I(N__69902));
    LocalMux I__15422 (
            .O(N__69905),
            .I(N__69888));
    LocalMux I__15421 (
            .O(N__69902),
            .I(N__69885));
    CEMux I__15420 (
            .O(N__69901),
            .I(N__69858));
    CEMux I__15419 (
            .O(N__69900),
            .I(N__69858));
    CEMux I__15418 (
            .O(N__69899),
            .I(N__69858));
    CEMux I__15417 (
            .O(N__69898),
            .I(N__69858));
    CEMux I__15416 (
            .O(N__69897),
            .I(N__69858));
    CEMux I__15415 (
            .O(N__69896),
            .I(N__69858));
    CEMux I__15414 (
            .O(N__69895),
            .I(N__69858));
    CEMux I__15413 (
            .O(N__69894),
            .I(N__69858));
    CEMux I__15412 (
            .O(N__69893),
            .I(N__69858));
    CEMux I__15411 (
            .O(N__69892),
            .I(N__69858));
    CEMux I__15410 (
            .O(N__69891),
            .I(N__69858));
    Glb2LocalMux I__15409 (
            .O(N__69888),
            .I(N__69858));
    Glb2LocalMux I__15408 (
            .O(N__69885),
            .I(N__69858));
    GlobalMux I__15407 (
            .O(N__69858),
            .I(N__69855));
    gio2CtrlBuf I__15406 (
            .O(N__69855),
            .I(\pid_side.N_838_g ));
    InMux I__15405 (
            .O(N__69852),
            .I(N__69849));
    LocalMux I__15404 (
            .O(N__69849),
            .I(N__69846));
    Span4Mux_v I__15403 (
            .O(N__69846),
            .I(N__69843));
    Odrv4 I__15402 (
            .O(N__69843),
            .I(\pid_side.un1_pid_prereg_370_1 ));
    InMux I__15401 (
            .O(N__69840),
            .I(N__69837));
    LocalMux I__15400 (
            .O(N__69837),
            .I(N__69833));
    InMux I__15399 (
            .O(N__69836),
            .I(N__69830));
    Span4Mux_v I__15398 (
            .O(N__69833),
            .I(N__69827));
    LocalMux I__15397 (
            .O(N__69830),
            .I(N__69823));
    Span4Mux_v I__15396 (
            .O(N__69827),
            .I(N__69820));
    InMux I__15395 (
            .O(N__69826),
            .I(N__69817));
    Span4Mux_h I__15394 (
            .O(N__69823),
            .I(N__69814));
    Odrv4 I__15393 (
            .O(N__69820),
            .I(\pid_side.error_i_reg_esr_RNIM5PSZ0Z_22 ));
    LocalMux I__15392 (
            .O(N__69817),
            .I(\pid_side.error_i_reg_esr_RNIM5PSZ0Z_22 ));
    Odrv4 I__15391 (
            .O(N__69814),
            .I(\pid_side.error_i_reg_esr_RNIM5PSZ0Z_22 ));
    CascadeMux I__15390 (
            .O(N__69807),
            .I(\pid_side.un1_pid_prereg_0_1_cascade_ ));
    CascadeMux I__15389 (
            .O(N__69804),
            .I(N__69801));
    InMux I__15388 (
            .O(N__69801),
            .I(N__69798));
    LocalMux I__15387 (
            .O(N__69798),
            .I(N__69795));
    Odrv4 I__15386 (
            .O(N__69795),
            .I(\pid_side.error_d_reg_prev_esr_RNIMFTP4Z0Z_14 ));
    InMux I__15385 (
            .O(N__69792),
            .I(N__69789));
    LocalMux I__15384 (
            .O(N__69789),
            .I(N__69784));
    InMux I__15383 (
            .O(N__69788),
            .I(N__69779));
    InMux I__15382 (
            .O(N__69787),
            .I(N__69779));
    Odrv12 I__15381 (
            .O(N__69784),
            .I(\pid_side.error_i_reg_esr_RNISCPRZ0Z_16 ));
    LocalMux I__15380 (
            .O(N__69779),
            .I(\pid_side.error_i_reg_esr_RNISCPRZ0Z_16 ));
    CascadeMux I__15379 (
            .O(N__69774),
            .I(\pid_side.un1_pid_prereg_0_2_cascade_ ));
    InMux I__15378 (
            .O(N__69771),
            .I(N__69768));
    LocalMux I__15377 (
            .O(N__69768),
            .I(N__69765));
    Odrv4 I__15376 (
            .O(N__69765),
            .I(\pid_side.error_d_reg_prev_esr_RNISHTJ9Z0Z_14 ));
    InMux I__15375 (
            .O(N__69762),
            .I(N__69759));
    LocalMux I__15374 (
            .O(N__69759),
            .I(N__69756));
    Span4Mux_h I__15373 (
            .O(N__69756),
            .I(N__69753));
    Odrv4 I__15372 (
            .O(N__69753),
            .I(\pid_side.pid_preregZ0Z_21 ));
    InMux I__15371 (
            .O(N__69750),
            .I(\pid_side.un1_pid_prereg_0_cry_20 ));
    InMux I__15370 (
            .O(N__69747),
            .I(N__69744));
    LocalMux I__15369 (
            .O(N__69744),
            .I(N__69741));
    Span4Mux_h I__15368 (
            .O(N__69741),
            .I(N__69738));
    Odrv4 I__15367 (
            .O(N__69738),
            .I(\pid_side.pid_preregZ0Z_22 ));
    InMux I__15366 (
            .O(N__69735),
            .I(\pid_side.un1_pid_prereg_0_cry_21 ));
    CascadeMux I__15365 (
            .O(N__69732),
            .I(N__69729));
    InMux I__15364 (
            .O(N__69729),
            .I(N__69726));
    LocalMux I__15363 (
            .O(N__69726),
            .I(N__69723));
    Span4Mux_v I__15362 (
            .O(N__69723),
            .I(N__69720));
    Odrv4 I__15361 (
            .O(N__69720),
            .I(\pid_side.error_d_reg_prev_esr_RNIK1TV8Z0Z_22 ));
    CascadeMux I__15360 (
            .O(N__69717),
            .I(N__69714));
    InMux I__15359 (
            .O(N__69714),
            .I(N__69711));
    LocalMux I__15358 (
            .O(N__69711),
            .I(N__69708));
    Span4Mux_h I__15357 (
            .O(N__69708),
            .I(N__69705));
    Odrv4 I__15356 (
            .O(N__69705),
            .I(\pid_side.pid_preregZ0Z_23 ));
    InMux I__15355 (
            .O(N__69702),
            .I(bfn_17_14_0_));
    InMux I__15354 (
            .O(N__69699),
            .I(N__69696));
    LocalMux I__15353 (
            .O(N__69696),
            .I(N__69693));
    Odrv4 I__15352 (
            .O(N__69693),
            .I(\pid_side.error_d_reg_prev_esr_RNIFQK34Z0Z_22 ));
    CascadeMux I__15351 (
            .O(N__69690),
            .I(N__69687));
    InMux I__15350 (
            .O(N__69687),
            .I(N__69684));
    LocalMux I__15349 (
            .O(N__69684),
            .I(N__69681));
    Odrv12 I__15348 (
            .O(N__69681),
            .I(\pid_side.error_d_reg_prev_esr_RNI33ME7Z0Z_22 ));
    InMux I__15347 (
            .O(N__69678),
            .I(N__69675));
    LocalMux I__15346 (
            .O(N__69675),
            .I(N__69672));
    Span4Mux_v I__15345 (
            .O(N__69672),
            .I(N__69669));
    Span4Mux_v I__15344 (
            .O(N__69669),
            .I(N__69666));
    Odrv4 I__15343 (
            .O(N__69666),
            .I(\pid_side.pid_preregZ0Z_24 ));
    InMux I__15342 (
            .O(N__69663),
            .I(\pid_side.un1_pid_prereg_0_cry_23 ));
    InMux I__15341 (
            .O(N__69660),
            .I(N__69657));
    LocalMux I__15340 (
            .O(N__69657),
            .I(N__69654));
    Odrv12 I__15339 (
            .O(N__69654),
            .I(\pid_side.error_d_reg_prev_esr_RNICN4M6Z0Z_22 ));
    CascadeMux I__15338 (
            .O(N__69651),
            .I(N__69648));
    InMux I__15337 (
            .O(N__69648),
            .I(N__69645));
    LocalMux I__15336 (
            .O(N__69645),
            .I(N__69642));
    Odrv12 I__15335 (
            .O(N__69642),
            .I(\pid_side.error_d_reg_prev_esr_RNIK81B3Z0Z_22 ));
    InMux I__15334 (
            .O(N__69639),
            .I(N__69636));
    LocalMux I__15333 (
            .O(N__69636),
            .I(N__69633));
    Span4Mux_h I__15332 (
            .O(N__69633),
            .I(N__69630));
    Span4Mux_v I__15331 (
            .O(N__69630),
            .I(N__69627));
    Odrv4 I__15330 (
            .O(N__69627),
            .I(\pid_side.pid_preregZ0Z_25 ));
    InMux I__15329 (
            .O(N__69624),
            .I(\pid_side.un1_pid_prereg_0_cry_24 ));
    CascadeMux I__15328 (
            .O(N__69621),
            .I(N__69618));
    InMux I__15327 (
            .O(N__69618),
            .I(N__69615));
    LocalMux I__15326 (
            .O(N__69615),
            .I(N__69612));
    Span4Mux_v I__15325 (
            .O(N__69612),
            .I(N__69609));
    Odrv4 I__15324 (
            .O(N__69609),
            .I(\pid_side.error_d_reg_prev_esr_RNIOE3B3Z0Z_22 ));
    InMux I__15323 (
            .O(N__69606),
            .I(N__69603));
    LocalMux I__15322 (
            .O(N__69603),
            .I(N__69600));
    Span4Mux_h I__15321 (
            .O(N__69600),
            .I(N__69597));
    Span4Mux_v I__15320 (
            .O(N__69597),
            .I(N__69594));
    Odrv4 I__15319 (
            .O(N__69594),
            .I(\pid_side.pid_preregZ0Z_26 ));
    InMux I__15318 (
            .O(N__69591),
            .I(\pid_side.un1_pid_prereg_0_cry_25 ));
    CascadeMux I__15317 (
            .O(N__69588),
            .I(N__69585));
    InMux I__15316 (
            .O(N__69585),
            .I(N__69582));
    LocalMux I__15315 (
            .O(N__69582),
            .I(N__69579));
    Odrv12 I__15314 (
            .O(N__69579),
            .I(\pid_side.error_d_reg_prev_esr_RNISFDM6Z0Z_22 ));
    CascadeMux I__15313 (
            .O(N__69576),
            .I(N__69573));
    InMux I__15312 (
            .O(N__69573),
            .I(N__69570));
    LocalMux I__15311 (
            .O(N__69570),
            .I(N__69567));
    Span4Mux_v I__15310 (
            .O(N__69567),
            .I(N__69564));
    Span4Mux_v I__15309 (
            .O(N__69564),
            .I(N__69561));
    Odrv4 I__15308 (
            .O(N__69561),
            .I(\pid_side.pid_preregZ0Z_27 ));
    InMux I__15307 (
            .O(N__69558),
            .I(\pid_side.un1_pid_prereg_0_cry_26 ));
    InMux I__15306 (
            .O(N__69555),
            .I(N__69552));
    LocalMux I__15305 (
            .O(N__69552),
            .I(N__69549));
    Odrv4 I__15304 (
            .O(N__69549),
            .I(\pid_side.error_d_reg_prev_esr_RNI3RHM6Z0Z_22 ));
    CascadeMux I__15303 (
            .O(N__69546),
            .I(N__69543));
    InMux I__15302 (
            .O(N__69543),
            .I(N__69540));
    LocalMux I__15301 (
            .O(N__69540),
            .I(N__69537));
    Odrv4 I__15300 (
            .O(N__69537),
            .I(\pid_side.error_d_reg_prev_esr_RNI0R7B3Z0Z_22 ));
    InMux I__15299 (
            .O(N__69534),
            .I(N__69531));
    LocalMux I__15298 (
            .O(N__69531),
            .I(N__69528));
    Span4Mux_h I__15297 (
            .O(N__69528),
            .I(N__69525));
    Odrv4 I__15296 (
            .O(N__69525),
            .I(\pid_side.pid_preregZ0Z_28 ));
    InMux I__15295 (
            .O(N__69522),
            .I(\pid_side.un1_pid_prereg_0_cry_27 ));
    CascadeMux I__15294 (
            .O(N__69519),
            .I(N__69516));
    InMux I__15293 (
            .O(N__69516),
            .I(N__69513));
    LocalMux I__15292 (
            .O(N__69513),
            .I(N__69510));
    Span4Mux_h I__15291 (
            .O(N__69510),
            .I(N__69507));
    Span4Mux_h I__15290 (
            .O(N__69507),
            .I(N__69504));
    Odrv4 I__15289 (
            .O(N__69504),
            .I(\pid_side.error_d_reg_prev_esr_RNITU3P4Z0Z_10 ));
    InMux I__15288 (
            .O(N__69501),
            .I(N__69494));
    InMux I__15287 (
            .O(N__69500),
            .I(N__69489));
    InMux I__15286 (
            .O(N__69499),
            .I(N__69489));
    InMux I__15285 (
            .O(N__69498),
            .I(N__69484));
    InMux I__15284 (
            .O(N__69497),
            .I(N__69484));
    LocalMux I__15283 (
            .O(N__69494),
            .I(N__69479));
    LocalMux I__15282 (
            .O(N__69489),
            .I(N__69479));
    LocalMux I__15281 (
            .O(N__69484),
            .I(N__69476));
    Span4Mux_v I__15280 (
            .O(N__69479),
            .I(N__69473));
    Span4Mux_h I__15279 (
            .O(N__69476),
            .I(N__69470));
    Odrv4 I__15278 (
            .O(N__69473),
            .I(\pid_side.pid_preregZ0Z_12 ));
    Odrv4 I__15277 (
            .O(N__69470),
            .I(\pid_side.pid_preregZ0Z_12 ));
    InMux I__15276 (
            .O(N__69465),
            .I(\pid_side.un1_pid_prereg_0_cry_11 ));
    InMux I__15275 (
            .O(N__69462),
            .I(\pid_side.un1_pid_prereg_0_cry_12 ));
    InMux I__15274 (
            .O(N__69459),
            .I(N__69456));
    LocalMux I__15273 (
            .O(N__69456),
            .I(N__69453));
    Odrv12 I__15272 (
            .O(N__69453),
            .I(\pid_side.un1_pid_prereg_0_cry_13_THRU_CO ));
    InMux I__15271 (
            .O(N__69450),
            .I(\pid_side.un1_pid_prereg_0_cry_13 ));
    InMux I__15270 (
            .O(N__69447),
            .I(bfn_17_13_0_));
    InMux I__15269 (
            .O(N__69444),
            .I(\pid_side.un1_pid_prereg_0_cry_15 ));
    InMux I__15268 (
            .O(N__69441),
            .I(\pid_side.un1_pid_prereg_0_cry_16 ));
    InMux I__15267 (
            .O(N__69438),
            .I(\pid_side.un1_pid_prereg_0_cry_17 ));
    InMux I__15266 (
            .O(N__69435),
            .I(\pid_side.un1_pid_prereg_0_cry_18 ));
    InMux I__15265 (
            .O(N__69432),
            .I(N__69429));
    LocalMux I__15264 (
            .O(N__69429),
            .I(N__69426));
    Span4Mux_v I__15263 (
            .O(N__69426),
            .I(N__69423));
    Odrv4 I__15262 (
            .O(N__69423),
            .I(\pid_side.pid_preregZ0Z_20 ));
    InMux I__15261 (
            .O(N__69420),
            .I(\pid_side.un1_pid_prereg_0_cry_19 ));
    CascadeMux I__15260 (
            .O(N__69417),
            .I(N__69413));
    InMux I__15259 (
            .O(N__69416),
            .I(N__69408));
    InMux I__15258 (
            .O(N__69413),
            .I(N__69405));
    InMux I__15257 (
            .O(N__69412),
            .I(N__69402));
    InMux I__15256 (
            .O(N__69411),
            .I(N__69399));
    LocalMux I__15255 (
            .O(N__69408),
            .I(N__69396));
    LocalMux I__15254 (
            .O(N__69405),
            .I(N__69389));
    LocalMux I__15253 (
            .O(N__69402),
            .I(N__69389));
    LocalMux I__15252 (
            .O(N__69399),
            .I(N__69389));
    Span4Mux_h I__15251 (
            .O(N__69396),
            .I(N__69386));
    Span4Mux_v I__15250 (
            .O(N__69389),
            .I(N__69383));
    Odrv4 I__15249 (
            .O(N__69386),
            .I(\pid_side.pid_preregZ0Z_4 ));
    Odrv4 I__15248 (
            .O(N__69383),
            .I(\pid_side.pid_preregZ0Z_4 ));
    InMux I__15247 (
            .O(N__69378),
            .I(\pid_side.un1_pid_prereg_0_cry_3 ));
    InMux I__15246 (
            .O(N__69375),
            .I(N__69370));
    InMux I__15245 (
            .O(N__69374),
            .I(N__69367));
    InMux I__15244 (
            .O(N__69373),
            .I(N__69363));
    LocalMux I__15243 (
            .O(N__69370),
            .I(N__69358));
    LocalMux I__15242 (
            .O(N__69367),
            .I(N__69358));
    InMux I__15241 (
            .O(N__69366),
            .I(N__69355));
    LocalMux I__15240 (
            .O(N__69363),
            .I(N__69348));
    Span4Mux_v I__15239 (
            .O(N__69358),
            .I(N__69348));
    LocalMux I__15238 (
            .O(N__69355),
            .I(N__69348));
    Span4Mux_h I__15237 (
            .O(N__69348),
            .I(N__69345));
    Odrv4 I__15236 (
            .O(N__69345),
            .I(\pid_side.pid_preregZ0Z_5 ));
    InMux I__15235 (
            .O(N__69342),
            .I(\pid_side.un1_pid_prereg_0_cry_4 ));
    InMux I__15234 (
            .O(N__69339),
            .I(\pid_side.un1_pid_prereg_0_cry_5 ));
    InMux I__15233 (
            .O(N__69336),
            .I(N__69333));
    LocalMux I__15232 (
            .O(N__69333),
            .I(N__69330));
    Odrv4 I__15231 (
            .O(N__69330),
            .I(\pid_side.error_p_reg_esr_RNIODMH3_0Z0Z_6 ));
    InMux I__15230 (
            .O(N__69327),
            .I(bfn_17_12_0_));
    InMux I__15229 (
            .O(N__69324),
            .I(N__69321));
    LocalMux I__15228 (
            .O(N__69321),
            .I(N__69318));
    Odrv12 I__15227 (
            .O(N__69318),
            .I(\pid_side.error_p_reg_esr_RNIKF8V6Z0Z_7 ));
    CascadeMux I__15226 (
            .O(N__69315),
            .I(N__69312));
    InMux I__15225 (
            .O(N__69312),
            .I(N__69308));
    InMux I__15224 (
            .O(N__69311),
            .I(N__69305));
    LocalMux I__15223 (
            .O(N__69308),
            .I(N__69302));
    LocalMux I__15222 (
            .O(N__69305),
            .I(\pid_side.error_p_reg_esr_RNIODMH3Z0Z_6 ));
    Odrv4 I__15221 (
            .O(N__69302),
            .I(\pid_side.error_p_reg_esr_RNIODMH3Z0Z_6 ));
    InMux I__15220 (
            .O(N__69297),
            .I(\pid_side.un1_pid_prereg_0_cry_7 ));
    InMux I__15219 (
            .O(N__69294),
            .I(N__69291));
    LocalMux I__15218 (
            .O(N__69291),
            .I(N__69288));
    Odrv12 I__15217 (
            .O(N__69288),
            .I(\pid_side.error_p_reg_esr_RNIECBV6Z0Z_8 ));
    InMux I__15216 (
            .O(N__69285),
            .I(N__69281));
    CascadeMux I__15215 (
            .O(N__69284),
            .I(N__69278));
    LocalMux I__15214 (
            .O(N__69281),
            .I(N__69275));
    InMux I__15213 (
            .O(N__69278),
            .I(N__69272));
    Span4Mux_v I__15212 (
            .O(N__69275),
            .I(N__69269));
    LocalMux I__15211 (
            .O(N__69272),
            .I(N__69266));
    Odrv4 I__15210 (
            .O(N__69269),
            .I(\pid_side.error_p_reg_esr_RNIS1ID3Z0Z_7 ));
    Odrv4 I__15209 (
            .O(N__69266),
            .I(\pid_side.error_p_reg_esr_RNIS1ID3Z0Z_7 ));
    InMux I__15208 (
            .O(N__69261),
            .I(\pid_side.un1_pid_prereg_0_cry_8 ));
    InMux I__15207 (
            .O(N__69258),
            .I(\pid_side.un1_pid_prereg_0_cry_9 ));
    InMux I__15206 (
            .O(N__69255),
            .I(\pid_side.un1_pid_prereg_0_cry_10 ));
    InMux I__15205 (
            .O(N__69252),
            .I(N__69248));
    InMux I__15204 (
            .O(N__69251),
            .I(N__69245));
    LocalMux I__15203 (
            .O(N__69248),
            .I(\pid_side.un1_pid_prereg_0_17 ));
    LocalMux I__15202 (
            .O(N__69245),
            .I(\pid_side.un1_pid_prereg_0_17 ));
    CascadeMux I__15201 (
            .O(N__69240),
            .I(\pid_side.un1_pid_prereg_0_18_cascade_ ));
    InMux I__15200 (
            .O(N__69237),
            .I(N__69232));
    InMux I__15199 (
            .O(N__69236),
            .I(N__69229));
    InMux I__15198 (
            .O(N__69235),
            .I(N__69226));
    LocalMux I__15197 (
            .O(N__69232),
            .I(N__69223));
    LocalMux I__15196 (
            .O(N__69229),
            .I(N__69218));
    LocalMux I__15195 (
            .O(N__69226),
            .I(N__69218));
    Span4Mux_v I__15194 (
            .O(N__69223),
            .I(N__69213));
    Span4Mux_v I__15193 (
            .O(N__69218),
            .I(N__69213));
    Odrv4 I__15192 (
            .O(N__69213),
            .I(\pid_side.error_i_reg_esr_RNIO8QSZ0Z_23 ));
    InMux I__15191 (
            .O(N__69210),
            .I(N__69201));
    InMux I__15190 (
            .O(N__69209),
            .I(N__69201));
    InMux I__15189 (
            .O(N__69208),
            .I(N__69201));
    LocalMux I__15188 (
            .O(N__69201),
            .I(\pid_side.un1_pid_prereg_0_16 ));
    CascadeMux I__15187 (
            .O(N__69198),
            .I(\pid_side.un1_pid_prereg_0_19_cascade_ ));
    InMux I__15186 (
            .O(N__69195),
            .I(N__69191));
    InMux I__15185 (
            .O(N__69194),
            .I(N__69188));
    LocalMux I__15184 (
            .O(N__69191),
            .I(N__69185));
    LocalMux I__15183 (
            .O(N__69188),
            .I(N__69181));
    Span4Mux_v I__15182 (
            .O(N__69185),
            .I(N__69178));
    InMux I__15181 (
            .O(N__69184),
            .I(N__69175));
    Span4Mux_v I__15180 (
            .O(N__69181),
            .I(N__69172));
    Span4Mux_h I__15179 (
            .O(N__69178),
            .I(N__69167));
    LocalMux I__15178 (
            .O(N__69175),
            .I(N__69167));
    Span4Mux_h I__15177 (
            .O(N__69172),
            .I(N__69164));
    Span4Mux_h I__15176 (
            .O(N__69167),
            .I(N__69161));
    Odrv4 I__15175 (
            .O(N__69164),
            .I(\pid_side.pid_preregZ0Z_0 ));
    Odrv4 I__15174 (
            .O(N__69161),
            .I(\pid_side.pid_preregZ0Z_0 ));
    InMux I__15173 (
            .O(N__69156),
            .I(\pid_side.un1_pid_prereg_0_cry_0_c_THRU_CO ));
    CascadeMux I__15172 (
            .O(N__69153),
            .I(N__69150));
    InMux I__15171 (
            .O(N__69150),
            .I(N__69147));
    LocalMux I__15170 (
            .O(N__69147),
            .I(N__69142));
    InMux I__15169 (
            .O(N__69146),
            .I(N__69139));
    InMux I__15168 (
            .O(N__69145),
            .I(N__69136));
    Span4Mux_v I__15167 (
            .O(N__69142),
            .I(N__69131));
    LocalMux I__15166 (
            .O(N__69139),
            .I(N__69131));
    LocalMux I__15165 (
            .O(N__69136),
            .I(N__69128));
    Span4Mux_h I__15164 (
            .O(N__69131),
            .I(N__69125));
    Odrv4 I__15163 (
            .O(N__69128),
            .I(\pid_side.pid_preregZ0Z_1 ));
    Odrv4 I__15162 (
            .O(N__69125),
            .I(\pid_side.pid_preregZ0Z_1 ));
    InMux I__15161 (
            .O(N__69120),
            .I(\pid_side.un1_pid_prereg_0_cry_0 ));
    InMux I__15160 (
            .O(N__69117),
            .I(N__69110));
    InMux I__15159 (
            .O(N__69116),
            .I(N__69110));
    InMux I__15158 (
            .O(N__69115),
            .I(N__69107));
    LocalMux I__15157 (
            .O(N__69110),
            .I(N__69104));
    LocalMux I__15156 (
            .O(N__69107),
            .I(N__69101));
    Span4Mux_h I__15155 (
            .O(N__69104),
            .I(N__69098));
    Odrv4 I__15154 (
            .O(N__69101),
            .I(\pid_side.pid_preregZ0Z_2 ));
    Odrv4 I__15153 (
            .O(N__69098),
            .I(\pid_side.pid_preregZ0Z_2 ));
    InMux I__15152 (
            .O(N__69093),
            .I(\pid_side.un1_pid_prereg_0_cry_1 ));
    CascadeMux I__15151 (
            .O(N__69090),
            .I(N__69086));
    CascadeMux I__15150 (
            .O(N__69089),
            .I(N__69082));
    InMux I__15149 (
            .O(N__69086),
            .I(N__69079));
    CascadeMux I__15148 (
            .O(N__69085),
            .I(N__69076));
    InMux I__15147 (
            .O(N__69082),
            .I(N__69073));
    LocalMux I__15146 (
            .O(N__69079),
            .I(N__69070));
    InMux I__15145 (
            .O(N__69076),
            .I(N__69067));
    LocalMux I__15144 (
            .O(N__69073),
            .I(N__69064));
    Span4Mux_v I__15143 (
            .O(N__69070),
            .I(N__69061));
    LocalMux I__15142 (
            .O(N__69067),
            .I(N__69058));
    Span4Mux_v I__15141 (
            .O(N__69064),
            .I(N__69055));
    Odrv4 I__15140 (
            .O(N__69061),
            .I(\pid_side.pid_preregZ0Z_3 ));
    Odrv12 I__15139 (
            .O(N__69058),
            .I(\pid_side.pid_preregZ0Z_3 ));
    Odrv4 I__15138 (
            .O(N__69055),
            .I(\pid_side.pid_preregZ0Z_3 ));
    InMux I__15137 (
            .O(N__69048),
            .I(\pid_side.un1_pid_prereg_0_cry_2 ));
    InMux I__15136 (
            .O(N__69045),
            .I(N__69039));
    InMux I__15135 (
            .O(N__69044),
            .I(N__69039));
    LocalMux I__15134 (
            .O(N__69039),
            .I(\pid_side.error_i_acumm_preregZ0Z_22 ));
    InMux I__15133 (
            .O(N__69036),
            .I(N__69030));
    InMux I__15132 (
            .O(N__69035),
            .I(N__69030));
    LocalMux I__15131 (
            .O(N__69030),
            .I(\pid_side.error_i_acumm_preregZ0Z_23 ));
    CascadeMux I__15130 (
            .O(N__69027),
            .I(N__69024));
    InMux I__15129 (
            .O(N__69024),
            .I(N__69018));
    InMux I__15128 (
            .O(N__69023),
            .I(N__69018));
    LocalMux I__15127 (
            .O(N__69018),
            .I(\pid_side.error_i_acumm_preregZ0Z_24 ));
    CascadeMux I__15126 (
            .O(N__69015),
            .I(N__69011));
    CascadeMux I__15125 (
            .O(N__69014),
            .I(N__69008));
    InMux I__15124 (
            .O(N__69011),
            .I(N__69005));
    InMux I__15123 (
            .O(N__69008),
            .I(N__69002));
    LocalMux I__15122 (
            .O(N__69005),
            .I(N__68999));
    LocalMux I__15121 (
            .O(N__69002),
            .I(\pid_side.error_i_acumm_preregZ0Z_17 ));
    Odrv4 I__15120 (
            .O(N__68999),
            .I(\pid_side.error_i_acumm_preregZ0Z_17 ));
    CascadeMux I__15119 (
            .O(N__68994),
            .I(N__68991));
    InMux I__15118 (
            .O(N__68991),
            .I(N__68986));
    InMux I__15117 (
            .O(N__68990),
            .I(N__68983));
    InMux I__15116 (
            .O(N__68989),
            .I(N__68980));
    LocalMux I__15115 (
            .O(N__68986),
            .I(N__68973));
    LocalMux I__15114 (
            .O(N__68983),
            .I(N__68973));
    LocalMux I__15113 (
            .O(N__68980),
            .I(N__68973));
    Span4Mux_h I__15112 (
            .O(N__68973),
            .I(N__68970));
    Odrv4 I__15111 (
            .O(N__68970),
            .I(\pid_side.error_i_acumm_preregZ0Z_5 ));
    CascadeMux I__15110 (
            .O(N__68967),
            .I(\pid_side.un1_pid_prereg_0_17_cascade_ ));
    InMux I__15109 (
            .O(N__68964),
            .I(N__68961));
    LocalMux I__15108 (
            .O(N__68961),
            .I(N__68957));
    InMux I__15107 (
            .O(N__68960),
            .I(N__68954));
    Odrv4 I__15106 (
            .O(N__68957),
            .I(\pid_side.un1_pid_prereg_0_14 ));
    LocalMux I__15105 (
            .O(N__68954),
            .I(\pid_side.un1_pid_prereg_0_14 ));
    CascadeMux I__15104 (
            .O(N__68949),
            .I(N__68946));
    InMux I__15103 (
            .O(N__68946),
            .I(N__68943));
    LocalMux I__15102 (
            .O(N__68943),
            .I(N__68940));
    Span4Mux_v I__15101 (
            .O(N__68940),
            .I(N__68936));
    InMux I__15100 (
            .O(N__68939),
            .I(N__68933));
    Odrv4 I__15099 (
            .O(N__68936),
            .I(\pid_side.un1_pid_prereg_0_15 ));
    LocalMux I__15098 (
            .O(N__68933),
            .I(\pid_side.un1_pid_prereg_0_15 ));
    InMux I__15097 (
            .O(N__68928),
            .I(N__68925));
    LocalMux I__15096 (
            .O(N__68925),
            .I(N__68920));
    InMux I__15095 (
            .O(N__68924),
            .I(N__68915));
    InMux I__15094 (
            .O(N__68923),
            .I(N__68915));
    Span4Mux_h I__15093 (
            .O(N__68920),
            .I(N__68910));
    LocalMux I__15092 (
            .O(N__68915),
            .I(N__68910));
    Span4Mux_v I__15091 (
            .O(N__68910),
            .I(N__68907));
    Odrv4 I__15090 (
            .O(N__68907),
            .I(\pid_side.error_i_reg_esr_RNIQBRSZ0Z_24 ));
    InMux I__15089 (
            .O(N__68904),
            .I(N__68896));
    InMux I__15088 (
            .O(N__68903),
            .I(N__68896));
    InMux I__15087 (
            .O(N__68902),
            .I(N__68891));
    InMux I__15086 (
            .O(N__68901),
            .I(N__68891));
    LocalMux I__15085 (
            .O(N__68896),
            .I(N__68888));
    LocalMux I__15084 (
            .O(N__68891),
            .I(N__68884));
    Span4Mux_v I__15083 (
            .O(N__68888),
            .I(N__68881));
    InMux I__15082 (
            .O(N__68887),
            .I(N__68878));
    Span4Mux_v I__15081 (
            .O(N__68884),
            .I(N__68875));
    Span4Mux_h I__15080 (
            .O(N__68881),
            .I(N__68870));
    LocalMux I__15079 (
            .O(N__68878),
            .I(N__68870));
    Span4Mux_h I__15078 (
            .O(N__68875),
            .I(N__68867));
    Span4Mux_h I__15077 (
            .O(N__68870),
            .I(N__68864));
    Odrv4 I__15076 (
            .O(N__68867),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_RNIUCMNZ0Z_1 ));
    Odrv4 I__15075 (
            .O(N__68864),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_RNIUCMNZ0Z_1 ));
    InMux I__15074 (
            .O(N__68859),
            .I(N__68856));
    LocalMux I__15073 (
            .O(N__68856),
            .I(\ppm_encoder_1.pulses2count_9_i_3_2 ));
    CascadeMux I__15072 (
            .O(N__68853),
            .I(N__68850));
    InMux I__15071 (
            .O(N__68850),
            .I(N__68847));
    LocalMux I__15070 (
            .O(N__68847),
            .I(N__68844));
    Span4Mux_v I__15069 (
            .O(N__68844),
            .I(N__68840));
    InMux I__15068 (
            .O(N__68843),
            .I(N__68837));
    Span4Mux_h I__15067 (
            .O(N__68840),
            .I(N__68831));
    LocalMux I__15066 (
            .O(N__68837),
            .I(N__68831));
    InMux I__15065 (
            .O(N__68836),
            .I(N__68828));
    Span4Mux_h I__15064 (
            .O(N__68831),
            .I(N__68825));
    LocalMux I__15063 (
            .O(N__68828),
            .I(\ppm_encoder_1.aileronZ0Z_2 ));
    Odrv4 I__15062 (
            .O(N__68825),
            .I(\ppm_encoder_1.aileronZ0Z_2 ));
    CascadeMux I__15061 (
            .O(N__68820),
            .I(N__68816));
    InMux I__15060 (
            .O(N__68819),
            .I(N__68808));
    InMux I__15059 (
            .O(N__68816),
            .I(N__68808));
    InMux I__15058 (
            .O(N__68815),
            .I(N__68805));
    InMux I__15057 (
            .O(N__68814),
            .I(N__68800));
    InMux I__15056 (
            .O(N__68813),
            .I(N__68800));
    LocalMux I__15055 (
            .O(N__68808),
            .I(N__68795));
    LocalMux I__15054 (
            .O(N__68805),
            .I(N__68795));
    LocalMux I__15053 (
            .O(N__68800),
            .I(N__68792));
    Span4Mux_v I__15052 (
            .O(N__68795),
            .I(N__68789));
    Span12Mux_s5_v I__15051 (
            .O(N__68792),
            .I(N__68786));
    Span4Mux_h I__15050 (
            .O(N__68789),
            .I(N__68783));
    Odrv12 I__15049 (
            .O(N__68786),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_RNIC2521Z0Z_3 ));
    Odrv4 I__15048 (
            .O(N__68783),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_RNIC2521Z0Z_3 ));
    InMux I__15047 (
            .O(N__68778),
            .I(N__68775));
    LocalMux I__15046 (
            .O(N__68775),
            .I(N__68772));
    Odrv4 I__15045 (
            .O(N__68772),
            .I(\ppm_encoder_1.pulses2countZ0Z_2 ));
    CEMux I__15044 (
            .O(N__68769),
            .I(N__68763));
    CEMux I__15043 (
            .O(N__68768),
            .I(N__68759));
    CEMux I__15042 (
            .O(N__68767),
            .I(N__68755));
    CEMux I__15041 (
            .O(N__68766),
            .I(N__68752));
    LocalMux I__15040 (
            .O(N__68763),
            .I(N__68748));
    CEMux I__15039 (
            .O(N__68762),
            .I(N__68745));
    LocalMux I__15038 (
            .O(N__68759),
            .I(N__68741));
    CEMux I__15037 (
            .O(N__68758),
            .I(N__68738));
    LocalMux I__15036 (
            .O(N__68755),
            .I(N__68735));
    LocalMux I__15035 (
            .O(N__68752),
            .I(N__68732));
    CEMux I__15034 (
            .O(N__68751),
            .I(N__68729));
    Span4Mux_s3_v I__15033 (
            .O(N__68748),
            .I(N__68724));
    LocalMux I__15032 (
            .O(N__68745),
            .I(N__68724));
    CEMux I__15031 (
            .O(N__68744),
            .I(N__68721));
    Span4Mux_s0_v I__15030 (
            .O(N__68741),
            .I(N__68716));
    LocalMux I__15029 (
            .O(N__68738),
            .I(N__68716));
    Span4Mux_v I__15028 (
            .O(N__68735),
            .I(N__68711));
    Span4Mux_v I__15027 (
            .O(N__68732),
            .I(N__68711));
    LocalMux I__15026 (
            .O(N__68729),
            .I(N__68708));
    Span4Mux_h I__15025 (
            .O(N__68724),
            .I(N__68703));
    LocalMux I__15024 (
            .O(N__68721),
            .I(N__68703));
    Span4Mux_v I__15023 (
            .O(N__68716),
            .I(N__68700));
    Span4Mux_h I__15022 (
            .O(N__68711),
            .I(N__68697));
    Span4Mux_v I__15021 (
            .O(N__68708),
            .I(N__68694));
    Span4Mux_v I__15020 (
            .O(N__68703),
            .I(N__68691));
    Span4Mux_h I__15019 (
            .O(N__68700),
            .I(N__68686));
    Span4Mux_h I__15018 (
            .O(N__68697),
            .I(N__68686));
    Span4Mux_h I__15017 (
            .O(N__68694),
            .I(N__68681));
    Span4Mux_h I__15016 (
            .O(N__68691),
            .I(N__68681));
    Odrv4 I__15015 (
            .O(N__68686),
            .I(\ppm_encoder_1.N_295_i_0 ));
    Odrv4 I__15014 (
            .O(N__68681),
            .I(\ppm_encoder_1.N_295_i_0 ));
    InMux I__15013 (
            .O(N__68676),
            .I(N__68671));
    CascadeMux I__15012 (
            .O(N__68675),
            .I(N__68667));
    CascadeMux I__15011 (
            .O(N__68674),
            .I(N__68664));
    LocalMux I__15010 (
            .O(N__68671),
            .I(N__68661));
    CascadeMux I__15009 (
            .O(N__68670),
            .I(N__68657));
    InMux I__15008 (
            .O(N__68667),
            .I(N__68654));
    InMux I__15007 (
            .O(N__68664),
            .I(N__68651));
    Span4Mux_v I__15006 (
            .O(N__68661),
            .I(N__68648));
    InMux I__15005 (
            .O(N__68660),
            .I(N__68645));
    InMux I__15004 (
            .O(N__68657),
            .I(N__68642));
    LocalMux I__15003 (
            .O(N__68654),
            .I(N__68637));
    LocalMux I__15002 (
            .O(N__68651),
            .I(N__68637));
    Span4Mux_h I__15001 (
            .O(N__68648),
            .I(N__68632));
    LocalMux I__15000 (
            .O(N__68645),
            .I(N__68632));
    LocalMux I__14999 (
            .O(N__68642),
            .I(N__68629));
    Span4Mux_h I__14998 (
            .O(N__68637),
            .I(N__68626));
    Span4Mux_v I__14997 (
            .O(N__68632),
            .I(N__68620));
    Span4Mux_h I__14996 (
            .O(N__68629),
            .I(N__68620));
    Span4Mux_v I__14995 (
            .O(N__68626),
            .I(N__68617));
    InMux I__14994 (
            .O(N__68625),
            .I(N__68614));
    Odrv4 I__14993 (
            .O(N__68620),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNIUTMRZ0 ));
    Odrv4 I__14992 (
            .O(N__68617),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNIUTMRZ0 ));
    LocalMux I__14991 (
            .O(N__68614),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNIUTMRZ0 ));
    InMux I__14990 (
            .O(N__68607),
            .I(N__68604));
    LocalMux I__14989 (
            .O(N__68604),
            .I(N__68601));
    Span4Mux_h I__14988 (
            .O(N__68601),
            .I(N__68598));
    Odrv4 I__14987 (
            .O(N__68598),
            .I(\ppm_encoder_1.pulses2count_9_0_0_1_3 ));
    CascadeMux I__14986 (
            .O(N__68595),
            .I(N__68591));
    InMux I__14985 (
            .O(N__68594),
            .I(N__68588));
    InMux I__14984 (
            .O(N__68591),
            .I(N__68585));
    LocalMux I__14983 (
            .O(N__68588),
            .I(N__68581));
    LocalMux I__14982 (
            .O(N__68585),
            .I(N__68578));
    InMux I__14981 (
            .O(N__68584),
            .I(N__68575));
    Span12Mux_s6_v I__14980 (
            .O(N__68581),
            .I(N__68572));
    Span4Mux_h I__14979 (
            .O(N__68578),
            .I(N__68569));
    LocalMux I__14978 (
            .O(N__68575),
            .I(\ppm_encoder_1.throttleZ0Z_3 ));
    Odrv12 I__14977 (
            .O(N__68572),
            .I(\ppm_encoder_1.throttleZ0Z_3 ));
    Odrv4 I__14976 (
            .O(N__68569),
            .I(\ppm_encoder_1.throttleZ0Z_3 ));
    InMux I__14975 (
            .O(N__68562),
            .I(N__68559));
    LocalMux I__14974 (
            .O(N__68559),
            .I(\ppm_encoder_1.pulses2count_9_0_0_3_3 ));
    InMux I__14973 (
            .O(N__68556),
            .I(N__68551));
    InMux I__14972 (
            .O(N__68555),
            .I(N__68548));
    InMux I__14971 (
            .O(N__68554),
            .I(N__68545));
    LocalMux I__14970 (
            .O(N__68551),
            .I(\ppm_encoder_1.counterZ0Z_14 ));
    LocalMux I__14969 (
            .O(N__68548),
            .I(\ppm_encoder_1.counterZ0Z_14 ));
    LocalMux I__14968 (
            .O(N__68545),
            .I(\ppm_encoder_1.counterZ0Z_14 ));
    InMux I__14967 (
            .O(N__68538),
            .I(N__68535));
    LocalMux I__14966 (
            .O(N__68535),
            .I(N__68532));
    Span4Mux_v I__14965 (
            .O(N__68532),
            .I(N__68529));
    Odrv4 I__14964 (
            .O(N__68529),
            .I(\ppm_encoder_1.pulses2countZ0Z_14 ));
    CascadeMux I__14963 (
            .O(N__68526),
            .I(N__68523));
    InMux I__14962 (
            .O(N__68523),
            .I(N__68520));
    LocalMux I__14961 (
            .O(N__68520),
            .I(\ppm_encoder_1.pulses2countZ0Z_15 ));
    CascadeMux I__14960 (
            .O(N__68517),
            .I(N__68513));
    InMux I__14959 (
            .O(N__68516),
            .I(N__68510));
    InMux I__14958 (
            .O(N__68513),
            .I(N__68507));
    LocalMux I__14957 (
            .O(N__68510),
            .I(N__68501));
    LocalMux I__14956 (
            .O(N__68507),
            .I(N__68501));
    InMux I__14955 (
            .O(N__68506),
            .I(N__68498));
    Odrv4 I__14954 (
            .O(N__68501),
            .I(\ppm_encoder_1.counterZ0Z_15 ));
    LocalMux I__14953 (
            .O(N__68498),
            .I(\ppm_encoder_1.counterZ0Z_15 ));
    InMux I__14952 (
            .O(N__68493),
            .I(N__68490));
    LocalMux I__14951 (
            .O(N__68490),
            .I(N__68487));
    Span4Mux_h I__14950 (
            .O(N__68487),
            .I(N__68484));
    Odrv4 I__14949 (
            .O(N__68484),
            .I(\ppm_encoder_1.counter24_0_I_45_c_RNOZ0 ));
    InMux I__14948 (
            .O(N__68481),
            .I(N__68476));
    InMux I__14947 (
            .O(N__68480),
            .I(N__68473));
    InMux I__14946 (
            .O(N__68479),
            .I(N__68470));
    LocalMux I__14945 (
            .O(N__68476),
            .I(N__68467));
    LocalMux I__14944 (
            .O(N__68473),
            .I(N__68464));
    LocalMux I__14943 (
            .O(N__68470),
            .I(\ppm_encoder_1.counterZ0Z_16 ));
    Odrv4 I__14942 (
            .O(N__68467),
            .I(\ppm_encoder_1.counterZ0Z_16 ));
    Odrv4 I__14941 (
            .O(N__68464),
            .I(\ppm_encoder_1.counterZ0Z_16 ));
    InMux I__14940 (
            .O(N__68457),
            .I(N__68452));
    InMux I__14939 (
            .O(N__68456),
            .I(N__68449));
    InMux I__14938 (
            .O(N__68455),
            .I(N__68446));
    LocalMux I__14937 (
            .O(N__68452),
            .I(\ppm_encoder_1.counterZ0Z_3 ));
    LocalMux I__14936 (
            .O(N__68449),
            .I(\ppm_encoder_1.counterZ0Z_3 ));
    LocalMux I__14935 (
            .O(N__68446),
            .I(\ppm_encoder_1.counterZ0Z_3 ));
    CascadeMux I__14934 (
            .O(N__68439),
            .I(N__68436));
    InMux I__14933 (
            .O(N__68436),
            .I(N__68431));
    InMux I__14932 (
            .O(N__68435),
            .I(N__68428));
    InMux I__14931 (
            .O(N__68434),
            .I(N__68425));
    LocalMux I__14930 (
            .O(N__68431),
            .I(N__68422));
    LocalMux I__14929 (
            .O(N__68428),
            .I(N__68419));
    LocalMux I__14928 (
            .O(N__68425),
            .I(\ppm_encoder_1.counterZ0Z_17 ));
    Odrv4 I__14927 (
            .O(N__68422),
            .I(\ppm_encoder_1.counterZ0Z_17 ));
    Odrv4 I__14926 (
            .O(N__68419),
            .I(\ppm_encoder_1.counterZ0Z_17 ));
    InMux I__14925 (
            .O(N__68412),
            .I(N__68407));
    InMux I__14924 (
            .O(N__68411),
            .I(N__68404));
    InMux I__14923 (
            .O(N__68410),
            .I(N__68401));
    LocalMux I__14922 (
            .O(N__68407),
            .I(\ppm_encoder_1.counterZ0Z_2 ));
    LocalMux I__14921 (
            .O(N__68404),
            .I(\ppm_encoder_1.counterZ0Z_2 ));
    LocalMux I__14920 (
            .O(N__68401),
            .I(\ppm_encoder_1.counterZ0Z_2 ));
    InMux I__14919 (
            .O(N__68394),
            .I(N__68391));
    LocalMux I__14918 (
            .O(N__68391),
            .I(N__68388));
    Span4Mux_h I__14917 (
            .O(N__68388),
            .I(N__68385));
    Odrv4 I__14916 (
            .O(N__68385),
            .I(\ppm_encoder_1.un1_PPM_STATE_0_sqmuxa_0_i_a2_18_9 ));
    CascadeMux I__14915 (
            .O(N__68382),
            .I(N__68379));
    InMux I__14914 (
            .O(N__68379),
            .I(N__68376));
    LocalMux I__14913 (
            .O(N__68376),
            .I(N__68373));
    Span4Mux_v I__14912 (
            .O(N__68373),
            .I(N__68370));
    Odrv4 I__14911 (
            .O(N__68370),
            .I(\pid_side.source_pid_1_sqmuxa_1_0_a4_4 ));
    InMux I__14910 (
            .O(N__68367),
            .I(N__68362));
    InMux I__14909 (
            .O(N__68366),
            .I(N__68359));
    InMux I__14908 (
            .O(N__68365),
            .I(N__68356));
    LocalMux I__14907 (
            .O(N__68362),
            .I(N__68353));
    LocalMux I__14906 (
            .O(N__68359),
            .I(N__68348));
    LocalMux I__14905 (
            .O(N__68356),
            .I(N__68348));
    Span4Mux_v I__14904 (
            .O(N__68353),
            .I(N__68345));
    Span4Mux_h I__14903 (
            .O(N__68348),
            .I(N__68342));
    Odrv4 I__14902 (
            .O(N__68345),
            .I(\pid_side.un10lto12 ));
    Odrv4 I__14901 (
            .O(N__68342),
            .I(\pid_side.un10lto12 ));
    CascadeMux I__14900 (
            .O(N__68337),
            .I(N__68333));
    InMux I__14899 (
            .O(N__68336),
            .I(N__68330));
    InMux I__14898 (
            .O(N__68333),
            .I(N__68327));
    LocalMux I__14897 (
            .O(N__68330),
            .I(\pid_side.error_i_acumm_preregZ0Z_21 ));
    LocalMux I__14896 (
            .O(N__68327),
            .I(\pid_side.error_i_acumm_preregZ0Z_21 ));
    InMux I__14895 (
            .O(N__68322),
            .I(N__68319));
    LocalMux I__14894 (
            .O(N__68319),
            .I(N__68314));
    InMux I__14893 (
            .O(N__68318),
            .I(N__68309));
    InMux I__14892 (
            .O(N__68317),
            .I(N__68309));
    Odrv4 I__14891 (
            .O(N__68314),
            .I(\pid_side.error_i_acumm_preregZ0Z_13 ));
    LocalMux I__14890 (
            .O(N__68309),
            .I(\pid_side.error_i_acumm_preregZ0Z_13 ));
    CascadeMux I__14889 (
            .O(N__68304),
            .I(\pid_front.m1_0_03_cascade_ ));
    InMux I__14888 (
            .O(N__68301),
            .I(N__68298));
    LocalMux I__14887 (
            .O(N__68298),
            .I(\pid_front.m1_2_03 ));
    InMux I__14886 (
            .O(N__68295),
            .I(N__68291));
    InMux I__14885 (
            .O(N__68294),
            .I(N__68287));
    LocalMux I__14884 (
            .O(N__68291),
            .I(N__68284));
    InMux I__14883 (
            .O(N__68290),
            .I(N__68281));
    LocalMux I__14882 (
            .O(N__68287),
            .I(N__68277));
    Span4Mux_h I__14881 (
            .O(N__68284),
            .I(N__68274));
    LocalMux I__14880 (
            .O(N__68281),
            .I(N__68271));
    InMux I__14879 (
            .O(N__68280),
            .I(N__68268));
    Span4Mux_v I__14878 (
            .O(N__68277),
            .I(N__68265));
    Sp12to4 I__14877 (
            .O(N__68274),
            .I(N__68260));
    Span12Mux_h I__14876 (
            .O(N__68271),
            .I(N__68260));
    LocalMux I__14875 (
            .O(N__68268),
            .I(pid_side_error_i_reg_9_sn_27));
    Odrv4 I__14874 (
            .O(N__68265),
            .I(pid_side_error_i_reg_9_sn_27));
    Odrv12 I__14873 (
            .O(N__68260),
            .I(pid_side_error_i_reg_9_sn_27));
    InMux I__14872 (
            .O(N__68253),
            .I(N__68250));
    LocalMux I__14871 (
            .O(N__68250),
            .I(N__68246));
    InMux I__14870 (
            .O(N__68249),
            .I(N__68243));
    Sp12to4 I__14869 (
            .O(N__68246),
            .I(N__68240));
    LocalMux I__14868 (
            .O(N__68243),
            .I(N__68237));
    Span12Mux_s10_v I__14867 (
            .O(N__68240),
            .I(N__68234));
    Span4Mux_v I__14866 (
            .O(N__68237),
            .I(N__68231));
    Odrv12 I__14865 (
            .O(N__68234),
            .I(\pid_front.m61_0_bm_0 ));
    Odrv4 I__14864 (
            .O(N__68231),
            .I(\pid_front.m61_0_bm_0 ));
    InMux I__14863 (
            .O(N__68226),
            .I(N__68223));
    LocalMux I__14862 (
            .O(N__68223),
            .I(N__68220));
    Odrv4 I__14861 (
            .O(N__68220),
            .I(\pid_front.error_cry_3_0_c_RNI76FZ0Z08 ));
    CascadeMux I__14860 (
            .O(N__68217),
            .I(N__68214));
    InMux I__14859 (
            .O(N__68214),
            .I(N__68211));
    LocalMux I__14858 (
            .O(N__68211),
            .I(N__68208));
    Span4Mux_h I__14857 (
            .O(N__68208),
            .I(N__68205));
    Odrv4 I__14856 (
            .O(N__68205),
            .I(\pid_front.error_i_regZ0Z_4 ));
    InMux I__14855 (
            .O(N__68202),
            .I(N__68199));
    LocalMux I__14854 (
            .O(N__68199),
            .I(N__68196));
    Span4Mux_v I__14853 (
            .O(N__68196),
            .I(N__68193));
    Odrv4 I__14852 (
            .O(N__68193),
            .I(\pid_side.error_i_reg_9_sn_17 ));
    InMux I__14851 (
            .O(N__68190),
            .I(N__68187));
    LocalMux I__14850 (
            .O(N__68187),
            .I(N__68184));
    Span12Mux_s9_h I__14849 (
            .O(N__68184),
            .I(N__68181));
    Odrv12 I__14848 (
            .O(N__68181),
            .I(\pid_side.error_i_reg_9_sn_25 ));
    CascadeMux I__14847 (
            .O(N__68178),
            .I(N__68175));
    InMux I__14846 (
            .O(N__68175),
            .I(N__68172));
    LocalMux I__14845 (
            .O(N__68172),
            .I(N__68167));
    InMux I__14844 (
            .O(N__68171),
            .I(N__68164));
    CascadeMux I__14843 (
            .O(N__68170),
            .I(N__68161));
    Span4Mux_v I__14842 (
            .O(N__68167),
            .I(N__68158));
    LocalMux I__14841 (
            .O(N__68164),
            .I(N__68155));
    InMux I__14840 (
            .O(N__68161),
            .I(N__68152));
    Span4Mux_h I__14839 (
            .O(N__68158),
            .I(N__68149));
    Span4Mux_h I__14838 (
            .O(N__68155),
            .I(N__68146));
    LocalMux I__14837 (
            .O(N__68152),
            .I(\ppm_encoder_1.aileronZ0Z_3 ));
    Odrv4 I__14836 (
            .O(N__68149),
            .I(\ppm_encoder_1.aileronZ0Z_3 ));
    Odrv4 I__14835 (
            .O(N__68146),
            .I(\ppm_encoder_1.aileronZ0Z_3 ));
    CascadeMux I__14834 (
            .O(N__68139),
            .I(N__68136));
    InMux I__14833 (
            .O(N__68136),
            .I(N__68133));
    LocalMux I__14832 (
            .O(N__68133),
            .I(N__68130));
    Odrv4 I__14831 (
            .O(N__68130),
            .I(\ppm_encoder_1.pulses2countZ0Z_3 ));
    CascadeMux I__14830 (
            .O(N__68127),
            .I(N__68124));
    InMux I__14829 (
            .O(N__68124),
            .I(N__68121));
    LocalMux I__14828 (
            .O(N__68121),
            .I(N__68118));
    Span4Mux_h I__14827 (
            .O(N__68118),
            .I(N__68115));
    Odrv4 I__14826 (
            .O(N__68115),
            .I(\pid_front.error_i_regZ0Z_9 ));
    InMux I__14825 (
            .O(N__68112),
            .I(N__68109));
    LocalMux I__14824 (
            .O(N__68109),
            .I(N__68106));
    Span4Mux_v I__14823 (
            .O(N__68106),
            .I(N__68103));
    Odrv4 I__14822 (
            .O(N__68103),
            .I(\pid_front.error_i_reg_esr_RNO_2Z0Z_25 ));
    CascadeMux I__14821 (
            .O(N__68100),
            .I(\pid_front.error_i_reg_esr_RNO_1Z0Z_25_cascade_ ));
    InMux I__14820 (
            .O(N__68097),
            .I(N__68091));
    InMux I__14819 (
            .O(N__68096),
            .I(N__68091));
    LocalMux I__14818 (
            .O(N__68091),
            .I(N__68088));
    Odrv4 I__14817 (
            .O(N__68088),
            .I(\pid_front.N_93_0 ));
    CascadeMux I__14816 (
            .O(N__68085),
            .I(\pid_front.error_i_reg_9_rn_1_25_cascade_ ));
    InMux I__14815 (
            .O(N__68082),
            .I(N__68079));
    LocalMux I__14814 (
            .O(N__68079),
            .I(N__68076));
    Span4Mux_h I__14813 (
            .O(N__68076),
            .I(N__68073));
    Odrv4 I__14812 (
            .O(N__68073),
            .I(\pid_front.error_i_regZ0Z_25 ));
    InMux I__14811 (
            .O(N__68070),
            .I(N__68067));
    LocalMux I__14810 (
            .O(N__68067),
            .I(\pid_front.N_29_1 ));
    InMux I__14809 (
            .O(N__68064),
            .I(N__68060));
    InMux I__14808 (
            .O(N__68063),
            .I(N__68057));
    LocalMux I__14807 (
            .O(N__68060),
            .I(\pid_front.N_32_0 ));
    LocalMux I__14806 (
            .O(N__68057),
            .I(\pid_front.N_32_0 ));
    CascadeMux I__14805 (
            .O(N__68052),
            .I(N__68049));
    InMux I__14804 (
            .O(N__68049),
            .I(N__68046));
    LocalMux I__14803 (
            .O(N__68046),
            .I(N__68043));
    Span4Mux_h I__14802 (
            .O(N__68043),
            .I(N__68040));
    Odrv4 I__14801 (
            .O(N__68040),
            .I(\pid_front.error_i_regZ0Z_8 ));
    InMux I__14800 (
            .O(N__68037),
            .I(N__68034));
    LocalMux I__14799 (
            .O(N__68034),
            .I(N__68031));
    Odrv12 I__14798 (
            .O(N__68031),
            .I(\pid_front.N_88_0_1 ));
    InMux I__14797 (
            .O(N__68028),
            .I(N__68025));
    LocalMux I__14796 (
            .O(N__68025),
            .I(\pid_front.N_126_1 ));
    InMux I__14795 (
            .O(N__68022),
            .I(N__68019));
    LocalMux I__14794 (
            .O(N__68019),
            .I(N__68016));
    Span4Mux_h I__14793 (
            .O(N__68016),
            .I(N__68013));
    Odrv4 I__14792 (
            .O(N__68013),
            .I(\pid_front.N_116_0 ));
    CascadeMux I__14791 (
            .O(N__68010),
            .I(\pid_front.error_i_reg_9_rn_1_13_cascade_ ));
    InMux I__14790 (
            .O(N__68007),
            .I(N__68004));
    LocalMux I__14789 (
            .O(N__68004),
            .I(\pid_front.N_127 ));
    CascadeMux I__14788 (
            .O(N__68001),
            .I(N__67998));
    InMux I__14787 (
            .O(N__67998),
            .I(N__67995));
    LocalMux I__14786 (
            .O(N__67995),
            .I(N__67992));
    Odrv4 I__14785 (
            .O(N__67992),
            .I(\pid_front.error_i_regZ0Z_13 ));
    InMux I__14784 (
            .O(N__67989),
            .I(N__67983));
    InMux I__14783 (
            .O(N__67988),
            .I(N__67983));
    LocalMux I__14782 (
            .O(N__67983),
            .I(N__67980));
    Span4Mux_v I__14781 (
            .O(N__67980),
            .I(N__67977));
    Odrv4 I__14780 (
            .O(N__67977),
            .I(\pid_front.error_i_regZ0Z_27 ));
    CascadeMux I__14779 (
            .O(N__67974),
            .I(\pid_front.m7_2_03_cascade_ ));
    CascadeMux I__14778 (
            .O(N__67971),
            .I(\pid_front.error_i_reg_9_rn_0_19_cascade_ ));
    InMux I__14777 (
            .O(N__67968),
            .I(N__67965));
    LocalMux I__14776 (
            .O(N__67965),
            .I(N__67962));
    Span4Mux_h I__14775 (
            .O(N__67962),
            .I(N__67959));
    Odrv4 I__14774 (
            .O(N__67959),
            .I(\pid_front.error_i_regZ0Z_19 ));
    CascadeMux I__14773 (
            .O(N__67956),
            .I(pid_front_error_i_reg_9_sn_19_cascade_));
    InMux I__14772 (
            .O(N__67953),
            .I(N__67950));
    LocalMux I__14771 (
            .O(N__67950),
            .I(\pid_front.error_i_reg_esr_RNO_2Z0Z_19 ));
    InMux I__14770 (
            .O(N__67947),
            .I(N__67944));
    LocalMux I__14769 (
            .O(N__67944),
            .I(N__67941));
    Span4Mux_h I__14768 (
            .O(N__67941),
            .I(N__67938));
    Odrv4 I__14767 (
            .O(N__67938),
            .I(\pid_front.N_55_0 ));
    InMux I__14766 (
            .O(N__67935),
            .I(N__67932));
    LocalMux I__14765 (
            .O(N__67932),
            .I(N__67929));
    Span4Mux_h I__14764 (
            .O(N__67929),
            .I(N__67925));
    InMux I__14763 (
            .O(N__67928),
            .I(N__67922));
    Odrv4 I__14762 (
            .O(N__67925),
            .I(\pid_front.N_110 ));
    LocalMux I__14761 (
            .O(N__67922),
            .I(\pid_front.N_110 ));
    CascadeMux I__14760 (
            .O(N__67917),
            .I(N__67914));
    InMux I__14759 (
            .O(N__67914),
            .I(N__67911));
    LocalMux I__14758 (
            .O(N__67911),
            .I(N__67908));
    Span4Mux_h I__14757 (
            .O(N__67908),
            .I(N__67905));
    Odrv4 I__14756 (
            .O(N__67905),
            .I(\pid_front.error_i_regZ0Z_6 ));
    InMux I__14755 (
            .O(N__67902),
            .I(N__67899));
    LocalMux I__14754 (
            .O(N__67899),
            .I(\pid_front.N_103_0 ));
    CascadeMux I__14753 (
            .O(N__67896),
            .I(N__67893));
    InMux I__14752 (
            .O(N__67893),
            .I(N__67890));
    LocalMux I__14751 (
            .O(N__67890),
            .I(N__67887));
    Span4Mux_h I__14750 (
            .O(N__67887),
            .I(N__67884));
    Odrv4 I__14749 (
            .O(N__67884),
            .I(\pid_front.error_i_regZ0Z_7 ));
    CascadeMux I__14748 (
            .O(N__67881),
            .I(\pid_side.error_i_reg_9_rn_1_12_cascade_ ));
    InMux I__14747 (
            .O(N__67878),
            .I(N__67875));
    LocalMux I__14746 (
            .O(N__67875),
            .I(\pid_side.N_129 ));
    CascadeMux I__14745 (
            .O(N__67872),
            .I(N__67869));
    InMux I__14744 (
            .O(N__67869),
            .I(N__67866));
    LocalMux I__14743 (
            .O(N__67866),
            .I(N__67863));
    Span12Mux_s9_h I__14742 (
            .O(N__67863),
            .I(N__67860));
    Odrv12 I__14741 (
            .O(N__67860),
            .I(\pid_side.error_i_regZ0Z_12 ));
    InMux I__14740 (
            .O(N__67857),
            .I(N__67854));
    LocalMux I__14739 (
            .O(N__67854),
            .I(N__67851));
    Span4Mux_s2_h I__14738 (
            .O(N__67851),
            .I(N__67847));
    InMux I__14737 (
            .O(N__67850),
            .I(N__67842));
    Span4Mux_v I__14736 (
            .O(N__67847),
            .I(N__67839));
    InMux I__14735 (
            .O(N__67846),
            .I(N__67835));
    InMux I__14734 (
            .O(N__67845),
            .I(N__67832));
    LocalMux I__14733 (
            .O(N__67842),
            .I(N__67829));
    Span4Mux_h I__14732 (
            .O(N__67839),
            .I(N__67826));
    InMux I__14731 (
            .O(N__67838),
            .I(N__67823));
    LocalMux I__14730 (
            .O(N__67835),
            .I(N__67816));
    LocalMux I__14729 (
            .O(N__67832),
            .I(N__67816));
    Span12Mux_s9_v I__14728 (
            .O(N__67829),
            .I(N__67816));
    Span4Mux_h I__14727 (
            .O(N__67826),
            .I(N__67813));
    LocalMux I__14726 (
            .O(N__67823),
            .I(\pid_front.error_4 ));
    Odrv12 I__14725 (
            .O(N__67816),
            .I(\pid_front.error_4 ));
    Odrv4 I__14724 (
            .O(N__67813),
            .I(\pid_front.error_4 ));
    InMux I__14723 (
            .O(N__67806),
            .I(N__67802));
    InMux I__14722 (
            .O(N__67805),
            .I(N__67799));
    LocalMux I__14721 (
            .O(N__67802),
            .I(N__67796));
    LocalMux I__14720 (
            .O(N__67799),
            .I(N__67793));
    Span4Mux_v I__14719 (
            .O(N__67796),
            .I(N__67790));
    Span12Mux_v I__14718 (
            .O(N__67793),
            .I(N__67785));
    Span4Mux_h I__14717 (
            .O(N__67790),
            .I(N__67781));
    InMux I__14716 (
            .O(N__67789),
            .I(N__67778));
    InMux I__14715 (
            .O(N__67788),
            .I(N__67775));
    Span12Mux_h I__14714 (
            .O(N__67785),
            .I(N__67772));
    InMux I__14713 (
            .O(N__67784),
            .I(N__67769));
    Span4Mux_h I__14712 (
            .O(N__67781),
            .I(N__67762));
    LocalMux I__14711 (
            .O(N__67778),
            .I(N__67762));
    LocalMux I__14710 (
            .O(N__67775),
            .I(N__67762));
    Odrv12 I__14709 (
            .O(N__67772),
            .I(\pid_front.error_5 ));
    LocalMux I__14708 (
            .O(N__67769),
            .I(\pid_front.error_5 ));
    Odrv4 I__14707 (
            .O(N__67762),
            .I(\pid_front.error_5 ));
    InMux I__14706 (
            .O(N__67755),
            .I(N__67751));
    InMux I__14705 (
            .O(N__67754),
            .I(N__67748));
    LocalMux I__14704 (
            .O(N__67751),
            .I(N__67743));
    LocalMux I__14703 (
            .O(N__67748),
            .I(N__67740));
    CascadeMux I__14702 (
            .O(N__67747),
            .I(N__67736));
    CascadeMux I__14701 (
            .O(N__67746),
            .I(N__67733));
    Span4Mux_h I__14700 (
            .O(N__67743),
            .I(N__67730));
    Span4Mux_s1_h I__14699 (
            .O(N__67740),
            .I(N__67727));
    InMux I__14698 (
            .O(N__67739),
            .I(N__67723));
    InMux I__14697 (
            .O(N__67736),
            .I(N__67718));
    InMux I__14696 (
            .O(N__67733),
            .I(N__67718));
    Span4Mux_v I__14695 (
            .O(N__67730),
            .I(N__67715));
    Span4Mux_h I__14694 (
            .O(N__67727),
            .I(N__67712));
    InMux I__14693 (
            .O(N__67726),
            .I(N__67709));
    LocalMux I__14692 (
            .O(N__67723),
            .I(N__67706));
    LocalMux I__14691 (
            .O(N__67718),
            .I(N__67703));
    Span4Mux_h I__14690 (
            .O(N__67715),
            .I(N__67700));
    Span4Mux_h I__14689 (
            .O(N__67712),
            .I(N__67697));
    LocalMux I__14688 (
            .O(N__67709),
            .I(N__67686));
    Span4Mux_v I__14687 (
            .O(N__67706),
            .I(N__67686));
    Span4Mux_h I__14686 (
            .O(N__67703),
            .I(N__67686));
    Span4Mux_h I__14685 (
            .O(N__67700),
            .I(N__67686));
    Span4Mux_v I__14684 (
            .O(N__67697),
            .I(N__67686));
    Odrv4 I__14683 (
            .O(N__67686),
            .I(\pid_front.error_6 ));
    InMux I__14682 (
            .O(N__67683),
            .I(N__67679));
    InMux I__14681 (
            .O(N__67682),
            .I(N__67676));
    LocalMux I__14680 (
            .O(N__67679),
            .I(N__67673));
    LocalMux I__14679 (
            .O(N__67676),
            .I(N__67670));
    Span4Mux_s3_h I__14678 (
            .O(N__67673),
            .I(N__67664));
    Span4Mux_s2_h I__14677 (
            .O(N__67670),
            .I(N__67659));
    InMux I__14676 (
            .O(N__67669),
            .I(N__67656));
    InMux I__14675 (
            .O(N__67668),
            .I(N__67651));
    InMux I__14674 (
            .O(N__67667),
            .I(N__67651));
    Span4Mux_v I__14673 (
            .O(N__67664),
            .I(N__67648));
    InMux I__14672 (
            .O(N__67663),
            .I(N__67645));
    InMux I__14671 (
            .O(N__67662),
            .I(N__67642));
    Span4Mux_h I__14670 (
            .O(N__67659),
            .I(N__67639));
    LocalMux I__14669 (
            .O(N__67656),
            .I(N__67635));
    LocalMux I__14668 (
            .O(N__67651),
            .I(N__67632));
    Span4Mux_h I__14667 (
            .O(N__67648),
            .I(N__67629));
    LocalMux I__14666 (
            .O(N__67645),
            .I(N__67622));
    LocalMux I__14665 (
            .O(N__67642),
            .I(N__67622));
    Span4Mux_h I__14664 (
            .O(N__67639),
            .I(N__67622));
    InMux I__14663 (
            .O(N__67638),
            .I(N__67619));
    Span4Mux_h I__14662 (
            .O(N__67635),
            .I(N__67616));
    Span4Mux_h I__14661 (
            .O(N__67632),
            .I(N__67609));
    Span4Mux_h I__14660 (
            .O(N__67629),
            .I(N__67609));
    Span4Mux_v I__14659 (
            .O(N__67622),
            .I(N__67609));
    LocalMux I__14658 (
            .O(N__67619),
            .I(\pid_front.error_7 ));
    Odrv4 I__14657 (
            .O(N__67616),
            .I(\pid_front.error_7 ));
    Odrv4 I__14656 (
            .O(N__67609),
            .I(\pid_front.error_7 ));
    InMux I__14655 (
            .O(N__67602),
            .I(N__67599));
    LocalMux I__14654 (
            .O(N__67599),
            .I(\pid_front.N_9_1 ));
    CascadeMux I__14653 (
            .O(N__67596),
            .I(\pid_front.error_cry_1_0_c_RNIDPRQ1Z0Z_0_cascade_ ));
    InMux I__14652 (
            .O(N__67593),
            .I(N__67590));
    LocalMux I__14651 (
            .O(N__67590),
            .I(\pid_front.error_cry_1_0_c_RNIDPRQZ0Z1 ));
    InMux I__14650 (
            .O(N__67587),
            .I(N__67583));
    InMux I__14649 (
            .O(N__67586),
            .I(N__67580));
    LocalMux I__14648 (
            .O(N__67583),
            .I(N__67574));
    LocalMux I__14647 (
            .O(N__67580),
            .I(N__67574));
    InMux I__14646 (
            .O(N__67579),
            .I(N__67571));
    Span4Mux_v I__14645 (
            .O(N__67574),
            .I(N__67566));
    LocalMux I__14644 (
            .O(N__67571),
            .I(N__67563));
    InMux I__14643 (
            .O(N__67570),
            .I(N__67558));
    InMux I__14642 (
            .O(N__67569),
            .I(N__67558));
    Span4Mux_v I__14641 (
            .O(N__67566),
            .I(N__67555));
    Span4Mux_v I__14640 (
            .O(N__67563),
            .I(N__67550));
    LocalMux I__14639 (
            .O(N__67558),
            .I(N__67550));
    Span4Mux_v I__14638 (
            .O(N__67555),
            .I(N__67547));
    Span4Mux_h I__14637 (
            .O(N__67550),
            .I(N__67544));
    Odrv4 I__14636 (
            .O(N__67547),
            .I(xy_ki_fast_3));
    Odrv4 I__14635 (
            .O(N__67544),
            .I(xy_ki_fast_3));
    CascadeMux I__14634 (
            .O(N__67539),
            .I(\pid_front.N_39_0_cascade_ ));
    CascadeMux I__14633 (
            .O(N__67536),
            .I(\pid_front.m53_0_ns_1_cascade_ ));
    InMux I__14632 (
            .O(N__67533),
            .I(N__67529));
    InMux I__14631 (
            .O(N__67532),
            .I(N__67526));
    LocalMux I__14630 (
            .O(N__67529),
            .I(N__67523));
    LocalMux I__14629 (
            .O(N__67526),
            .I(N__67520));
    Span4Mux_v I__14628 (
            .O(N__67523),
            .I(N__67516));
    Span4Mux_v I__14627 (
            .O(N__67520),
            .I(N__67513));
    InMux I__14626 (
            .O(N__67519),
            .I(N__67510));
    Span4Mux_h I__14625 (
            .O(N__67516),
            .I(N__67507));
    Sp12to4 I__14624 (
            .O(N__67513),
            .I(N__67502));
    LocalMux I__14623 (
            .O(N__67510),
            .I(N__67502));
    Odrv4 I__14622 (
            .O(N__67507),
            .I(\pid_front.state_ns_0 ));
    Odrv12 I__14621 (
            .O(N__67502),
            .I(\pid_front.state_ns_0 ));
    CascadeMux I__14620 (
            .O(N__67497),
            .I(\pid_front.N_54_0_cascade_ ));
    CascadeMux I__14619 (
            .O(N__67494),
            .I(N__67491));
    InMux I__14618 (
            .O(N__67491),
            .I(N__67488));
    LocalMux I__14617 (
            .O(N__67488),
            .I(N__67484));
    InMux I__14616 (
            .O(N__67487),
            .I(N__67481));
    Span4Mux_h I__14615 (
            .O(N__67484),
            .I(N__67478));
    LocalMux I__14614 (
            .O(N__67481),
            .I(\pid_front.error_i_regZ0Z_11 ));
    Odrv4 I__14613 (
            .O(N__67478),
            .I(\pid_front.error_i_regZ0Z_11 ));
    InMux I__14612 (
            .O(N__67473),
            .I(N__67470));
    LocalMux I__14611 (
            .O(N__67470),
            .I(\pid_front.N_54_0 ));
    InMux I__14610 (
            .O(N__67467),
            .I(N__67464));
    LocalMux I__14609 (
            .O(N__67464),
            .I(\pid_side.error_i_reg_9_rn_1_17 ));
    InMux I__14608 (
            .O(N__67461),
            .I(N__67458));
    LocalMux I__14607 (
            .O(N__67458),
            .I(N__67455));
    Odrv12 I__14606 (
            .O(N__67455),
            .I(\pid_side.error_i_regZ0Z_17 ));
    InMux I__14605 (
            .O(N__67452),
            .I(N__67449));
    LocalMux I__14604 (
            .O(N__67449),
            .I(\pid_side.error_i_reg_9_rn_1_25 ));
    InMux I__14603 (
            .O(N__67446),
            .I(N__67443));
    LocalMux I__14602 (
            .O(N__67443),
            .I(N__67440));
    Span4Mux_v I__14601 (
            .O(N__67440),
            .I(N__67437));
    Odrv4 I__14600 (
            .O(N__67437),
            .I(\pid_side.error_i_regZ0Z_25 ));
    InMux I__14599 (
            .O(N__67434),
            .I(N__67431));
    LocalMux I__14598 (
            .O(N__67431),
            .I(N__67427));
    InMux I__14597 (
            .O(N__67430),
            .I(N__67424));
    Span4Mux_h I__14596 (
            .O(N__67427),
            .I(N__67421));
    LocalMux I__14595 (
            .O(N__67424),
            .I(\pid_side.m61_0_bmZ0 ));
    Odrv4 I__14594 (
            .O(N__67421),
            .I(\pid_side.m61_0_bmZ0 ));
    InMux I__14593 (
            .O(N__67416),
            .I(N__67412));
    InMux I__14592 (
            .O(N__67415),
            .I(N__67409));
    LocalMux I__14591 (
            .O(N__67412),
            .I(N__67406));
    LocalMux I__14590 (
            .O(N__67409),
            .I(N__67401));
    Span4Mux_v I__14589 (
            .O(N__67406),
            .I(N__67398));
    InMux I__14588 (
            .O(N__67405),
            .I(N__67392));
    InMux I__14587 (
            .O(N__67404),
            .I(N__67392));
    Span4Mux_s3_h I__14586 (
            .O(N__67401),
            .I(N__67387));
    Span4Mux_h I__14585 (
            .O(N__67398),
            .I(N__67384));
    CascadeMux I__14584 (
            .O(N__67397),
            .I(N__67381));
    LocalMux I__14583 (
            .O(N__67392),
            .I(N__67377));
    InMux I__14582 (
            .O(N__67391),
            .I(N__67374));
    InMux I__14581 (
            .O(N__67390),
            .I(N__67371));
    Span4Mux_h I__14580 (
            .O(N__67387),
            .I(N__67368));
    Span4Mux_h I__14579 (
            .O(N__67384),
            .I(N__67365));
    InMux I__14578 (
            .O(N__67381),
            .I(N__67360));
    InMux I__14577 (
            .O(N__67380),
            .I(N__67360));
    Span4Mux_v I__14576 (
            .O(N__67377),
            .I(N__67357));
    LocalMux I__14575 (
            .O(N__67374),
            .I(N__67350));
    LocalMux I__14574 (
            .O(N__67371),
            .I(N__67350));
    Span4Mux_h I__14573 (
            .O(N__67368),
            .I(N__67350));
    Span4Mux_h I__14572 (
            .O(N__67365),
            .I(N__67347));
    LocalMux I__14571 (
            .O(N__67360),
            .I(\pid_front.error_11 ));
    Odrv4 I__14570 (
            .O(N__67357),
            .I(\pid_front.error_11 ));
    Odrv4 I__14569 (
            .O(N__67350),
            .I(\pid_front.error_11 ));
    Odrv4 I__14568 (
            .O(N__67347),
            .I(\pid_front.error_11 ));
    InMux I__14567 (
            .O(N__67338),
            .I(N__67335));
    LocalMux I__14566 (
            .O(N__67335),
            .I(N__67331));
    InMux I__14565 (
            .O(N__67334),
            .I(N__67327));
    Span4Mux_s2_h I__14564 (
            .O(N__67331),
            .I(N__67324));
    CascadeMux I__14563 (
            .O(N__67330),
            .I(N__67321));
    LocalMux I__14562 (
            .O(N__67327),
            .I(N__67317));
    Span4Mux_h I__14561 (
            .O(N__67324),
            .I(N__67314));
    InMux I__14560 (
            .O(N__67321),
            .I(N__67308));
    InMux I__14559 (
            .O(N__67320),
            .I(N__67308));
    Span4Mux_s3_h I__14558 (
            .O(N__67317),
            .I(N__67302));
    Span4Mux_v I__14557 (
            .O(N__67314),
            .I(N__67299));
    InMux I__14556 (
            .O(N__67313),
            .I(N__67296));
    LocalMux I__14555 (
            .O(N__67308),
            .I(N__67293));
    InMux I__14554 (
            .O(N__67307),
            .I(N__67290));
    InMux I__14553 (
            .O(N__67306),
            .I(N__67287));
    InMux I__14552 (
            .O(N__67305),
            .I(N__67284));
    Span4Mux_h I__14551 (
            .O(N__67302),
            .I(N__67281));
    Span4Mux_h I__14550 (
            .O(N__67299),
            .I(N__67278));
    LocalMux I__14549 (
            .O(N__67296),
            .I(N__67273));
    Span4Mux_v I__14548 (
            .O(N__67293),
            .I(N__67273));
    LocalMux I__14547 (
            .O(N__67290),
            .I(N__67262));
    LocalMux I__14546 (
            .O(N__67287),
            .I(N__67262));
    LocalMux I__14545 (
            .O(N__67284),
            .I(N__67262));
    Span4Mux_h I__14544 (
            .O(N__67281),
            .I(N__67262));
    Span4Mux_h I__14543 (
            .O(N__67278),
            .I(N__67262));
    Odrv4 I__14542 (
            .O(N__67273),
            .I(\pid_front.error_10 ));
    Odrv4 I__14541 (
            .O(N__67262),
            .I(\pid_front.error_10 ));
    InMux I__14540 (
            .O(N__67257),
            .I(N__67254));
    LocalMux I__14539 (
            .O(N__67254),
            .I(N__67250));
    InMux I__14538 (
            .O(N__67253),
            .I(N__67247));
    Span4Mux_v I__14537 (
            .O(N__67250),
            .I(N__67244));
    LocalMux I__14536 (
            .O(N__67247),
            .I(N__67241));
    Span4Mux_h I__14535 (
            .O(N__67244),
            .I(N__67238));
    Span4Mux_s3_h I__14534 (
            .O(N__67241),
            .I(N__67234));
    Span4Mux_h I__14533 (
            .O(N__67238),
            .I(N__67230));
    InMux I__14532 (
            .O(N__67237),
            .I(N__67227));
    Span4Mux_h I__14531 (
            .O(N__67234),
            .I(N__67224));
    InMux I__14530 (
            .O(N__67233),
            .I(N__67221));
    Span4Mux_h I__14529 (
            .O(N__67230),
            .I(N__67216));
    LocalMux I__14528 (
            .O(N__67227),
            .I(N__67216));
    Span4Mux_h I__14527 (
            .O(N__67224),
            .I(N__67209));
    LocalMux I__14526 (
            .O(N__67221),
            .I(N__67209));
    Span4Mux_h I__14525 (
            .O(N__67216),
            .I(N__67206));
    InMux I__14524 (
            .O(N__67215),
            .I(N__67201));
    InMux I__14523 (
            .O(N__67214),
            .I(N__67201));
    Odrv4 I__14522 (
            .O(N__67209),
            .I(\pid_front.error_13 ));
    Odrv4 I__14521 (
            .O(N__67206),
            .I(\pid_front.error_13 ));
    LocalMux I__14520 (
            .O(N__67201),
            .I(\pid_front.error_13 ));
    CascadeMux I__14519 (
            .O(N__67194),
            .I(\pid_front.g0_15_1_cascade_ ));
    InMux I__14518 (
            .O(N__67191),
            .I(N__67188));
    LocalMux I__14517 (
            .O(N__67188),
            .I(N__67185));
    Span4Mux_v I__14516 (
            .O(N__67185),
            .I(N__67180));
    InMux I__14515 (
            .O(N__67184),
            .I(N__67176));
    InMux I__14514 (
            .O(N__67183),
            .I(N__67173));
    Span4Mux_h I__14513 (
            .O(N__67180),
            .I(N__67170));
    InMux I__14512 (
            .O(N__67179),
            .I(N__67167));
    LocalMux I__14511 (
            .O(N__67176),
            .I(N__67160));
    LocalMux I__14510 (
            .O(N__67173),
            .I(N__67157));
    Span4Mux_h I__14509 (
            .O(N__67170),
            .I(N__67154));
    LocalMux I__14508 (
            .O(N__67167),
            .I(N__67151));
    InMux I__14507 (
            .O(N__67166),
            .I(N__67146));
    InMux I__14506 (
            .O(N__67165),
            .I(N__67146));
    InMux I__14505 (
            .O(N__67164),
            .I(N__67141));
    InMux I__14504 (
            .O(N__67163),
            .I(N__67141));
    Span12Mux_s8_v I__14503 (
            .O(N__67160),
            .I(N__67138));
    Span4Mux_h I__14502 (
            .O(N__67157),
            .I(N__67133));
    Span4Mux_h I__14501 (
            .O(N__67154),
            .I(N__67133));
    Odrv4 I__14500 (
            .O(N__67151),
            .I(\pid_front.error_12 ));
    LocalMux I__14499 (
            .O(N__67146),
            .I(\pid_front.error_12 ));
    LocalMux I__14498 (
            .O(N__67141),
            .I(\pid_front.error_12 ));
    Odrv12 I__14497 (
            .O(N__67138),
            .I(\pid_front.error_12 ));
    Odrv4 I__14496 (
            .O(N__67133),
            .I(\pid_front.error_12 ));
    InMux I__14495 (
            .O(N__67122),
            .I(N__67119));
    LocalMux I__14494 (
            .O(N__67119),
            .I(\pid_side.N_9_1_0 ));
    InMux I__14493 (
            .O(N__67116),
            .I(N__67112));
    InMux I__14492 (
            .O(N__67115),
            .I(N__67109));
    LocalMux I__14491 (
            .O(N__67112),
            .I(N__67104));
    LocalMux I__14490 (
            .O(N__67109),
            .I(N__67101));
    InMux I__14489 (
            .O(N__67108),
            .I(N__67098));
    CascadeMux I__14488 (
            .O(N__67107),
            .I(N__67095));
    Span4Mux_v I__14487 (
            .O(N__67104),
            .I(N__67092));
    Span4Mux_h I__14486 (
            .O(N__67101),
            .I(N__67087));
    LocalMux I__14485 (
            .O(N__67098),
            .I(N__67087));
    InMux I__14484 (
            .O(N__67095),
            .I(N__67084));
    Span4Mux_v I__14483 (
            .O(N__67092),
            .I(N__67081));
    Span4Mux_v I__14482 (
            .O(N__67087),
            .I(N__67078));
    LocalMux I__14481 (
            .O(N__67084),
            .I(\pid_side.N_15_0 ));
    Odrv4 I__14480 (
            .O(N__67081),
            .I(\pid_side.N_15_0 ));
    Odrv4 I__14479 (
            .O(N__67078),
            .I(\pid_side.N_15_0 ));
    InMux I__14478 (
            .O(N__67071),
            .I(N__67068));
    LocalMux I__14477 (
            .O(N__67068),
            .I(N__67062));
    InMux I__14476 (
            .O(N__67067),
            .I(N__67055));
    InMux I__14475 (
            .O(N__67066),
            .I(N__67055));
    InMux I__14474 (
            .O(N__67065),
            .I(N__67055));
    Odrv4 I__14473 (
            .O(N__67062),
            .I(\pid_side.N_28_1 ));
    LocalMux I__14472 (
            .O(N__67055),
            .I(\pid_side.N_28_1 ));
    CascadeMux I__14471 (
            .O(N__67050),
            .I(\pid_side.N_60_0_cascade_ ));
    InMux I__14470 (
            .O(N__67047),
            .I(N__67044));
    LocalMux I__14469 (
            .O(N__67044),
            .I(N__67040));
    InMux I__14468 (
            .O(N__67043),
            .I(N__67037));
    Span4Mux_v I__14467 (
            .O(N__67040),
            .I(N__67034));
    LocalMux I__14466 (
            .O(N__67037),
            .I(\pid_side.N_11_0 ));
    Odrv4 I__14465 (
            .O(N__67034),
            .I(\pid_side.N_11_0 ));
    InMux I__14464 (
            .O(N__67029),
            .I(N__67026));
    LocalMux I__14463 (
            .O(N__67026),
            .I(N__67023));
    Span4Mux_h I__14462 (
            .O(N__67023),
            .I(N__67020));
    Span4Mux_v I__14461 (
            .O(N__67020),
            .I(N__67016));
    InMux I__14460 (
            .O(N__67019),
            .I(N__67013));
    Odrv4 I__14459 (
            .O(N__67016),
            .I(\pid_side.N_12_1 ));
    LocalMux I__14458 (
            .O(N__67013),
            .I(\pid_side.N_12_1 ));
    CascadeMux I__14457 (
            .O(N__67008),
            .I(\pid_side.N_12_1_cascade_ ));
    CascadeMux I__14456 (
            .O(N__67005),
            .I(\pid_side.N_93_0_cascade_ ));
    CascadeMux I__14455 (
            .O(N__67002),
            .I(\pid_side.un4_error_i_reg_35_am_1_cascade_ ));
    InMux I__14454 (
            .O(N__66999),
            .I(N__66996));
    LocalMux I__14453 (
            .O(N__66996),
            .I(\pid_side.error_i_reg_esr_RNO_2_0_25 ));
    InMux I__14452 (
            .O(N__66993),
            .I(N__66990));
    LocalMux I__14451 (
            .O(N__66990),
            .I(\pid_side.N_93_0 ));
    CascadeMux I__14450 (
            .O(N__66987),
            .I(N__66984));
    InMux I__14449 (
            .O(N__66984),
            .I(N__66981));
    LocalMux I__14448 (
            .O(N__66981),
            .I(N__66978));
    Span4Mux_v I__14447 (
            .O(N__66978),
            .I(N__66975));
    Odrv4 I__14446 (
            .O(N__66975),
            .I(\pid_side.error_i_regZ0Z_9 ));
    CascadeMux I__14445 (
            .O(N__66972),
            .I(pid_side_N_166_cascade_));
    InMux I__14444 (
            .O(N__66969),
            .I(N__66966));
    LocalMux I__14443 (
            .O(N__66966),
            .I(N__66963));
    Odrv4 I__14442 (
            .O(N__66963),
            .I(\pid_side.error_cry_0_c_RNI94FZ0Z58 ));
    CascadeMux I__14441 (
            .O(N__66960),
            .I(N__66957));
    InMux I__14440 (
            .O(N__66957),
            .I(N__66954));
    LocalMux I__14439 (
            .O(N__66954),
            .I(N__66951));
    Odrv12 I__14438 (
            .O(N__66951),
            .I(\pid_side.error_i_regZ0Z_4 ));
    CascadeMux I__14437 (
            .O(N__66948),
            .I(\pid_side.m32_0_ns_1_cascade_ ));
    CascadeMux I__14436 (
            .O(N__66945),
            .I(\pid_side.N_89_i_cascade_ ));
    InMux I__14435 (
            .O(N__66942),
            .I(N__66939));
    LocalMux I__14434 (
            .O(N__66939),
            .I(N__66936));
    Span12Mux_v I__14433 (
            .O(N__66936),
            .I(N__66933));
    Odrv12 I__14432 (
            .O(N__66933),
            .I(\pid_side.state_ns_0 ));
    CascadeMux I__14431 (
            .O(N__66930),
            .I(N__66927));
    InMux I__14430 (
            .O(N__66927),
            .I(N__66923));
    InMux I__14429 (
            .O(N__66926),
            .I(N__66920));
    LocalMux I__14428 (
            .O(N__66923),
            .I(N__66917));
    LocalMux I__14427 (
            .O(N__66920),
            .I(\pid_side.error_i_regZ0Z_8 ));
    Odrv4 I__14426 (
            .O(N__66917),
            .I(\pid_side.error_i_regZ0Z_8 ));
    CascadeMux I__14425 (
            .O(N__66912),
            .I(\pid_side.N_22_0_cascade_ ));
    InMux I__14424 (
            .O(N__66909),
            .I(N__66903));
    InMux I__14423 (
            .O(N__66908),
            .I(N__66903));
    LocalMux I__14422 (
            .O(N__66903),
            .I(\pid_side.N_22_0 ));
    CascadeMux I__14421 (
            .O(N__66900),
            .I(\pid_side.error_i_reg_esr_RNO_4Z0Z_16_cascade_ ));
    InMux I__14420 (
            .O(N__66897),
            .I(N__66894));
    LocalMux I__14419 (
            .O(N__66894),
            .I(\pid_side.error_i_reg_esr_RNO_3Z0Z_16 ));
    InMux I__14418 (
            .O(N__66891),
            .I(N__66888));
    LocalMux I__14417 (
            .O(N__66888),
            .I(N__66885));
    Span4Mux_v I__14416 (
            .O(N__66885),
            .I(N__66882));
    Odrv4 I__14415 (
            .O(N__66882),
            .I(\pid_side.m20_2_03_0 ));
    InMux I__14414 (
            .O(N__66879),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_21 ));
    InMux I__14413 (
            .O(N__66876),
            .I(N__66873));
    LocalMux I__14412 (
            .O(N__66873),
            .I(\pid_side.error_i_regZ0Z_23 ));
    InMux I__14411 (
            .O(N__66870),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_22 ));
    InMux I__14410 (
            .O(N__66867),
            .I(bfn_16_16_0_));
    InMux I__14409 (
            .O(N__66864),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_24 ));
    CascadeMux I__14408 (
            .O(N__66861),
            .I(N__66858));
    InMux I__14407 (
            .O(N__66858),
            .I(N__66855));
    LocalMux I__14406 (
            .O(N__66855),
            .I(N__66852));
    Span4Mux_v I__14405 (
            .O(N__66852),
            .I(N__66849));
    Odrv4 I__14404 (
            .O(N__66849),
            .I(\pid_side.error_i_regZ0Z_26 ));
    InMux I__14403 (
            .O(N__66846),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_25 ));
    InMux I__14402 (
            .O(N__66843),
            .I(N__66838));
    InMux I__14401 (
            .O(N__66842),
            .I(N__66833));
    InMux I__14400 (
            .O(N__66841),
            .I(N__66833));
    LocalMux I__14399 (
            .O(N__66838),
            .I(N__66830));
    LocalMux I__14398 (
            .O(N__66833),
            .I(N__66827));
    Odrv12 I__14397 (
            .O(N__66830),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_26_c_RNI0LUS ));
    Odrv4 I__14396 (
            .O(N__66827),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_26_c_RNI0LUS ));
    InMux I__14395 (
            .O(N__66822),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_26 ));
    InMux I__14394 (
            .O(N__66819),
            .I(N__66813));
    InMux I__14393 (
            .O(N__66818),
            .I(N__66813));
    LocalMux I__14392 (
            .O(N__66813),
            .I(N__66810));
    Odrv4 I__14391 (
            .O(N__66810),
            .I(\pid_side.error_i_regZ0Z_27 ));
    CascadeMux I__14390 (
            .O(N__66807),
            .I(N__66797));
    CascadeMux I__14389 (
            .O(N__66806),
            .I(N__66793));
    CascadeMux I__14388 (
            .O(N__66805),
            .I(N__66789));
    CascadeMux I__14387 (
            .O(N__66804),
            .I(N__66785));
    CascadeMux I__14386 (
            .O(N__66803),
            .I(N__66781));
    CascadeMux I__14385 (
            .O(N__66802),
            .I(N__66777));
    CascadeMux I__14384 (
            .O(N__66801),
            .I(N__66772));
    InMux I__14383 (
            .O(N__66800),
            .I(N__66760));
    InMux I__14382 (
            .O(N__66797),
            .I(N__66760));
    InMux I__14381 (
            .O(N__66796),
            .I(N__66760));
    InMux I__14380 (
            .O(N__66793),
            .I(N__66760));
    InMux I__14379 (
            .O(N__66792),
            .I(N__66760));
    InMux I__14378 (
            .O(N__66789),
            .I(N__66743));
    InMux I__14377 (
            .O(N__66788),
            .I(N__66743));
    InMux I__14376 (
            .O(N__66785),
            .I(N__66743));
    InMux I__14375 (
            .O(N__66784),
            .I(N__66743));
    InMux I__14374 (
            .O(N__66781),
            .I(N__66743));
    InMux I__14373 (
            .O(N__66780),
            .I(N__66743));
    InMux I__14372 (
            .O(N__66777),
            .I(N__66743));
    InMux I__14371 (
            .O(N__66776),
            .I(N__66743));
    InMux I__14370 (
            .O(N__66775),
            .I(N__66736));
    InMux I__14369 (
            .O(N__66772),
            .I(N__66736));
    InMux I__14368 (
            .O(N__66771),
            .I(N__66736));
    LocalMux I__14367 (
            .O(N__66760),
            .I(N__66729));
    LocalMux I__14366 (
            .O(N__66743),
            .I(N__66729));
    LocalMux I__14365 (
            .O(N__66736),
            .I(N__66729));
    Odrv12 I__14364 (
            .O(N__66729),
            .I(\pid_side.error_i_acummZ0Z_13 ));
    InMux I__14363 (
            .O(N__66726),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_27 ));
    InMux I__14362 (
            .O(N__66723),
            .I(N__66718));
    InMux I__14361 (
            .O(N__66722),
            .I(N__66715));
    InMux I__14360 (
            .O(N__66721),
            .I(N__66712));
    LocalMux I__14359 (
            .O(N__66718),
            .I(N__66709));
    LocalMux I__14358 (
            .O(N__66715),
            .I(N__66706));
    LocalMux I__14357 (
            .O(N__66712),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_27_c_RNI1NVS ));
    Odrv4 I__14356 (
            .O(N__66709),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_27_c_RNI1NVS ));
    Odrv12 I__14355 (
            .O(N__66706),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_27_c_RNI1NVS ));
    CascadeMux I__14354 (
            .O(N__66699),
            .I(N__66695));
    InMux I__14353 (
            .O(N__66698),
            .I(N__66690));
    InMux I__14352 (
            .O(N__66695),
            .I(N__66690));
    LocalMux I__14351 (
            .O(N__66690),
            .I(N__66687));
    Span12Mux_s10_v I__14350 (
            .O(N__66687),
            .I(N__66684));
    Odrv12 I__14349 (
            .O(N__66684),
            .I(\pid_side.error_i_acumm_preregZ0Z_25 ));
    InMux I__14348 (
            .O(N__66681),
            .I(N__66678));
    LocalMux I__14347 (
            .O(N__66678),
            .I(N__66675));
    Span4Mux_h I__14346 (
            .O(N__66675),
            .I(N__66672));
    Odrv4 I__14345 (
            .O(N__66672),
            .I(\pid_side.error_i_regZ0Z_14 ));
    InMux I__14344 (
            .O(N__66669),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_13 ));
    CascadeMux I__14343 (
            .O(N__66666),
            .I(N__66663));
    InMux I__14342 (
            .O(N__66663),
            .I(N__66660));
    LocalMux I__14341 (
            .O(N__66660),
            .I(N__66657));
    Span4Mux_h I__14340 (
            .O(N__66657),
            .I(N__66654));
    Odrv4 I__14339 (
            .O(N__66654),
            .I(\pid_side.error_i_regZ0Z_15 ));
    InMux I__14338 (
            .O(N__66651),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_14 ));
    CascadeMux I__14337 (
            .O(N__66648),
            .I(N__66645));
    InMux I__14336 (
            .O(N__66645),
            .I(N__66642));
    LocalMux I__14335 (
            .O(N__66642),
            .I(N__66639));
    Odrv4 I__14334 (
            .O(N__66639),
            .I(\pid_side.error_i_regZ0Z_16 ));
    InMux I__14333 (
            .O(N__66636),
            .I(bfn_16_15_0_));
    InMux I__14332 (
            .O(N__66633),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_16 ));
    CascadeMux I__14331 (
            .O(N__66630),
            .I(N__66627));
    InMux I__14330 (
            .O(N__66627),
            .I(N__66624));
    LocalMux I__14329 (
            .O(N__66624),
            .I(N__66621));
    Odrv12 I__14328 (
            .O(N__66621),
            .I(\pid_side.error_i_regZ0Z_18 ));
    InMux I__14327 (
            .O(N__66618),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_17 ));
    InMux I__14326 (
            .O(N__66615),
            .I(N__66612));
    LocalMux I__14325 (
            .O(N__66612),
            .I(N__66609));
    Span4Mux_h I__14324 (
            .O(N__66609),
            .I(N__66606));
    Odrv4 I__14323 (
            .O(N__66606),
            .I(\pid_side.error_i_regZ0Z_19 ));
    InMux I__14322 (
            .O(N__66603),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_18 ));
    CascadeMux I__14321 (
            .O(N__66600),
            .I(N__66597));
    InMux I__14320 (
            .O(N__66597),
            .I(N__66594));
    LocalMux I__14319 (
            .O(N__66594),
            .I(N__66591));
    Span4Mux_h I__14318 (
            .O(N__66591),
            .I(N__66588));
    Odrv4 I__14317 (
            .O(N__66588),
            .I(\pid_side.error_i_regZ0Z_20 ));
    InMux I__14316 (
            .O(N__66585),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_19 ));
    InMux I__14315 (
            .O(N__66582),
            .I(N__66579));
    LocalMux I__14314 (
            .O(N__66579),
            .I(N__66576));
    Span4Mux_h I__14313 (
            .O(N__66576),
            .I(N__66573));
    Odrv4 I__14312 (
            .O(N__66573),
            .I(\pid_side.error_i_regZ0Z_21 ));
    InMux I__14311 (
            .O(N__66570),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_20 ));
    CascadeMux I__14310 (
            .O(N__66567),
            .I(N__66564));
    InMux I__14309 (
            .O(N__66564),
            .I(N__66561));
    LocalMux I__14308 (
            .O(N__66561),
            .I(N__66558));
    Span4Mux_h I__14307 (
            .O(N__66558),
            .I(N__66555));
    Odrv4 I__14306 (
            .O(N__66555),
            .I(\pid_side.error_i_regZ0Z_22 ));
    InMux I__14305 (
            .O(N__66552),
            .I(N__66549));
    LocalMux I__14304 (
            .O(N__66549),
            .I(N__66546));
    Odrv4 I__14303 (
            .O(N__66546),
            .I(\pid_side.error_i_acummZ0Z_6 ));
    CascadeMux I__14302 (
            .O(N__66543),
            .I(N__66540));
    InMux I__14301 (
            .O(N__66540),
            .I(N__66537));
    LocalMux I__14300 (
            .O(N__66537),
            .I(N__66534));
    Odrv4 I__14299 (
            .O(N__66534),
            .I(\pid_side.error_i_regZ0Z_6 ));
    InMux I__14298 (
            .O(N__66531),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_5 ));
    InMux I__14297 (
            .O(N__66528),
            .I(N__66525));
    LocalMux I__14296 (
            .O(N__66525),
            .I(\pid_side.error_i_acummZ0Z_7 ));
    CascadeMux I__14295 (
            .O(N__66522),
            .I(N__66519));
    InMux I__14294 (
            .O(N__66519),
            .I(N__66516));
    LocalMux I__14293 (
            .O(N__66516),
            .I(N__66513));
    Span4Mux_v I__14292 (
            .O(N__66513),
            .I(N__66510));
    Odrv4 I__14291 (
            .O(N__66510),
            .I(\pid_side.error_i_regZ0Z_7 ));
    InMux I__14290 (
            .O(N__66507),
            .I(N__66502));
    InMux I__14289 (
            .O(N__66506),
            .I(N__66497));
    InMux I__14288 (
            .O(N__66505),
            .I(N__66497));
    LocalMux I__14287 (
            .O(N__66502),
            .I(N__66494));
    LocalMux I__14286 (
            .O(N__66497),
            .I(N__66491));
    Span4Mux_h I__14285 (
            .O(N__66494),
            .I(N__66488));
    Span4Mux_h I__14284 (
            .O(N__66491),
            .I(N__66485));
    Odrv4 I__14283 (
            .O(N__66488),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_6_c_RNIF9RN ));
    Odrv4 I__14282 (
            .O(N__66485),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_6_c_RNIF9RN ));
    InMux I__14281 (
            .O(N__66480),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_6 ));
    InMux I__14280 (
            .O(N__66477),
            .I(N__66474));
    LocalMux I__14279 (
            .O(N__66474),
            .I(N__66471));
    Odrv4 I__14278 (
            .O(N__66471),
            .I(\pid_side.error_i_acummZ0Z_8 ));
    InMux I__14277 (
            .O(N__66468),
            .I(N__66463));
    InMux I__14276 (
            .O(N__66467),
            .I(N__66460));
    InMux I__14275 (
            .O(N__66466),
            .I(N__66457));
    LocalMux I__14274 (
            .O(N__66463),
            .I(N__66454));
    LocalMux I__14273 (
            .O(N__66460),
            .I(N__66449));
    LocalMux I__14272 (
            .O(N__66457),
            .I(N__66449));
    Span4Mux_h I__14271 (
            .O(N__66454),
            .I(N__66446));
    Span4Mux_h I__14270 (
            .O(N__66449),
            .I(N__66443));
    Odrv4 I__14269 (
            .O(N__66446),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_7_c_RNI9JMJ ));
    Odrv4 I__14268 (
            .O(N__66443),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_7_c_RNI9JMJ ));
    InMux I__14267 (
            .O(N__66438),
            .I(bfn_16_14_0_));
    InMux I__14266 (
            .O(N__66435),
            .I(N__66432));
    LocalMux I__14265 (
            .O(N__66432),
            .I(N__66429));
    Odrv4 I__14264 (
            .O(N__66429),
            .I(\pid_side.error_i_acummZ0Z_9 ));
    InMux I__14263 (
            .O(N__66426),
            .I(N__66419));
    InMux I__14262 (
            .O(N__66425),
            .I(N__66419));
    InMux I__14261 (
            .O(N__66424),
            .I(N__66416));
    LocalMux I__14260 (
            .O(N__66419),
            .I(N__66413));
    LocalMux I__14259 (
            .O(N__66416),
            .I(N__66410));
    Span4Mux_h I__14258 (
            .O(N__66413),
            .I(N__66407));
    Odrv12 I__14257 (
            .O(N__66410),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_8_c_RNILHTN ));
    Odrv4 I__14256 (
            .O(N__66407),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_8_c_RNILHTN ));
    InMux I__14255 (
            .O(N__66402),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_8 ));
    InMux I__14254 (
            .O(N__66399),
            .I(N__66396));
    LocalMux I__14253 (
            .O(N__66396),
            .I(N__66393));
    Span4Mux_v I__14252 (
            .O(N__66393),
            .I(N__66390));
    Odrv4 I__14251 (
            .O(N__66390),
            .I(\pid_side.error_i_acummZ0Z_10 ));
    CascadeMux I__14250 (
            .O(N__66387),
            .I(N__66384));
    InMux I__14249 (
            .O(N__66384),
            .I(N__66381));
    LocalMux I__14248 (
            .O(N__66381),
            .I(N__66378));
    Odrv4 I__14247 (
            .O(N__66378),
            .I(\pid_side.error_i_regZ0Z_10 ));
    InMux I__14246 (
            .O(N__66375),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_9 ));
    InMux I__14245 (
            .O(N__66372),
            .I(N__66369));
    LocalMux I__14244 (
            .O(N__66369),
            .I(N__66366));
    Odrv4 I__14243 (
            .O(N__66366),
            .I(\pid_side.error_i_acummZ0Z_11 ));
    CascadeMux I__14242 (
            .O(N__66363),
            .I(N__66360));
    InMux I__14241 (
            .O(N__66360),
            .I(N__66357));
    LocalMux I__14240 (
            .O(N__66357),
            .I(N__66354));
    Span4Mux_h I__14239 (
            .O(N__66354),
            .I(N__66351));
    Odrv4 I__14238 (
            .O(N__66351),
            .I(\pid_side.error_i_regZ0Z_11 ));
    InMux I__14237 (
            .O(N__66348),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_10 ));
    InMux I__14236 (
            .O(N__66345),
            .I(N__66342));
    LocalMux I__14235 (
            .O(N__66342),
            .I(N__66339));
    Span4Mux_h I__14234 (
            .O(N__66339),
            .I(N__66336));
    Odrv4 I__14233 (
            .O(N__66336),
            .I(\pid_side.error_i_acummZ0Z_12 ));
    InMux I__14232 (
            .O(N__66333),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_11 ));
    InMux I__14231 (
            .O(N__66330),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_12 ));
    InMux I__14230 (
            .O(N__66327),
            .I(N__66324));
    LocalMux I__14229 (
            .O(N__66324),
            .I(N__66320));
    InMux I__14228 (
            .O(N__66323),
            .I(N__66317));
    Odrv4 I__14227 (
            .O(N__66320),
            .I(\pid_side.un1_pid_prereg_0_24 ));
    LocalMux I__14226 (
            .O(N__66317),
            .I(\pid_side.un1_pid_prereg_0_24 ));
    CascadeMux I__14225 (
            .O(N__66312),
            .I(N__66308));
    CascadeMux I__14224 (
            .O(N__66311),
            .I(N__66304));
    InMux I__14223 (
            .O(N__66308),
            .I(N__66299));
    InMux I__14222 (
            .O(N__66307),
            .I(N__66299));
    InMux I__14221 (
            .O(N__66304),
            .I(N__66296));
    LocalMux I__14220 (
            .O(N__66299),
            .I(\pid_side.un1_pid_prereg_0_26 ));
    LocalMux I__14219 (
            .O(N__66296),
            .I(\pid_side.un1_pid_prereg_0_26 ));
    InMux I__14218 (
            .O(N__66291),
            .I(N__66281));
    InMux I__14217 (
            .O(N__66290),
            .I(N__66281));
    InMux I__14216 (
            .O(N__66289),
            .I(N__66276));
    InMux I__14215 (
            .O(N__66288),
            .I(N__66276));
    InMux I__14214 (
            .O(N__66287),
            .I(N__66271));
    InMux I__14213 (
            .O(N__66286),
            .I(N__66271));
    LocalMux I__14212 (
            .O(N__66281),
            .I(N__66266));
    LocalMux I__14211 (
            .O(N__66276),
            .I(N__66266));
    LocalMux I__14210 (
            .O(N__66271),
            .I(\pid_side.un1_pid_prereg_0_25 ));
    Odrv4 I__14209 (
            .O(N__66266),
            .I(\pid_side.un1_pid_prereg_0_25 ));
    InMux I__14208 (
            .O(N__66261),
            .I(N__66258));
    LocalMux I__14207 (
            .O(N__66258),
            .I(N__66255));
    Span12Mux_v I__14206 (
            .O(N__66255),
            .I(N__66251));
    InMux I__14205 (
            .O(N__66254),
            .I(N__66248));
    Odrv12 I__14204 (
            .O(N__66251),
            .I(\pid_side.error_i_acummZ0Z_0 ));
    LocalMux I__14203 (
            .O(N__66248),
            .I(\pid_side.error_i_acummZ0Z_0 ));
    InMux I__14202 (
            .O(N__66243),
            .I(N__66240));
    LocalMux I__14201 (
            .O(N__66240),
            .I(N__66236));
    CascadeMux I__14200 (
            .O(N__66239),
            .I(N__66233));
    Span12Mux_v I__14199 (
            .O(N__66236),
            .I(N__66230));
    InMux I__14198 (
            .O(N__66233),
            .I(N__66227));
    Odrv12 I__14197 (
            .O(N__66230),
            .I(\pid_side.error_i_regZ0Z_0 ));
    LocalMux I__14196 (
            .O(N__66227),
            .I(\pid_side.error_i_regZ0Z_0 ));
    InMux I__14195 (
            .O(N__66222),
            .I(N__66219));
    LocalMux I__14194 (
            .O(N__66219),
            .I(N__66216));
    Odrv4 I__14193 (
            .O(N__66216),
            .I(\pid_side.error_i_acummZ0Z_1 ));
    CascadeMux I__14192 (
            .O(N__66213),
            .I(N__66210));
    InMux I__14191 (
            .O(N__66210),
            .I(N__66207));
    LocalMux I__14190 (
            .O(N__66207),
            .I(N__66204));
    Odrv4 I__14189 (
            .O(N__66204),
            .I(\pid_side.error_i_regZ0Z_1 ));
    InMux I__14188 (
            .O(N__66201),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_0 ));
    InMux I__14187 (
            .O(N__66198),
            .I(N__66195));
    LocalMux I__14186 (
            .O(N__66195),
            .I(N__66192));
    Odrv4 I__14185 (
            .O(N__66192),
            .I(\pid_side.error_i_acummZ0Z_2 ));
    CascadeMux I__14184 (
            .O(N__66189),
            .I(N__66186));
    InMux I__14183 (
            .O(N__66186),
            .I(N__66183));
    LocalMux I__14182 (
            .O(N__66183),
            .I(\pid_side.error_i_regZ0Z_2 ));
    InMux I__14181 (
            .O(N__66180),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_1 ));
    InMux I__14180 (
            .O(N__66177),
            .I(N__66174));
    LocalMux I__14179 (
            .O(N__66174),
            .I(N__66171));
    Odrv4 I__14178 (
            .O(N__66171),
            .I(\pid_side.error_i_acummZ0Z_3 ));
    CascadeMux I__14177 (
            .O(N__66168),
            .I(N__66165));
    InMux I__14176 (
            .O(N__66165),
            .I(N__66162));
    LocalMux I__14175 (
            .O(N__66162),
            .I(N__66159));
    Odrv4 I__14174 (
            .O(N__66159),
            .I(\pid_side.error_i_regZ0Z_3 ));
    InMux I__14173 (
            .O(N__66156),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_2 ));
    InMux I__14172 (
            .O(N__66153),
            .I(N__66150));
    LocalMux I__14171 (
            .O(N__66150),
            .I(N__66147));
    Odrv4 I__14170 (
            .O(N__66147),
            .I(\pid_side.error_i_acummZ0Z_4 ));
    InMux I__14169 (
            .O(N__66144),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_3 ));
    InMux I__14168 (
            .O(N__66141),
            .I(N__66138));
    LocalMux I__14167 (
            .O(N__66138),
            .I(N__66135));
    Odrv4 I__14166 (
            .O(N__66135),
            .I(\pid_side.error_i_acummZ0Z_5 ));
    InMux I__14165 (
            .O(N__66132),
            .I(\pid_side.un1_error_i_acumm_prereg_cry_4 ));
    CascadeMux I__14164 (
            .O(N__66129),
            .I(N__66126));
    InMux I__14163 (
            .O(N__66126),
            .I(N__66119));
    InMux I__14162 (
            .O(N__66125),
            .I(N__66119));
    InMux I__14161 (
            .O(N__66124),
            .I(N__66116));
    LocalMux I__14160 (
            .O(N__66119),
            .I(N__66113));
    LocalMux I__14159 (
            .O(N__66116),
            .I(\pid_side.error_i_acumm_preregZ0Z_6 ));
    Odrv4 I__14158 (
            .O(N__66113),
            .I(\pid_side.error_i_acumm_preregZ0Z_6 ));
    CEMux I__14157 (
            .O(N__66108),
            .I(N__66104));
    CEMux I__14156 (
            .O(N__66107),
            .I(N__66101));
    LocalMux I__14155 (
            .O(N__66104),
            .I(N__66097));
    LocalMux I__14154 (
            .O(N__66101),
            .I(N__66094));
    CEMux I__14153 (
            .O(N__66100),
            .I(N__66090));
    Span4Mux_v I__14152 (
            .O(N__66097),
            .I(N__66085));
    Span4Mux_v I__14151 (
            .O(N__66094),
            .I(N__66085));
    CEMux I__14150 (
            .O(N__66093),
            .I(N__66082));
    LocalMux I__14149 (
            .O(N__66090),
            .I(N__66079));
    Span4Mux_h I__14148 (
            .O(N__66085),
            .I(N__66074));
    LocalMux I__14147 (
            .O(N__66082),
            .I(N__66074));
    Span4Mux_h I__14146 (
            .O(N__66079),
            .I(N__66071));
    Span4Mux_h I__14145 (
            .O(N__66074),
            .I(N__66068));
    Odrv4 I__14144 (
            .O(N__66071),
            .I(\pid_side.error_i_acumm_1_sqmuxa_1_i ));
    Odrv4 I__14143 (
            .O(N__66068),
            .I(\pid_side.error_i_acumm_1_sqmuxa_1_i ));
    InMux I__14142 (
            .O(N__66063),
            .I(N__66060));
    LocalMux I__14141 (
            .O(N__66060),
            .I(N__66057));
    Odrv12 I__14140 (
            .O(N__66057),
            .I(\pid_side.error_i_acumm16lto27_13 ));
    InMux I__14139 (
            .O(N__66054),
            .I(N__66051));
    LocalMux I__14138 (
            .O(N__66051),
            .I(N__66048));
    Odrv4 I__14137 (
            .O(N__66048),
            .I(\pid_side.error_i_acumm_prereg_esr_RNIBT1C4Z0Z_12 ));
    InMux I__14136 (
            .O(N__66045),
            .I(N__66040));
    CascadeMux I__14135 (
            .O(N__66044),
            .I(N__66034));
    InMux I__14134 (
            .O(N__66043),
            .I(N__66031));
    LocalMux I__14133 (
            .O(N__66040),
            .I(N__66028));
    InMux I__14132 (
            .O(N__66039),
            .I(N__66025));
    InMux I__14131 (
            .O(N__66038),
            .I(N__66022));
    InMux I__14130 (
            .O(N__66037),
            .I(N__66019));
    InMux I__14129 (
            .O(N__66034),
            .I(N__66016));
    LocalMux I__14128 (
            .O(N__66031),
            .I(N__66013));
    Span4Mux_v I__14127 (
            .O(N__66028),
            .I(N__66008));
    LocalMux I__14126 (
            .O(N__66025),
            .I(N__66008));
    LocalMux I__14125 (
            .O(N__66022),
            .I(N__66005));
    LocalMux I__14124 (
            .O(N__66019),
            .I(N__66001));
    LocalMux I__14123 (
            .O(N__66016),
            .I(N__65998));
    Span4Mux_v I__14122 (
            .O(N__66013),
            .I(N__65995));
    Span4Mux_h I__14121 (
            .O(N__66008),
            .I(N__65991));
    Span4Mux_v I__14120 (
            .O(N__66005),
            .I(N__65988));
    InMux I__14119 (
            .O(N__66004),
            .I(N__65984));
    Span4Mux_h I__14118 (
            .O(N__66001),
            .I(N__65979));
    Span4Mux_v I__14117 (
            .O(N__65998),
            .I(N__65979));
    Span4Mux_h I__14116 (
            .O(N__65995),
            .I(N__65976));
    InMux I__14115 (
            .O(N__65994),
            .I(N__65973));
    Sp12to4 I__14114 (
            .O(N__65991),
            .I(N__65970));
    Sp12to4 I__14113 (
            .O(N__65988),
            .I(N__65967));
    InMux I__14112 (
            .O(N__65987),
            .I(N__65964));
    LocalMux I__14111 (
            .O(N__65984),
            .I(N__65961));
    Span4Mux_v I__14110 (
            .O(N__65979),
            .I(N__65958));
    Sp12to4 I__14109 (
            .O(N__65976),
            .I(N__65951));
    LocalMux I__14108 (
            .O(N__65973),
            .I(N__65951));
    Span12Mux_v I__14107 (
            .O(N__65970),
            .I(N__65951));
    Span12Mux_h I__14106 (
            .O(N__65967),
            .I(N__65944));
    LocalMux I__14105 (
            .O(N__65964),
            .I(N__65944));
    Span12Mux_v I__14104 (
            .O(N__65961),
            .I(N__65944));
    Sp12to4 I__14103 (
            .O(N__65958),
            .I(N__65936));
    Span12Mux_v I__14102 (
            .O(N__65951),
            .I(N__65936));
    Span12Mux_v I__14101 (
            .O(N__65944),
            .I(N__65936));
    IoInMux I__14100 (
            .O(N__65943),
            .I(N__65933));
    Odrv12 I__14099 (
            .O(N__65936),
            .I(reset_system));
    LocalMux I__14098 (
            .O(N__65933),
            .I(reset_system));
    InMux I__14097 (
            .O(N__65928),
            .I(N__65920));
    InMux I__14096 (
            .O(N__65927),
            .I(N__65909));
    InMux I__14095 (
            .O(N__65926),
            .I(N__65909));
    InMux I__14094 (
            .O(N__65925),
            .I(N__65909));
    InMux I__14093 (
            .O(N__65924),
            .I(N__65909));
    InMux I__14092 (
            .O(N__65923),
            .I(N__65909));
    LocalMux I__14091 (
            .O(N__65920),
            .I(\pid_side.error_i_acumm_2_sqmuxa_1 ));
    LocalMux I__14090 (
            .O(N__65909),
            .I(\pid_side.error_i_acumm_2_sqmuxa_1 ));
    CascadeMux I__14089 (
            .O(N__65904),
            .I(\pid_side.error_i_acumm_2_sqmuxa_1_cascade_ ));
    InMux I__14088 (
            .O(N__65901),
            .I(N__65898));
    LocalMux I__14087 (
            .O(N__65898),
            .I(\pid_side.error_i_acumm_prereg_esr_RNIGIQP9Z0Z_12 ));
    CascadeMux I__14086 (
            .O(N__65895),
            .I(N__65886));
    InMux I__14085 (
            .O(N__65894),
            .I(N__65876));
    InMux I__14084 (
            .O(N__65893),
            .I(N__65865));
    InMux I__14083 (
            .O(N__65892),
            .I(N__65865));
    InMux I__14082 (
            .O(N__65891),
            .I(N__65865));
    InMux I__14081 (
            .O(N__65890),
            .I(N__65865));
    InMux I__14080 (
            .O(N__65889),
            .I(N__65865));
    InMux I__14079 (
            .O(N__65886),
            .I(N__65858));
    InMux I__14078 (
            .O(N__65885),
            .I(N__65858));
    InMux I__14077 (
            .O(N__65884),
            .I(N__65858));
    InMux I__14076 (
            .O(N__65883),
            .I(N__65847));
    InMux I__14075 (
            .O(N__65882),
            .I(N__65847));
    InMux I__14074 (
            .O(N__65881),
            .I(N__65847));
    InMux I__14073 (
            .O(N__65880),
            .I(N__65847));
    InMux I__14072 (
            .O(N__65879),
            .I(N__65847));
    LocalMux I__14071 (
            .O(N__65876),
            .I(\pid_side.error_i_acumm_2_sqmuxa ));
    LocalMux I__14070 (
            .O(N__65865),
            .I(\pid_side.error_i_acumm_2_sqmuxa ));
    LocalMux I__14069 (
            .O(N__65858),
            .I(\pid_side.error_i_acumm_2_sqmuxa ));
    LocalMux I__14068 (
            .O(N__65847),
            .I(\pid_side.error_i_acumm_2_sqmuxa ));
    CascadeMux I__14067 (
            .O(N__65838),
            .I(\pid_side.un1_pid_prereg_370_1_cascade_ ));
    CascadeMux I__14066 (
            .O(N__65835),
            .I(\pid_side.un1_pid_prereg_0_14_cascade_ ));
    CascadeMux I__14065 (
            .O(N__65832),
            .I(\pid_side.un1_pid_prereg_0_15_cascade_ ));
    InMux I__14064 (
            .O(N__65829),
            .I(N__65823));
    InMux I__14063 (
            .O(N__65828),
            .I(N__65823));
    LocalMux I__14062 (
            .O(N__65823),
            .I(\pid_side.error_i_acumm16lto3 ));
    InMux I__14061 (
            .O(N__65820),
            .I(N__65816));
    InMux I__14060 (
            .O(N__65819),
            .I(N__65813));
    LocalMux I__14059 (
            .O(N__65816),
            .I(N__65810));
    LocalMux I__14058 (
            .O(N__65813),
            .I(\pid_side.error_i_acumm_preregZ0Z_16 ));
    Odrv4 I__14057 (
            .O(N__65810),
            .I(\pid_side.error_i_acumm_preregZ0Z_16 ));
    CascadeMux I__14056 (
            .O(N__65805),
            .I(N__65801));
    InMux I__14055 (
            .O(N__65804),
            .I(N__65798));
    InMux I__14054 (
            .O(N__65801),
            .I(N__65795));
    LocalMux I__14053 (
            .O(N__65798),
            .I(N__65791));
    LocalMux I__14052 (
            .O(N__65795),
            .I(N__65788));
    InMux I__14051 (
            .O(N__65794),
            .I(N__65785));
    Span4Mux_h I__14050 (
            .O(N__65791),
            .I(N__65782));
    Odrv4 I__14049 (
            .O(N__65788),
            .I(\pid_side.error_i_acumm_preregZ0Z_9 ));
    LocalMux I__14048 (
            .O(N__65785),
            .I(\pid_side.error_i_acumm_preregZ0Z_9 ));
    Odrv4 I__14047 (
            .O(N__65782),
            .I(\pid_side.error_i_acumm_preregZ0Z_9 ));
    InMux I__14046 (
            .O(N__65775),
            .I(N__65769));
    InMux I__14045 (
            .O(N__65774),
            .I(N__65769));
    LocalMux I__14044 (
            .O(N__65769),
            .I(\pid_side.error_i_acumm_preregZ0Z_27 ));
    CascadeMux I__14043 (
            .O(N__65766),
            .I(N__65763));
    InMux I__14042 (
            .O(N__65763),
            .I(N__65760));
    LocalMux I__14041 (
            .O(N__65760),
            .I(N__65755));
    InMux I__14040 (
            .O(N__65759),
            .I(N__65750));
    InMux I__14039 (
            .O(N__65758),
            .I(N__65750));
    Odrv12 I__14038 (
            .O(N__65755),
            .I(\pid_side.error_i_acumm_preregZ0Z_11 ));
    LocalMux I__14037 (
            .O(N__65750),
            .I(\pid_side.error_i_acumm_preregZ0Z_11 ));
    InMux I__14036 (
            .O(N__65745),
            .I(N__65740));
    InMux I__14035 (
            .O(N__65744),
            .I(N__65735));
    InMux I__14034 (
            .O(N__65743),
            .I(N__65735));
    LocalMux I__14033 (
            .O(N__65740),
            .I(\pid_side.error_i_acumm_preregZ0Z_4 ));
    LocalMux I__14032 (
            .O(N__65735),
            .I(\pid_side.error_i_acumm_preregZ0Z_4 ));
    InMux I__14031 (
            .O(N__65730),
            .I(N__65727));
    LocalMux I__14030 (
            .O(N__65727),
            .I(\pid_side.error_i_acumm16lto27_9 ));
    CascadeMux I__14029 (
            .O(N__65724),
            .I(\pid_side.error_i_acumm16lto27_8_cascade_ ));
    InMux I__14028 (
            .O(N__65721),
            .I(N__65718));
    LocalMux I__14027 (
            .O(N__65718),
            .I(\pid_side.error_i_acumm16lto27_7 ));
    InMux I__14026 (
            .O(N__65715),
            .I(N__65711));
    InMux I__14025 (
            .O(N__65714),
            .I(N__65708));
    LocalMux I__14024 (
            .O(N__65711),
            .I(\pid_side.error_i_acumm_preregZ0Z_15 ));
    LocalMux I__14023 (
            .O(N__65708),
            .I(\pid_side.error_i_acumm_preregZ0Z_15 ));
    InMux I__14022 (
            .O(N__65703),
            .I(N__65699));
    InMux I__14021 (
            .O(N__65702),
            .I(N__65696));
    LocalMux I__14020 (
            .O(N__65699),
            .I(\pid_side.error_i_acumm_preregZ0Z_14 ));
    LocalMux I__14019 (
            .O(N__65696),
            .I(\pid_side.error_i_acumm_preregZ0Z_14 ));
    InMux I__14018 (
            .O(N__65691),
            .I(N__65688));
    LocalMux I__14017 (
            .O(N__65688),
            .I(\pid_side.error_i_acumm16lto27_10 ));
    CascadeMux I__14016 (
            .O(N__65685),
            .I(\pid_side.un10lto27_8_cascade_ ));
    InMux I__14015 (
            .O(N__65682),
            .I(N__65679));
    LocalMux I__14014 (
            .O(N__65679),
            .I(\pid_side.un10lto27_11 ));
    CascadeMux I__14013 (
            .O(N__65676),
            .I(N__65673));
    InMux I__14012 (
            .O(N__65673),
            .I(N__65667));
    InMux I__14011 (
            .O(N__65672),
            .I(N__65667));
    LocalMux I__14010 (
            .O(N__65667),
            .I(\pid_side.error_i_acumm_preregZ0Z_26 ));
    InMux I__14009 (
            .O(N__65664),
            .I(N__65658));
    InMux I__14008 (
            .O(N__65663),
            .I(N__65658));
    LocalMux I__14007 (
            .O(N__65658),
            .I(\pid_side.error_i_acumm_preregZ0Z_1 ));
    CascadeMux I__14006 (
            .O(N__65655),
            .I(N__65651));
    InMux I__14005 (
            .O(N__65654),
            .I(N__65648));
    InMux I__14004 (
            .O(N__65651),
            .I(N__65645));
    LocalMux I__14003 (
            .O(N__65648),
            .I(\pid_side.error_i_acumm_preregZ0Z_2 ));
    LocalMux I__14002 (
            .O(N__65645),
            .I(\pid_side.error_i_acumm_preregZ0Z_2 ));
    CascadeMux I__14001 (
            .O(N__65640),
            .I(\pid_side.un10lto27_10_cascade_ ));
    InMux I__14000 (
            .O(N__65637),
            .I(N__65634));
    LocalMux I__13999 (
            .O(N__65634),
            .I(N__65631));
    Span4Mux_v I__13998 (
            .O(N__65631),
            .I(N__65628));
    Odrv4 I__13997 (
            .O(N__65628),
            .I(\pid_side.error_i_acumm_prereg_esr_RNI5LOD5_0Z0Z_14 ));
    InMux I__13996 (
            .O(N__65625),
            .I(N__65622));
    LocalMux I__13995 (
            .O(N__65622),
            .I(\pid_side.un10lto27_9 ));
    InMux I__13994 (
            .O(N__65619),
            .I(N__65615));
    InMux I__13993 (
            .O(N__65618),
            .I(N__65612));
    LocalMux I__13992 (
            .O(N__65615),
            .I(\pid_side.error_i_acumm_preregZ0Z_20 ));
    LocalMux I__13991 (
            .O(N__65612),
            .I(\pid_side.error_i_acumm_preregZ0Z_20 ));
    InMux I__13990 (
            .O(N__65607),
            .I(N__65603));
    InMux I__13989 (
            .O(N__65606),
            .I(N__65600));
    LocalMux I__13988 (
            .O(N__65603),
            .I(\pid_side.error_i_acumm_preregZ0Z_19 ));
    LocalMux I__13987 (
            .O(N__65600),
            .I(\pid_side.error_i_acumm_preregZ0Z_19 ));
    CascadeMux I__13986 (
            .O(N__65595),
            .I(N__65592));
    InMux I__13985 (
            .O(N__65592),
            .I(N__65588));
    InMux I__13984 (
            .O(N__65591),
            .I(N__65585));
    LocalMux I__13983 (
            .O(N__65588),
            .I(\pid_side.error_i_acumm_preregZ0Z_18 ));
    LocalMux I__13982 (
            .O(N__65585),
            .I(\pid_side.error_i_acumm_preregZ0Z_18 ));
    InMux I__13981 (
            .O(N__65580),
            .I(\ppm_encoder_1.un1_counter_13_cry_10 ));
    InMux I__13980 (
            .O(N__65577),
            .I(N__65572));
    InMux I__13979 (
            .O(N__65576),
            .I(N__65569));
    InMux I__13978 (
            .O(N__65575),
            .I(N__65566));
    LocalMux I__13977 (
            .O(N__65572),
            .I(N__65563));
    LocalMux I__13976 (
            .O(N__65569),
            .I(\ppm_encoder_1.counterZ0Z_12 ));
    LocalMux I__13975 (
            .O(N__65566),
            .I(\ppm_encoder_1.counterZ0Z_12 ));
    Odrv4 I__13974 (
            .O(N__65563),
            .I(\ppm_encoder_1.counterZ0Z_12 ));
    InMux I__13973 (
            .O(N__65556),
            .I(\ppm_encoder_1.un1_counter_13_cry_11 ));
    InMux I__13972 (
            .O(N__65553),
            .I(N__65548));
    InMux I__13971 (
            .O(N__65552),
            .I(N__65545));
    InMux I__13970 (
            .O(N__65551),
            .I(N__65542));
    LocalMux I__13969 (
            .O(N__65548),
            .I(N__65539));
    LocalMux I__13968 (
            .O(N__65545),
            .I(\ppm_encoder_1.counterZ0Z_13 ));
    LocalMux I__13967 (
            .O(N__65542),
            .I(\ppm_encoder_1.counterZ0Z_13 ));
    Odrv4 I__13966 (
            .O(N__65539),
            .I(\ppm_encoder_1.counterZ0Z_13 ));
    InMux I__13965 (
            .O(N__65532),
            .I(\ppm_encoder_1.un1_counter_13_cry_12 ));
    InMux I__13964 (
            .O(N__65529),
            .I(\ppm_encoder_1.un1_counter_13_cry_13 ));
    InMux I__13963 (
            .O(N__65526),
            .I(\ppm_encoder_1.un1_counter_13_cry_14 ));
    InMux I__13962 (
            .O(N__65523),
            .I(bfn_16_6_0_));
    InMux I__13961 (
            .O(N__65520),
            .I(\ppm_encoder_1.un1_counter_13_cry_16 ));
    InMux I__13960 (
            .O(N__65517),
            .I(\ppm_encoder_1.un1_counter_13_cry_17 ));
    InMux I__13959 (
            .O(N__65514),
            .I(N__65511));
    LocalMux I__13958 (
            .O(N__65511),
            .I(N__65505));
    InMux I__13957 (
            .O(N__65510),
            .I(N__65502));
    InMux I__13956 (
            .O(N__65509),
            .I(N__65497));
    InMux I__13955 (
            .O(N__65508),
            .I(N__65497));
    Span4Mux_h I__13954 (
            .O(N__65505),
            .I(N__65494));
    LocalMux I__13953 (
            .O(N__65502),
            .I(\ppm_encoder_1.counterZ0Z_18 ));
    LocalMux I__13952 (
            .O(N__65497),
            .I(\ppm_encoder_1.counterZ0Z_18 ));
    Odrv4 I__13951 (
            .O(N__65494),
            .I(\ppm_encoder_1.counterZ0Z_18 ));
    SRMux I__13950 (
            .O(N__65487),
            .I(N__65483));
    SRMux I__13949 (
            .O(N__65486),
            .I(N__65480));
    LocalMux I__13948 (
            .O(N__65483),
            .I(N__65476));
    LocalMux I__13947 (
            .O(N__65480),
            .I(N__65473));
    SRMux I__13946 (
            .O(N__65479),
            .I(N__65470));
    Span4Mux_h I__13945 (
            .O(N__65476),
            .I(N__65467));
    Span4Mux_s3_v I__13944 (
            .O(N__65473),
            .I(N__65462));
    LocalMux I__13943 (
            .O(N__65470),
            .I(N__65462));
    Odrv4 I__13942 (
            .O(N__65467),
            .I(\ppm_encoder_1.counter24_0_I_57_c_RNIGCOZ0Z83 ));
    Odrv4 I__13941 (
            .O(N__65462),
            .I(\ppm_encoder_1.counter24_0_I_57_c_RNIGCOZ0Z83 ));
    InMux I__13940 (
            .O(N__65457),
            .I(N__65451));
    CascadeMux I__13939 (
            .O(N__65456),
            .I(N__65446));
    CascadeMux I__13938 (
            .O(N__65455),
            .I(N__65443));
    CascadeMux I__13937 (
            .O(N__65454),
            .I(N__65440));
    LocalMux I__13936 (
            .O(N__65451),
            .I(N__65433));
    InMux I__13935 (
            .O(N__65450),
            .I(N__65415));
    InMux I__13934 (
            .O(N__65449),
            .I(N__65415));
    InMux I__13933 (
            .O(N__65446),
            .I(N__65415));
    InMux I__13932 (
            .O(N__65443),
            .I(N__65415));
    InMux I__13931 (
            .O(N__65440),
            .I(N__65415));
    InMux I__13930 (
            .O(N__65439),
            .I(N__65415));
    InMux I__13929 (
            .O(N__65438),
            .I(N__65415));
    InMux I__13928 (
            .O(N__65437),
            .I(N__65415));
    InMux I__13927 (
            .O(N__65436),
            .I(N__65412));
    Span4Mux_v I__13926 (
            .O(N__65433),
            .I(N__65409));
    CascadeMux I__13925 (
            .O(N__65432),
            .I(N__65404));
    LocalMux I__13924 (
            .O(N__65415),
            .I(N__65393));
    LocalMux I__13923 (
            .O(N__65412),
            .I(N__65390));
    Span4Mux_v I__13922 (
            .O(N__65409),
            .I(N__65387));
    InMux I__13921 (
            .O(N__65408),
            .I(N__65372));
    InMux I__13920 (
            .O(N__65407),
            .I(N__65372));
    InMux I__13919 (
            .O(N__65404),
            .I(N__65372));
    InMux I__13918 (
            .O(N__65403),
            .I(N__65372));
    InMux I__13917 (
            .O(N__65402),
            .I(N__65372));
    InMux I__13916 (
            .O(N__65401),
            .I(N__65372));
    InMux I__13915 (
            .O(N__65400),
            .I(N__65372));
    InMux I__13914 (
            .O(N__65399),
            .I(N__65365));
    InMux I__13913 (
            .O(N__65398),
            .I(N__65365));
    InMux I__13912 (
            .O(N__65397),
            .I(N__65365));
    InMux I__13911 (
            .O(N__65396),
            .I(N__65362));
    Span4Mux_h I__13910 (
            .O(N__65393),
            .I(N__65359));
    Span4Mux_v I__13909 (
            .O(N__65390),
            .I(N__65356));
    Span4Mux_v I__13908 (
            .O(N__65387),
            .I(N__65351));
    LocalMux I__13907 (
            .O(N__65372),
            .I(N__65351));
    LocalMux I__13906 (
            .O(N__65365),
            .I(N__65348));
    LocalMux I__13905 (
            .O(N__65362),
            .I(N__65344));
    Sp12to4 I__13904 (
            .O(N__65359),
            .I(N__65341));
    Span4Mux_h I__13903 (
            .O(N__65356),
            .I(N__65333));
    Span4Mux_h I__13902 (
            .O(N__65351),
            .I(N__65333));
    Span4Mux_h I__13901 (
            .O(N__65348),
            .I(N__65333));
    InMux I__13900 (
            .O(N__65347),
            .I(N__65330));
    Span4Mux_v I__13899 (
            .O(N__65344),
            .I(N__65327));
    Span12Mux_v I__13898 (
            .O(N__65341),
            .I(N__65324));
    InMux I__13897 (
            .O(N__65340),
            .I(N__65321));
    Span4Mux_h I__13896 (
            .O(N__65333),
            .I(N__65318));
    LocalMux I__13895 (
            .O(N__65330),
            .I(\pid_alt.N_72_i ));
    Odrv4 I__13894 (
            .O(N__65327),
            .I(\pid_alt.N_72_i ));
    Odrv12 I__13893 (
            .O(N__65324),
            .I(\pid_alt.N_72_i ));
    LocalMux I__13892 (
            .O(N__65321),
            .I(\pid_alt.N_72_i ));
    Odrv4 I__13891 (
            .O(N__65318),
            .I(\pid_alt.N_72_i ));
    CascadeMux I__13890 (
            .O(N__65307),
            .I(N__65300));
    CascadeMux I__13889 (
            .O(N__65306),
            .I(N__65292));
    CascadeMux I__13888 (
            .O(N__65305),
            .I(N__65280));
    CascadeMux I__13887 (
            .O(N__65304),
            .I(N__65274));
    CascadeMux I__13886 (
            .O(N__65303),
            .I(N__65268));
    InMux I__13885 (
            .O(N__65300),
            .I(N__65261));
    CascadeMux I__13884 (
            .O(N__65299),
            .I(N__65258));
    CascadeMux I__13883 (
            .O(N__65298),
            .I(N__65255));
    CascadeMux I__13882 (
            .O(N__65297),
            .I(N__65252));
    CascadeMux I__13881 (
            .O(N__65296),
            .I(N__65249));
    CascadeMux I__13880 (
            .O(N__65295),
            .I(N__65244));
    InMux I__13879 (
            .O(N__65292),
            .I(N__65240));
    CascadeMux I__13878 (
            .O(N__65291),
            .I(N__65237));
    CascadeMux I__13877 (
            .O(N__65290),
            .I(N__65234));
    CascadeMux I__13876 (
            .O(N__65289),
            .I(N__65231));
    CascadeMux I__13875 (
            .O(N__65288),
            .I(N__65228));
    CascadeMux I__13874 (
            .O(N__65287),
            .I(N__65225));
    CascadeMux I__13873 (
            .O(N__65286),
            .I(N__65219));
    CascadeMux I__13872 (
            .O(N__65285),
            .I(N__65214));
    CascadeMux I__13871 (
            .O(N__65284),
            .I(N__65210));
    InMux I__13870 (
            .O(N__65283),
            .I(N__65197));
    InMux I__13869 (
            .O(N__65280),
            .I(N__65197));
    InMux I__13868 (
            .O(N__65279),
            .I(N__65197));
    InMux I__13867 (
            .O(N__65278),
            .I(N__65197));
    InMux I__13866 (
            .O(N__65277),
            .I(N__65197));
    InMux I__13865 (
            .O(N__65274),
            .I(N__65197));
    CascadeMux I__13864 (
            .O(N__65273),
            .I(N__65194));
    CascadeMux I__13863 (
            .O(N__65272),
            .I(N__65191));
    CascadeMux I__13862 (
            .O(N__65271),
            .I(N__65184));
    InMux I__13861 (
            .O(N__65268),
            .I(N__65177));
    InMux I__13860 (
            .O(N__65267),
            .I(N__65177));
    CascadeMux I__13859 (
            .O(N__65266),
            .I(N__65174));
    CascadeMux I__13858 (
            .O(N__65265),
            .I(N__65169));
    CascadeMux I__13857 (
            .O(N__65264),
            .I(N__65164));
    LocalMux I__13856 (
            .O(N__65261),
            .I(N__65161));
    InMux I__13855 (
            .O(N__65258),
            .I(N__65156));
    InMux I__13854 (
            .O(N__65255),
            .I(N__65156));
    InMux I__13853 (
            .O(N__65252),
            .I(N__65149));
    InMux I__13852 (
            .O(N__65249),
            .I(N__65149));
    InMux I__13851 (
            .O(N__65248),
            .I(N__65149));
    InMux I__13850 (
            .O(N__65247),
            .I(N__65142));
    InMux I__13849 (
            .O(N__65244),
            .I(N__65142));
    InMux I__13848 (
            .O(N__65243),
            .I(N__65142));
    LocalMux I__13847 (
            .O(N__65240),
            .I(N__65139));
    InMux I__13846 (
            .O(N__65237),
            .I(N__65134));
    InMux I__13845 (
            .O(N__65234),
            .I(N__65134));
    InMux I__13844 (
            .O(N__65231),
            .I(N__65121));
    InMux I__13843 (
            .O(N__65228),
            .I(N__65121));
    InMux I__13842 (
            .O(N__65225),
            .I(N__65121));
    InMux I__13841 (
            .O(N__65224),
            .I(N__65121));
    InMux I__13840 (
            .O(N__65223),
            .I(N__65121));
    InMux I__13839 (
            .O(N__65222),
            .I(N__65121));
    InMux I__13838 (
            .O(N__65219),
            .I(N__65108));
    InMux I__13837 (
            .O(N__65218),
            .I(N__65108));
    InMux I__13836 (
            .O(N__65217),
            .I(N__65108));
    InMux I__13835 (
            .O(N__65214),
            .I(N__65108));
    InMux I__13834 (
            .O(N__65213),
            .I(N__65108));
    InMux I__13833 (
            .O(N__65210),
            .I(N__65108));
    LocalMux I__13832 (
            .O(N__65197),
            .I(N__65105));
    InMux I__13831 (
            .O(N__65194),
            .I(N__65100));
    InMux I__13830 (
            .O(N__65191),
            .I(N__65100));
    CascadeMux I__13829 (
            .O(N__65190),
            .I(N__65096));
    CascadeMux I__13828 (
            .O(N__65189),
            .I(N__65093));
    InMux I__13827 (
            .O(N__65188),
            .I(N__65082));
    InMux I__13826 (
            .O(N__65187),
            .I(N__65082));
    InMux I__13825 (
            .O(N__65184),
            .I(N__65082));
    InMux I__13824 (
            .O(N__65183),
            .I(N__65082));
    InMux I__13823 (
            .O(N__65182),
            .I(N__65082));
    LocalMux I__13822 (
            .O(N__65177),
            .I(N__65078));
    InMux I__13821 (
            .O(N__65174),
            .I(N__65069));
    InMux I__13820 (
            .O(N__65173),
            .I(N__65069));
    InMux I__13819 (
            .O(N__65172),
            .I(N__65069));
    InMux I__13818 (
            .O(N__65169),
            .I(N__65069));
    InMux I__13817 (
            .O(N__65168),
            .I(N__65062));
    InMux I__13816 (
            .O(N__65167),
            .I(N__65062));
    InMux I__13815 (
            .O(N__65164),
            .I(N__65062));
    Span4Mux_s2_v I__13814 (
            .O(N__65161),
            .I(N__65055));
    LocalMux I__13813 (
            .O(N__65156),
            .I(N__65055));
    LocalMux I__13812 (
            .O(N__65149),
            .I(N__65055));
    LocalMux I__13811 (
            .O(N__65142),
            .I(N__65051));
    Span4Mux_s2_v I__13810 (
            .O(N__65139),
            .I(N__65048));
    LocalMux I__13809 (
            .O(N__65134),
            .I(N__65045));
    LocalMux I__13808 (
            .O(N__65121),
            .I(N__65036));
    LocalMux I__13807 (
            .O(N__65108),
            .I(N__65036));
    Span4Mux_v I__13806 (
            .O(N__65105),
            .I(N__65036));
    LocalMux I__13805 (
            .O(N__65100),
            .I(N__65036));
    InMux I__13804 (
            .O(N__65099),
            .I(N__65029));
    InMux I__13803 (
            .O(N__65096),
            .I(N__65029));
    InMux I__13802 (
            .O(N__65093),
            .I(N__65029));
    LocalMux I__13801 (
            .O(N__65082),
            .I(N__65026));
    InMux I__13800 (
            .O(N__65081),
            .I(N__65023));
    Span4Mux_v I__13799 (
            .O(N__65078),
            .I(N__65014));
    LocalMux I__13798 (
            .O(N__65069),
            .I(N__65014));
    LocalMux I__13797 (
            .O(N__65062),
            .I(N__65014));
    Span4Mux_v I__13796 (
            .O(N__65055),
            .I(N__65014));
    InMux I__13795 (
            .O(N__65054),
            .I(N__65011));
    Span4Mux_h I__13794 (
            .O(N__65051),
            .I(N__65008));
    Span4Mux_v I__13793 (
            .O(N__65048),
            .I(N__65001));
    Span4Mux_h I__13792 (
            .O(N__65045),
            .I(N__65001));
    Span4Mux_v I__13791 (
            .O(N__65036),
            .I(N__65001));
    LocalMux I__13790 (
            .O(N__65029),
            .I(N__64998));
    Span4Mux_v I__13789 (
            .O(N__65026),
            .I(N__64991));
    LocalMux I__13788 (
            .O(N__65023),
            .I(N__64991));
    Span4Mux_h I__13787 (
            .O(N__65014),
            .I(N__64991));
    LocalMux I__13786 (
            .O(N__65011),
            .I(N__64988));
    Span4Mux_s2_v I__13785 (
            .O(N__65008),
            .I(N__64985));
    Sp12to4 I__13784 (
            .O(N__65001),
            .I(N__64976));
    Span12Mux_s6_v I__13783 (
            .O(N__64998),
            .I(N__64976));
    Sp12to4 I__13782 (
            .O(N__64991),
            .I(N__64976));
    Span12Mux_h I__13781 (
            .O(N__64988),
            .I(N__64976));
    Odrv4 I__13780 (
            .O(N__64985),
            .I(pid_altitude_dv));
    Odrv12 I__13779 (
            .O(N__64976),
            .I(pid_altitude_dv));
    CEMux I__13778 (
            .O(N__64971),
            .I(N__64968));
    LocalMux I__13777 (
            .O(N__64968),
            .I(N__64965));
    Span4Mux_h I__13776 (
            .O(N__64965),
            .I(N__64962));
    Span4Mux_h I__13775 (
            .O(N__64962),
            .I(N__64959));
    Odrv4 I__13774 (
            .O(N__64959),
            .I(\pid_alt.state_1_0_0 ));
    InMux I__13773 (
            .O(N__64956),
            .I(\ppm_encoder_1.un1_counter_13_cry_2 ));
    InMux I__13772 (
            .O(N__64953),
            .I(N__64950));
    LocalMux I__13771 (
            .O(N__64950),
            .I(N__64947));
    Span4Mux_v I__13770 (
            .O(N__64947),
            .I(N__64942));
    InMux I__13769 (
            .O(N__64946),
            .I(N__64939));
    InMux I__13768 (
            .O(N__64945),
            .I(N__64936));
    Span4Mux_h I__13767 (
            .O(N__64942),
            .I(N__64931));
    LocalMux I__13766 (
            .O(N__64939),
            .I(N__64931));
    LocalMux I__13765 (
            .O(N__64936),
            .I(\ppm_encoder_1.counterZ0Z_4 ));
    Odrv4 I__13764 (
            .O(N__64931),
            .I(\ppm_encoder_1.counterZ0Z_4 ));
    InMux I__13763 (
            .O(N__64926),
            .I(\ppm_encoder_1.un1_counter_13_cry_3 ));
    InMux I__13762 (
            .O(N__64923),
            .I(N__64920));
    LocalMux I__13761 (
            .O(N__64920),
            .I(N__64917));
    Span4Mux_v I__13760 (
            .O(N__64917),
            .I(N__64912));
    InMux I__13759 (
            .O(N__64916),
            .I(N__64909));
    InMux I__13758 (
            .O(N__64915),
            .I(N__64906));
    Span4Mux_h I__13757 (
            .O(N__64912),
            .I(N__64901));
    LocalMux I__13756 (
            .O(N__64909),
            .I(N__64901));
    LocalMux I__13755 (
            .O(N__64906),
            .I(\ppm_encoder_1.counterZ0Z_5 ));
    Odrv4 I__13754 (
            .O(N__64901),
            .I(\ppm_encoder_1.counterZ0Z_5 ));
    InMux I__13753 (
            .O(N__64896),
            .I(\ppm_encoder_1.un1_counter_13_cry_4 ));
    InMux I__13752 (
            .O(N__64893),
            .I(N__64890));
    LocalMux I__13751 (
            .O(N__64890),
            .I(N__64886));
    InMux I__13750 (
            .O(N__64889),
            .I(N__64883));
    Span4Mux_v I__13749 (
            .O(N__64886),
            .I(N__64879));
    LocalMux I__13748 (
            .O(N__64883),
            .I(N__64876));
    InMux I__13747 (
            .O(N__64882),
            .I(N__64873));
    Span4Mux_h I__13746 (
            .O(N__64879),
            .I(N__64868));
    Span4Mux_h I__13745 (
            .O(N__64876),
            .I(N__64868));
    LocalMux I__13744 (
            .O(N__64873),
            .I(\ppm_encoder_1.counterZ0Z_6 ));
    Odrv4 I__13743 (
            .O(N__64868),
            .I(\ppm_encoder_1.counterZ0Z_6 ));
    InMux I__13742 (
            .O(N__64863),
            .I(\ppm_encoder_1.un1_counter_13_cry_5 ));
    CascadeMux I__13741 (
            .O(N__64860),
            .I(N__64857));
    InMux I__13740 (
            .O(N__64857),
            .I(N__64854));
    LocalMux I__13739 (
            .O(N__64854),
            .I(N__64851));
    Span4Mux_v I__13738 (
            .O(N__64851),
            .I(N__64847));
    InMux I__13737 (
            .O(N__64850),
            .I(N__64844));
    Span4Mux_h I__13736 (
            .O(N__64847),
            .I(N__64838));
    LocalMux I__13735 (
            .O(N__64844),
            .I(N__64838));
    InMux I__13734 (
            .O(N__64843),
            .I(N__64835));
    Span4Mux_h I__13733 (
            .O(N__64838),
            .I(N__64832));
    LocalMux I__13732 (
            .O(N__64835),
            .I(\ppm_encoder_1.counterZ0Z_7 ));
    Odrv4 I__13731 (
            .O(N__64832),
            .I(\ppm_encoder_1.counterZ0Z_7 ));
    InMux I__13730 (
            .O(N__64827),
            .I(\ppm_encoder_1.un1_counter_13_cry_6 ));
    InMux I__13729 (
            .O(N__64824),
            .I(N__64819));
    InMux I__13728 (
            .O(N__64823),
            .I(N__64816));
    InMux I__13727 (
            .O(N__64822),
            .I(N__64813));
    LocalMux I__13726 (
            .O(N__64819),
            .I(\ppm_encoder_1.counterZ0Z_8 ));
    LocalMux I__13725 (
            .O(N__64816),
            .I(\ppm_encoder_1.counterZ0Z_8 ));
    LocalMux I__13724 (
            .O(N__64813),
            .I(\ppm_encoder_1.counterZ0Z_8 ));
    InMux I__13723 (
            .O(N__64806),
            .I(bfn_16_5_0_));
    InMux I__13722 (
            .O(N__64803),
            .I(N__64798));
    InMux I__13721 (
            .O(N__64802),
            .I(N__64795));
    InMux I__13720 (
            .O(N__64801),
            .I(N__64792));
    LocalMux I__13719 (
            .O(N__64798),
            .I(\ppm_encoder_1.counterZ0Z_9 ));
    LocalMux I__13718 (
            .O(N__64795),
            .I(\ppm_encoder_1.counterZ0Z_9 ));
    LocalMux I__13717 (
            .O(N__64792),
            .I(\ppm_encoder_1.counterZ0Z_9 ));
    InMux I__13716 (
            .O(N__64785),
            .I(\ppm_encoder_1.un1_counter_13_cry_8 ));
    CascadeMux I__13715 (
            .O(N__64782),
            .I(N__64777));
    InMux I__13714 (
            .O(N__64781),
            .I(N__64774));
    InMux I__13713 (
            .O(N__64780),
            .I(N__64771));
    InMux I__13712 (
            .O(N__64777),
            .I(N__64768));
    LocalMux I__13711 (
            .O(N__64774),
            .I(\ppm_encoder_1.counterZ0Z_10 ));
    LocalMux I__13710 (
            .O(N__64771),
            .I(\ppm_encoder_1.counterZ0Z_10 ));
    LocalMux I__13709 (
            .O(N__64768),
            .I(\ppm_encoder_1.counterZ0Z_10 ));
    InMux I__13708 (
            .O(N__64761),
            .I(\ppm_encoder_1.un1_counter_13_cry_9 ));
    CascadeMux I__13707 (
            .O(N__64758),
            .I(N__64754));
    InMux I__13706 (
            .O(N__64757),
            .I(N__64750));
    InMux I__13705 (
            .O(N__64754),
            .I(N__64747));
    InMux I__13704 (
            .O(N__64753),
            .I(N__64744));
    LocalMux I__13703 (
            .O(N__64750),
            .I(\ppm_encoder_1.counterZ0Z_11 ));
    LocalMux I__13702 (
            .O(N__64747),
            .I(\ppm_encoder_1.counterZ0Z_11 ));
    LocalMux I__13701 (
            .O(N__64744),
            .I(\ppm_encoder_1.counterZ0Z_11 ));
    InMux I__13700 (
            .O(N__64737),
            .I(N__64734));
    LocalMux I__13699 (
            .O(N__64734),
            .I(\ppm_encoder_1.pulses2countZ0Z_0 ));
    InMux I__13698 (
            .O(N__64731),
            .I(N__64728));
    LocalMux I__13697 (
            .O(N__64728),
            .I(N__64725));
    Span4Mux_s2_v I__13696 (
            .O(N__64725),
            .I(N__64722));
    Odrv4 I__13695 (
            .O(N__64722),
            .I(\ppm_encoder_1.counter24_0_I_1_c_RNOZ0 ));
    InMux I__13694 (
            .O(N__64719),
            .I(N__64716));
    LocalMux I__13693 (
            .O(N__64716),
            .I(N__64713));
    Span4Mux_s3_v I__13692 (
            .O(N__64713),
            .I(N__64710));
    Span4Mux_h I__13691 (
            .O(N__64710),
            .I(N__64707));
    Odrv4 I__13690 (
            .O(N__64707),
            .I(\ppm_encoder_1.pulses2count_9_0_3_1 ));
    CascadeMux I__13689 (
            .O(N__64704),
            .I(N__64701));
    InMux I__13688 (
            .O(N__64701),
            .I(N__64698));
    LocalMux I__13687 (
            .O(N__64698),
            .I(N__64695));
    Span4Mux_h I__13686 (
            .O(N__64695),
            .I(N__64692));
    Odrv4 I__13685 (
            .O(N__64692),
            .I(\ppm_encoder_1.pulses2count_9_0_0_1 ));
    InMux I__13684 (
            .O(N__64689),
            .I(N__64686));
    LocalMux I__13683 (
            .O(N__64686),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_1 ));
    CascadeMux I__13682 (
            .O(N__64683),
            .I(N__64680));
    InMux I__13681 (
            .O(N__64680),
            .I(N__64677));
    LocalMux I__13680 (
            .O(N__64677),
            .I(\ppm_encoder_1.pulses2countZ0Z_1 ));
    InMux I__13679 (
            .O(N__64674),
            .I(N__64670));
    CascadeMux I__13678 (
            .O(N__64673),
            .I(N__64666));
    LocalMux I__13677 (
            .O(N__64670),
            .I(N__64663));
    InMux I__13676 (
            .O(N__64669),
            .I(N__64658));
    InMux I__13675 (
            .O(N__64666),
            .I(N__64658));
    Span4Mux_s3_v I__13674 (
            .O(N__64663),
            .I(N__64655));
    LocalMux I__13673 (
            .O(N__64658),
            .I(N__64651));
    Span4Mux_h I__13672 (
            .O(N__64655),
            .I(N__64648));
    InMux I__13671 (
            .O(N__64654),
            .I(N__64645));
    Span4Mux_s1_v I__13670 (
            .O(N__64651),
            .I(N__64642));
    Odrv4 I__13669 (
            .O(N__64648),
            .I(\ppm_encoder_1.init_pulsesZ0Z_15 ));
    LocalMux I__13668 (
            .O(N__64645),
            .I(\ppm_encoder_1.init_pulsesZ0Z_15 ));
    Odrv4 I__13667 (
            .O(N__64642),
            .I(\ppm_encoder_1.init_pulsesZ0Z_15 ));
    CascadeMux I__13666 (
            .O(N__64635),
            .I(N__64631));
    InMux I__13665 (
            .O(N__64634),
            .I(N__64628));
    InMux I__13664 (
            .O(N__64631),
            .I(N__64625));
    LocalMux I__13663 (
            .O(N__64628),
            .I(N__64622));
    LocalMux I__13662 (
            .O(N__64625),
            .I(N__64619));
    Span12Mux_s3_v I__13661 (
            .O(N__64622),
            .I(N__64615));
    Span4Mux_v I__13660 (
            .O(N__64619),
            .I(N__64612));
    InMux I__13659 (
            .O(N__64618),
            .I(N__64609));
    Odrv12 I__13658 (
            .O(N__64615),
            .I(\ppm_encoder_1.init_pulsesZ0Z_17 ));
    Odrv4 I__13657 (
            .O(N__64612),
            .I(\ppm_encoder_1.init_pulsesZ0Z_17 ));
    LocalMux I__13656 (
            .O(N__64609),
            .I(\ppm_encoder_1.init_pulsesZ0Z_17 ));
    CascadeMux I__13655 (
            .O(N__64602),
            .I(N__64592));
    CascadeMux I__13654 (
            .O(N__64601),
            .I(N__64587));
    InMux I__13653 (
            .O(N__64600),
            .I(N__64577));
    InMux I__13652 (
            .O(N__64599),
            .I(N__64577));
    InMux I__13651 (
            .O(N__64598),
            .I(N__64573));
    InMux I__13650 (
            .O(N__64597),
            .I(N__64570));
    InMux I__13649 (
            .O(N__64596),
            .I(N__64565));
    InMux I__13648 (
            .O(N__64595),
            .I(N__64565));
    InMux I__13647 (
            .O(N__64592),
            .I(N__64562));
    InMux I__13646 (
            .O(N__64591),
            .I(N__64557));
    InMux I__13645 (
            .O(N__64590),
            .I(N__64557));
    InMux I__13644 (
            .O(N__64587),
            .I(N__64552));
    InMux I__13643 (
            .O(N__64586),
            .I(N__64552));
    CascadeMux I__13642 (
            .O(N__64585),
            .I(N__64549));
    InMux I__13641 (
            .O(N__64584),
            .I(N__64543));
    InMux I__13640 (
            .O(N__64583),
            .I(N__64538));
    InMux I__13639 (
            .O(N__64582),
            .I(N__64538));
    LocalMux I__13638 (
            .O(N__64577),
            .I(N__64535));
    InMux I__13637 (
            .O(N__64576),
            .I(N__64532));
    LocalMux I__13636 (
            .O(N__64573),
            .I(N__64527));
    LocalMux I__13635 (
            .O(N__64570),
            .I(N__64527));
    LocalMux I__13634 (
            .O(N__64565),
            .I(N__64524));
    LocalMux I__13633 (
            .O(N__64562),
            .I(N__64521));
    LocalMux I__13632 (
            .O(N__64557),
            .I(N__64517));
    LocalMux I__13631 (
            .O(N__64552),
            .I(N__64514));
    InMux I__13630 (
            .O(N__64549),
            .I(N__64505));
    InMux I__13629 (
            .O(N__64548),
            .I(N__64505));
    InMux I__13628 (
            .O(N__64547),
            .I(N__64505));
    InMux I__13627 (
            .O(N__64546),
            .I(N__64505));
    LocalMux I__13626 (
            .O(N__64543),
            .I(N__64495));
    LocalMux I__13625 (
            .O(N__64538),
            .I(N__64495));
    Span4Mux_h I__13624 (
            .O(N__64535),
            .I(N__64495));
    LocalMux I__13623 (
            .O(N__64532),
            .I(N__64495));
    Span4Mux_v I__13622 (
            .O(N__64527),
            .I(N__64488));
    Span4Mux_v I__13621 (
            .O(N__64524),
            .I(N__64488));
    Span4Mux_s1_v I__13620 (
            .O(N__64521),
            .I(N__64488));
    CascadeMux I__13619 (
            .O(N__64520),
            .I(N__64484));
    Span4Mux_v I__13618 (
            .O(N__64517),
            .I(N__64479));
    Span4Mux_s1_v I__13617 (
            .O(N__64514),
            .I(N__64479));
    LocalMux I__13616 (
            .O(N__64505),
            .I(N__64476));
    InMux I__13615 (
            .O(N__64504),
            .I(N__64473));
    Span4Mux_v I__13614 (
            .O(N__64495),
            .I(N__64468));
    Span4Mux_h I__13613 (
            .O(N__64488),
            .I(N__64468));
    InMux I__13612 (
            .O(N__64487),
            .I(N__64463));
    InMux I__13611 (
            .O(N__64484),
            .I(N__64463));
    Span4Mux_h I__13610 (
            .O(N__64479),
            .I(N__64458));
    Span4Mux_h I__13609 (
            .O(N__64476),
            .I(N__64458));
    LocalMux I__13608 (
            .O(N__64473),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_3 ));
    Odrv4 I__13607 (
            .O(N__64468),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_3 ));
    LocalMux I__13606 (
            .O(N__64463),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_3 ));
    Odrv4 I__13605 (
            .O(N__64458),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_3 ));
    CascadeMux I__13604 (
            .O(N__64449),
            .I(N__64445));
    CascadeMux I__13603 (
            .O(N__64448),
            .I(N__64438));
    InMux I__13602 (
            .O(N__64445),
            .I(N__64432));
    InMux I__13601 (
            .O(N__64444),
            .I(N__64428));
    InMux I__13600 (
            .O(N__64443),
            .I(N__64423));
    InMux I__13599 (
            .O(N__64442),
            .I(N__64423));
    InMux I__13598 (
            .O(N__64441),
            .I(N__64420));
    InMux I__13597 (
            .O(N__64438),
            .I(N__64411));
    InMux I__13596 (
            .O(N__64437),
            .I(N__64411));
    InMux I__13595 (
            .O(N__64436),
            .I(N__64411));
    InMux I__13594 (
            .O(N__64435),
            .I(N__64411));
    LocalMux I__13593 (
            .O(N__64432),
            .I(N__64408));
    InMux I__13592 (
            .O(N__64431),
            .I(N__64405));
    LocalMux I__13591 (
            .O(N__64428),
            .I(N__64402));
    LocalMux I__13590 (
            .O(N__64423),
            .I(N__64399));
    LocalMux I__13589 (
            .O(N__64420),
            .I(N__64392));
    LocalMux I__13588 (
            .O(N__64411),
            .I(N__64377));
    Span4Mux_h I__13587 (
            .O(N__64408),
            .I(N__64377));
    LocalMux I__13586 (
            .O(N__64405),
            .I(N__64377));
    Span4Mux_h I__13585 (
            .O(N__64402),
            .I(N__64377));
    Span4Mux_h I__13584 (
            .O(N__64399),
            .I(N__64377));
    InMux I__13583 (
            .O(N__64398),
            .I(N__64374));
    InMux I__13582 (
            .O(N__64397),
            .I(N__64371));
    InMux I__13581 (
            .O(N__64396),
            .I(N__64366));
    InMux I__13580 (
            .O(N__64395),
            .I(N__64366));
    Span4Mux_v I__13579 (
            .O(N__64392),
            .I(N__64363));
    InMux I__13578 (
            .O(N__64391),
            .I(N__64358));
    InMux I__13577 (
            .O(N__64390),
            .I(N__64358));
    InMux I__13576 (
            .O(N__64389),
            .I(N__64353));
    InMux I__13575 (
            .O(N__64388),
            .I(N__64353));
    Span4Mux_v I__13574 (
            .O(N__64377),
            .I(N__64350));
    LocalMux I__13573 (
            .O(N__64374),
            .I(N__64347));
    LocalMux I__13572 (
            .O(N__64371),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNISSERZ0 ));
    LocalMux I__13571 (
            .O(N__64366),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNISSERZ0 ));
    Odrv4 I__13570 (
            .O(N__64363),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNISSERZ0 ));
    LocalMux I__13569 (
            .O(N__64358),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNISSERZ0 ));
    LocalMux I__13568 (
            .O(N__64353),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNISSERZ0 ));
    Odrv4 I__13567 (
            .O(N__64350),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNISSERZ0 ));
    Odrv4 I__13566 (
            .O(N__64347),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNISSERZ0 ));
    InMux I__13565 (
            .O(N__64332),
            .I(N__64329));
    LocalMux I__13564 (
            .O(N__64329),
            .I(N__64326));
    Odrv4 I__13563 (
            .O(N__64326),
            .I(\ppm_encoder_1.pulses2countZ0Z_16 ));
    CascadeMux I__13562 (
            .O(N__64323),
            .I(N__64320));
    InMux I__13561 (
            .O(N__64320),
            .I(N__64317));
    LocalMux I__13560 (
            .O(N__64317),
            .I(\ppm_encoder_1.pulses2countZ0Z_17 ));
    InMux I__13559 (
            .O(N__64314),
            .I(N__64311));
    LocalMux I__13558 (
            .O(N__64311),
            .I(N__64308));
    Odrv4 I__13557 (
            .O(N__64308),
            .I(\ppm_encoder_1.counter24_0_I_51_c_RNOZ0 ));
    CascadeMux I__13556 (
            .O(N__64305),
            .I(N__64299));
    CascadeMux I__13555 (
            .O(N__64304),
            .I(N__64296));
    InMux I__13554 (
            .O(N__64303),
            .I(N__64281));
    InMux I__13553 (
            .O(N__64302),
            .I(N__64281));
    InMux I__13552 (
            .O(N__64299),
            .I(N__64278));
    InMux I__13551 (
            .O(N__64296),
            .I(N__64275));
    InMux I__13550 (
            .O(N__64295),
            .I(N__64248));
    InMux I__13549 (
            .O(N__64294),
            .I(N__64248));
    InMux I__13548 (
            .O(N__64293),
            .I(N__64248));
    InMux I__13547 (
            .O(N__64292),
            .I(N__64243));
    InMux I__13546 (
            .O(N__64291),
            .I(N__64243));
    InMux I__13545 (
            .O(N__64290),
            .I(N__64240));
    InMux I__13544 (
            .O(N__64289),
            .I(N__64234));
    InMux I__13543 (
            .O(N__64288),
            .I(N__64234));
    InMux I__13542 (
            .O(N__64287),
            .I(N__64225));
    InMux I__13541 (
            .O(N__64286),
            .I(N__64225));
    LocalMux I__13540 (
            .O(N__64281),
            .I(N__64218));
    LocalMux I__13539 (
            .O(N__64278),
            .I(N__64218));
    LocalMux I__13538 (
            .O(N__64275),
            .I(N__64218));
    InMux I__13537 (
            .O(N__64274),
            .I(N__64211));
    InMux I__13536 (
            .O(N__64273),
            .I(N__64211));
    InMux I__13535 (
            .O(N__64272),
            .I(N__64211));
    InMux I__13534 (
            .O(N__64271),
            .I(N__64206));
    InMux I__13533 (
            .O(N__64270),
            .I(N__64206));
    InMux I__13532 (
            .O(N__64269),
            .I(N__64201));
    InMux I__13531 (
            .O(N__64268),
            .I(N__64201));
    InMux I__13530 (
            .O(N__64267),
            .I(N__64192));
    InMux I__13529 (
            .O(N__64266),
            .I(N__64192));
    InMux I__13528 (
            .O(N__64265),
            .I(N__64192));
    InMux I__13527 (
            .O(N__64264),
            .I(N__64192));
    InMux I__13526 (
            .O(N__64263),
            .I(N__64185));
    InMux I__13525 (
            .O(N__64262),
            .I(N__64185));
    InMux I__13524 (
            .O(N__64261),
            .I(N__64185));
    InMux I__13523 (
            .O(N__64260),
            .I(N__64176));
    InMux I__13522 (
            .O(N__64259),
            .I(N__64176));
    InMux I__13521 (
            .O(N__64258),
            .I(N__64176));
    InMux I__13520 (
            .O(N__64257),
            .I(N__64176));
    InMux I__13519 (
            .O(N__64256),
            .I(N__64173));
    CascadeMux I__13518 (
            .O(N__64255),
            .I(N__64169));
    LocalMux I__13517 (
            .O(N__64248),
            .I(N__64161));
    LocalMux I__13516 (
            .O(N__64243),
            .I(N__64158));
    LocalMux I__13515 (
            .O(N__64240),
            .I(N__64155));
    InMux I__13514 (
            .O(N__64239),
            .I(N__64152));
    LocalMux I__13513 (
            .O(N__64234),
            .I(N__64149));
    InMux I__13512 (
            .O(N__64233),
            .I(N__64137));
    InMux I__13511 (
            .O(N__64232),
            .I(N__64137));
    InMux I__13510 (
            .O(N__64231),
            .I(N__64137));
    InMux I__13509 (
            .O(N__64230),
            .I(N__64137));
    LocalMux I__13508 (
            .O(N__64225),
            .I(N__64128));
    Span4Mux_v I__13507 (
            .O(N__64218),
            .I(N__64128));
    LocalMux I__13506 (
            .O(N__64211),
            .I(N__64128));
    LocalMux I__13505 (
            .O(N__64206),
            .I(N__64128));
    LocalMux I__13504 (
            .O(N__64201),
            .I(N__64123));
    LocalMux I__13503 (
            .O(N__64192),
            .I(N__64123));
    LocalMux I__13502 (
            .O(N__64185),
            .I(N__64116));
    LocalMux I__13501 (
            .O(N__64176),
            .I(N__64116));
    LocalMux I__13500 (
            .O(N__64173),
            .I(N__64116));
    InMux I__13499 (
            .O(N__64172),
            .I(N__64113));
    InMux I__13498 (
            .O(N__64169),
            .I(N__64110));
    InMux I__13497 (
            .O(N__64168),
            .I(N__64105));
    InMux I__13496 (
            .O(N__64167),
            .I(N__64105));
    InMux I__13495 (
            .O(N__64166),
            .I(N__64094));
    InMux I__13494 (
            .O(N__64165),
            .I(N__64094));
    InMux I__13493 (
            .O(N__64164),
            .I(N__64094));
    Span4Mux_h I__13492 (
            .O(N__64161),
            .I(N__64091));
    Span4Mux_v I__13491 (
            .O(N__64158),
            .I(N__64082));
    Span4Mux_v I__13490 (
            .O(N__64155),
            .I(N__64082));
    LocalMux I__13489 (
            .O(N__64152),
            .I(N__64082));
    Span4Mux_s3_v I__13488 (
            .O(N__64149),
            .I(N__64082));
    InMux I__13487 (
            .O(N__64148),
            .I(N__64079));
    InMux I__13486 (
            .O(N__64147),
            .I(N__64074));
    InMux I__13485 (
            .O(N__64146),
            .I(N__64074));
    LocalMux I__13484 (
            .O(N__64137),
            .I(N__64067));
    Span4Mux_h I__13483 (
            .O(N__64128),
            .I(N__64067));
    Span4Mux_s0_v I__13482 (
            .O(N__64123),
            .I(N__64067));
    Span4Mux_s3_v I__13481 (
            .O(N__64116),
            .I(N__64064));
    LocalMux I__13480 (
            .O(N__64113),
            .I(N__64057));
    LocalMux I__13479 (
            .O(N__64110),
            .I(N__64057));
    LocalMux I__13478 (
            .O(N__64105),
            .I(N__64057));
    InMux I__13477 (
            .O(N__64104),
            .I(N__64050));
    InMux I__13476 (
            .O(N__64103),
            .I(N__64050));
    InMux I__13475 (
            .O(N__64102),
            .I(N__64050));
    InMux I__13474 (
            .O(N__64101),
            .I(N__64047));
    LocalMux I__13473 (
            .O(N__64094),
            .I(\ppm_encoder_1.PPM_STATE_RNIV4V5Z0Z_1 ));
    Odrv4 I__13472 (
            .O(N__64091),
            .I(\ppm_encoder_1.PPM_STATE_RNIV4V5Z0Z_1 ));
    Odrv4 I__13471 (
            .O(N__64082),
            .I(\ppm_encoder_1.PPM_STATE_RNIV4V5Z0Z_1 ));
    LocalMux I__13470 (
            .O(N__64079),
            .I(\ppm_encoder_1.PPM_STATE_RNIV4V5Z0Z_1 ));
    LocalMux I__13469 (
            .O(N__64074),
            .I(\ppm_encoder_1.PPM_STATE_RNIV4V5Z0Z_1 ));
    Odrv4 I__13468 (
            .O(N__64067),
            .I(\ppm_encoder_1.PPM_STATE_RNIV4V5Z0Z_1 ));
    Odrv4 I__13467 (
            .O(N__64064),
            .I(\ppm_encoder_1.PPM_STATE_RNIV4V5Z0Z_1 ));
    Odrv12 I__13466 (
            .O(N__64057),
            .I(\ppm_encoder_1.PPM_STATE_RNIV4V5Z0Z_1 ));
    LocalMux I__13465 (
            .O(N__64050),
            .I(\ppm_encoder_1.PPM_STATE_RNIV4V5Z0Z_1 ));
    LocalMux I__13464 (
            .O(N__64047),
            .I(\ppm_encoder_1.PPM_STATE_RNIV4V5Z0Z_1 ));
    InMux I__13463 (
            .O(N__64026),
            .I(N__64023));
    LocalMux I__13462 (
            .O(N__64023),
            .I(N__64020));
    Span4Mux_v I__13461 (
            .O(N__64020),
            .I(N__64016));
    InMux I__13460 (
            .O(N__64019),
            .I(N__64012));
    Span4Mux_v I__13459 (
            .O(N__64016),
            .I(N__64009));
    InMux I__13458 (
            .O(N__64015),
            .I(N__64006));
    LocalMux I__13457 (
            .O(N__64012),
            .I(\ppm_encoder_1.counterZ0Z_0 ));
    Odrv4 I__13456 (
            .O(N__64009),
            .I(\ppm_encoder_1.counterZ0Z_0 ));
    LocalMux I__13455 (
            .O(N__64006),
            .I(\ppm_encoder_1.counterZ0Z_0 ));
    InMux I__13454 (
            .O(N__63999),
            .I(N__63996));
    LocalMux I__13453 (
            .O(N__63996),
            .I(N__63993));
    Span4Mux_v I__13452 (
            .O(N__63993),
            .I(N__63989));
    InMux I__13451 (
            .O(N__63992),
            .I(N__63985));
    Span4Mux_v I__13450 (
            .O(N__63989),
            .I(N__63982));
    InMux I__13449 (
            .O(N__63988),
            .I(N__63979));
    LocalMux I__13448 (
            .O(N__63985),
            .I(\ppm_encoder_1.counterZ0Z_1 ));
    Odrv4 I__13447 (
            .O(N__63982),
            .I(\ppm_encoder_1.counterZ0Z_1 ));
    LocalMux I__13446 (
            .O(N__63979),
            .I(\ppm_encoder_1.counterZ0Z_1 ));
    InMux I__13445 (
            .O(N__63972),
            .I(\ppm_encoder_1.un1_counter_13_cry_0 ));
    InMux I__13444 (
            .O(N__63969),
            .I(\ppm_encoder_1.un1_counter_13_cry_1 ));
    InMux I__13443 (
            .O(N__63966),
            .I(N__63963));
    LocalMux I__13442 (
            .O(N__63963),
            .I(N__63960));
    Odrv12 I__13441 (
            .O(N__63960),
            .I(\pid_front.error_i_reg_9_rn_0_26 ));
    CascadeMux I__13440 (
            .O(N__63957),
            .I(N__63954));
    InMux I__13439 (
            .O(N__63954),
            .I(N__63951));
    LocalMux I__13438 (
            .O(N__63951),
            .I(N__63948));
    Span4Mux_h I__13437 (
            .O(N__63948),
            .I(N__63945));
    Odrv4 I__13436 (
            .O(N__63945),
            .I(\pid_front.error_i_regZ0Z_26 ));
    InMux I__13435 (
            .O(N__63942),
            .I(N__63939));
    LocalMux I__13434 (
            .O(N__63939),
            .I(N__63936));
    Span4Mux_s0_v I__13433 (
            .O(N__63936),
            .I(N__63932));
    CascadeMux I__13432 (
            .O(N__63935),
            .I(N__63929));
    Span4Mux_h I__13431 (
            .O(N__63932),
            .I(N__63925));
    InMux I__13430 (
            .O(N__63929),
            .I(N__63922));
    InMux I__13429 (
            .O(N__63928),
            .I(N__63919));
    Odrv4 I__13428 (
            .O(N__63925),
            .I(\ppm_encoder_1.init_pulsesZ0Z_16 ));
    LocalMux I__13427 (
            .O(N__63922),
            .I(\ppm_encoder_1.init_pulsesZ0Z_16 ));
    LocalMux I__13426 (
            .O(N__63919),
            .I(\ppm_encoder_1.init_pulsesZ0Z_16 ));
    CascadeMux I__13425 (
            .O(N__63912),
            .I(N__63909));
    InMux I__13424 (
            .O(N__63909),
            .I(N__63904));
    InMux I__13423 (
            .O(N__63908),
            .I(N__63900));
    InMux I__13422 (
            .O(N__63907),
            .I(N__63897));
    LocalMux I__13421 (
            .O(N__63904),
            .I(N__63894));
    CascadeMux I__13420 (
            .O(N__63903),
            .I(N__63891));
    LocalMux I__13419 (
            .O(N__63900),
            .I(N__63888));
    LocalMux I__13418 (
            .O(N__63897),
            .I(N__63885));
    Span4Mux_h I__13417 (
            .O(N__63894),
            .I(N__63882));
    InMux I__13416 (
            .O(N__63891),
            .I(N__63879));
    Span4Mux_h I__13415 (
            .O(N__63888),
            .I(N__63874));
    Span4Mux_h I__13414 (
            .O(N__63885),
            .I(N__63874));
    Span4Mux_v I__13413 (
            .O(N__63882),
            .I(N__63869));
    LocalMux I__13412 (
            .O(N__63879),
            .I(N__63869));
    Odrv4 I__13411 (
            .O(N__63874),
            .I(\ppm_encoder_1.m9_0_i ));
    Odrv4 I__13410 (
            .O(N__63869),
            .I(\ppm_encoder_1.m9_0_i ));
    InMux I__13409 (
            .O(N__63864),
            .I(N__63861));
    LocalMux I__13408 (
            .O(N__63861),
            .I(N__63854));
    InMux I__13407 (
            .O(N__63860),
            .I(N__63851));
    InMux I__13406 (
            .O(N__63859),
            .I(N__63848));
    InMux I__13405 (
            .O(N__63858),
            .I(N__63844));
    InMux I__13404 (
            .O(N__63857),
            .I(N__63841));
    Span4Mux_v I__13403 (
            .O(N__63854),
            .I(N__63836));
    LocalMux I__13402 (
            .O(N__63851),
            .I(N__63836));
    LocalMux I__13401 (
            .O(N__63848),
            .I(N__63833));
    CascadeMux I__13400 (
            .O(N__63847),
            .I(N__63830));
    LocalMux I__13399 (
            .O(N__63844),
            .I(N__63827));
    LocalMux I__13398 (
            .O(N__63841),
            .I(N__63824));
    Span4Mux_h I__13397 (
            .O(N__63836),
            .I(N__63819));
    Span4Mux_h I__13396 (
            .O(N__63833),
            .I(N__63819));
    InMux I__13395 (
            .O(N__63830),
            .I(N__63816));
    Odrv4 I__13394 (
            .O(N__63827),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIHO7DZ0Z_0 ));
    Odrv12 I__13393 (
            .O(N__63824),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIHO7DZ0Z_0 ));
    Odrv4 I__13392 (
            .O(N__63819),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIHO7DZ0Z_0 ));
    LocalMux I__13391 (
            .O(N__63816),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIHO7DZ0Z_0 ));
    InMux I__13390 (
            .O(N__63807),
            .I(N__63798));
    InMux I__13389 (
            .O(N__63806),
            .I(N__63798));
    InMux I__13388 (
            .O(N__63805),
            .I(N__63790));
    InMux I__13387 (
            .O(N__63804),
            .I(N__63783));
    InMux I__13386 (
            .O(N__63803),
            .I(N__63783));
    LocalMux I__13385 (
            .O(N__63798),
            .I(N__63780));
    InMux I__13384 (
            .O(N__63797),
            .I(N__63776));
    InMux I__13383 (
            .O(N__63796),
            .I(N__63771));
    InMux I__13382 (
            .O(N__63795),
            .I(N__63771));
    InMux I__13381 (
            .O(N__63794),
            .I(N__63766));
    InMux I__13380 (
            .O(N__63793),
            .I(N__63766));
    LocalMux I__13379 (
            .O(N__63790),
            .I(N__63763));
    InMux I__13378 (
            .O(N__63789),
            .I(N__63758));
    InMux I__13377 (
            .O(N__63788),
            .I(N__63758));
    LocalMux I__13376 (
            .O(N__63783),
            .I(N__63753));
    Span4Mux_s3_v I__13375 (
            .O(N__63780),
            .I(N__63750));
    InMux I__13374 (
            .O(N__63779),
            .I(N__63747));
    LocalMux I__13373 (
            .O(N__63776),
            .I(N__63742));
    LocalMux I__13372 (
            .O(N__63771),
            .I(N__63742));
    LocalMux I__13371 (
            .O(N__63766),
            .I(N__63738));
    Span4Mux_v I__13370 (
            .O(N__63763),
            .I(N__63733));
    LocalMux I__13369 (
            .O(N__63758),
            .I(N__63733));
    InMux I__13368 (
            .O(N__63757),
            .I(N__63730));
    InMux I__13367 (
            .O(N__63756),
            .I(N__63727));
    Span4Mux_s3_v I__13366 (
            .O(N__63753),
            .I(N__63722));
    Span4Mux_h I__13365 (
            .O(N__63750),
            .I(N__63722));
    LocalMux I__13364 (
            .O(N__63747),
            .I(N__63717));
    Span4Mux_h I__13363 (
            .O(N__63742),
            .I(N__63717));
    InMux I__13362 (
            .O(N__63741),
            .I(N__63714));
    Span4Mux_v I__13361 (
            .O(N__63738),
            .I(N__63709));
    Span4Mux_h I__13360 (
            .O(N__63733),
            .I(N__63709));
    LocalMux I__13359 (
            .O(N__63730),
            .I(N__63706));
    LocalMux I__13358 (
            .O(N__63727),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z1 ));
    Odrv4 I__13357 (
            .O(N__63722),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z1 ));
    Odrv4 I__13356 (
            .O(N__63717),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z1 ));
    LocalMux I__13355 (
            .O(N__63714),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z1 ));
    Odrv4 I__13354 (
            .O(N__63709),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z1 ));
    Odrv12 I__13353 (
            .O(N__63706),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z1 ));
    CascadeMux I__13352 (
            .O(N__63693),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNISSERZ0_cascade_ ));
    CascadeMux I__13351 (
            .O(N__63690),
            .I(N__63686));
    InMux I__13350 (
            .O(N__63689),
            .I(N__63683));
    InMux I__13349 (
            .O(N__63686),
            .I(N__63679));
    LocalMux I__13348 (
            .O(N__63683),
            .I(N__63676));
    InMux I__13347 (
            .O(N__63682),
            .I(N__63672));
    LocalMux I__13346 (
            .O(N__63679),
            .I(N__63669));
    Span4Mux_s3_v I__13345 (
            .O(N__63676),
            .I(N__63666));
    InMux I__13344 (
            .O(N__63675),
            .I(N__63663));
    LocalMux I__13343 (
            .O(N__63672),
            .I(N__63660));
    Span4Mux_h I__13342 (
            .O(N__63669),
            .I(N__63657));
    Sp12to4 I__13341 (
            .O(N__63666),
            .I(N__63652));
    LocalMux I__13340 (
            .O(N__63663),
            .I(N__63652));
    Odrv4 I__13339 (
            .O(N__63660),
            .I(\ppm_encoder_1.init_pulsesZ0Z_1 ));
    Odrv4 I__13338 (
            .O(N__63657),
            .I(\ppm_encoder_1.init_pulsesZ0Z_1 ));
    Odrv12 I__13337 (
            .O(N__63652),
            .I(\ppm_encoder_1.init_pulsesZ0Z_1 ));
    InMux I__13336 (
            .O(N__63645),
            .I(N__63641));
    CascadeMux I__13335 (
            .O(N__63644),
            .I(N__63638));
    LocalMux I__13334 (
            .O(N__63641),
            .I(N__63635));
    InMux I__13333 (
            .O(N__63638),
            .I(N__63632));
    Span4Mux_v I__13332 (
            .O(N__63635),
            .I(N__63629));
    LocalMux I__13331 (
            .O(N__63632),
            .I(N__63626));
    Odrv4 I__13330 (
            .O(N__63629),
            .I(\ppm_encoder_1.init_pulsesZ0Z_0 ));
    Odrv12 I__13329 (
            .O(N__63626),
            .I(\ppm_encoder_1.init_pulsesZ0Z_0 ));
    InMux I__13328 (
            .O(N__63621),
            .I(N__63618));
    LocalMux I__13327 (
            .O(N__63618),
            .I(N__63614));
    CascadeMux I__13326 (
            .O(N__63617),
            .I(N__63610));
    Span4Mux_s2_v I__13325 (
            .O(N__63614),
            .I(N__63607));
    InMux I__13324 (
            .O(N__63613),
            .I(N__63602));
    InMux I__13323 (
            .O(N__63610),
            .I(N__63602));
    Odrv4 I__13322 (
            .O(N__63607),
            .I(\ppm_encoder_1.elevatorZ0Z_0 ));
    LocalMux I__13321 (
            .O(N__63602),
            .I(\ppm_encoder_1.elevatorZ0Z_0 ));
    CascadeMux I__13320 (
            .O(N__63597),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_2Z0Z_0_cascade_ ));
    InMux I__13319 (
            .O(N__63594),
            .I(N__63585));
    InMux I__13318 (
            .O(N__63593),
            .I(N__63581));
    InMux I__13317 (
            .O(N__63592),
            .I(N__63576));
    InMux I__13316 (
            .O(N__63591),
            .I(N__63576));
    InMux I__13315 (
            .O(N__63590),
            .I(N__63573));
    InMux I__13314 (
            .O(N__63589),
            .I(N__63568));
    InMux I__13313 (
            .O(N__63588),
            .I(N__63568));
    LocalMux I__13312 (
            .O(N__63585),
            .I(N__63565));
    InMux I__13311 (
            .O(N__63584),
            .I(N__63562));
    LocalMux I__13310 (
            .O(N__63581),
            .I(N__63559));
    LocalMux I__13309 (
            .O(N__63576),
            .I(N__63556));
    LocalMux I__13308 (
            .O(N__63573),
            .I(N__63552));
    LocalMux I__13307 (
            .O(N__63568),
            .I(N__63549));
    Span4Mux_v I__13306 (
            .O(N__63565),
            .I(N__63546));
    LocalMux I__13305 (
            .O(N__63562),
            .I(N__63539));
    Span4Mux_h I__13304 (
            .O(N__63559),
            .I(N__63539));
    Span4Mux_h I__13303 (
            .O(N__63556),
            .I(N__63536));
    InMux I__13302 (
            .O(N__63555),
            .I(N__63533));
    Span4Mux_v I__13301 (
            .O(N__63552),
            .I(N__63526));
    Span4Mux_v I__13300 (
            .O(N__63549),
            .I(N__63526));
    Span4Mux_h I__13299 (
            .O(N__63546),
            .I(N__63526));
    InMux I__13298 (
            .O(N__63545),
            .I(N__63521));
    InMux I__13297 (
            .O(N__63544),
            .I(N__63521));
    Odrv4 I__13296 (
            .O(N__63539),
            .I(\ppm_encoder_1.m9_0_i_o2 ));
    Odrv4 I__13295 (
            .O(N__63536),
            .I(\ppm_encoder_1.m9_0_i_o2 ));
    LocalMux I__13294 (
            .O(N__63533),
            .I(\ppm_encoder_1.m9_0_i_o2 ));
    Odrv4 I__13293 (
            .O(N__63526),
            .I(\ppm_encoder_1.m9_0_i_o2 ));
    LocalMux I__13292 (
            .O(N__63521),
            .I(\ppm_encoder_1.m9_0_i_o2 ));
    InMux I__13291 (
            .O(N__63510),
            .I(N__63507));
    LocalMux I__13290 (
            .O(N__63507),
            .I(\ppm_encoder_1.pulses2count_9_0_2_0 ));
    InMux I__13289 (
            .O(N__63504),
            .I(N__63501));
    LocalMux I__13288 (
            .O(N__63501),
            .I(N__63495));
    CascadeMux I__13287 (
            .O(N__63500),
            .I(N__63492));
    CascadeMux I__13286 (
            .O(N__63499),
            .I(N__63489));
    InMux I__13285 (
            .O(N__63498),
            .I(N__63486));
    Span4Mux_h I__13284 (
            .O(N__63495),
            .I(N__63483));
    InMux I__13283 (
            .O(N__63492),
            .I(N__63478));
    InMux I__13282 (
            .O(N__63489),
            .I(N__63478));
    LocalMux I__13281 (
            .O(N__63486),
            .I(N__63475));
    Span4Mux_h I__13280 (
            .O(N__63483),
            .I(N__63470));
    LocalMux I__13279 (
            .O(N__63478),
            .I(N__63470));
    Odrv12 I__13278 (
            .O(N__63475),
            .I(\ppm_encoder_1.init_pulsesZ0Z_9 ));
    Odrv4 I__13277 (
            .O(N__63470),
            .I(\ppm_encoder_1.init_pulsesZ0Z_9 ));
    CascadeMux I__13276 (
            .O(N__63465),
            .I(N__63462));
    InMux I__13275 (
            .O(N__63462),
            .I(N__63451));
    InMux I__13274 (
            .O(N__63461),
            .I(N__63451));
    InMux I__13273 (
            .O(N__63460),
            .I(N__63442));
    InMux I__13272 (
            .O(N__63459),
            .I(N__63442));
    InMux I__13271 (
            .O(N__63458),
            .I(N__63442));
    CascadeMux I__13270 (
            .O(N__63457),
            .I(N__63435));
    CascadeMux I__13269 (
            .O(N__63456),
            .I(N__63432));
    LocalMux I__13268 (
            .O(N__63451),
            .I(N__63427));
    CascadeMux I__13267 (
            .O(N__63450),
            .I(N__63424));
    InMux I__13266 (
            .O(N__63449),
            .I(N__63419));
    LocalMux I__13265 (
            .O(N__63442),
            .I(N__63416));
    InMux I__13264 (
            .O(N__63441),
            .I(N__63407));
    InMux I__13263 (
            .O(N__63440),
            .I(N__63407));
    InMux I__13262 (
            .O(N__63439),
            .I(N__63407));
    InMux I__13261 (
            .O(N__63438),
            .I(N__63407));
    InMux I__13260 (
            .O(N__63435),
            .I(N__63400));
    InMux I__13259 (
            .O(N__63432),
            .I(N__63397));
    InMux I__13258 (
            .O(N__63431),
            .I(N__63392));
    InMux I__13257 (
            .O(N__63430),
            .I(N__63392));
    Span4Mux_h I__13256 (
            .O(N__63427),
            .I(N__63385));
    InMux I__13255 (
            .O(N__63424),
            .I(N__63382));
    InMux I__13254 (
            .O(N__63423),
            .I(N__63376));
    InMux I__13253 (
            .O(N__63422),
            .I(N__63376));
    LocalMux I__13252 (
            .O(N__63419),
            .I(N__63371));
    Span4Mux_h I__13251 (
            .O(N__63416),
            .I(N__63371));
    LocalMux I__13250 (
            .O(N__63407),
            .I(N__63368));
    InMux I__13249 (
            .O(N__63406),
            .I(N__63363));
    InMux I__13248 (
            .O(N__63405),
            .I(N__63363));
    CascadeMux I__13247 (
            .O(N__63404),
            .I(N__63360));
    CascadeMux I__13246 (
            .O(N__63403),
            .I(N__63356));
    LocalMux I__13245 (
            .O(N__63400),
            .I(N__63349));
    LocalMux I__13244 (
            .O(N__63397),
            .I(N__63349));
    LocalMux I__13243 (
            .O(N__63392),
            .I(N__63346));
    InMux I__13242 (
            .O(N__63391),
            .I(N__63341));
    InMux I__13241 (
            .O(N__63390),
            .I(N__63341));
    InMux I__13240 (
            .O(N__63389),
            .I(N__63338));
    InMux I__13239 (
            .O(N__63388),
            .I(N__63335));
    Span4Mux_v I__13238 (
            .O(N__63385),
            .I(N__63330));
    LocalMux I__13237 (
            .O(N__63382),
            .I(N__63330));
    InMux I__13236 (
            .O(N__63381),
            .I(N__63327));
    LocalMux I__13235 (
            .O(N__63376),
            .I(N__63320));
    Span4Mux_v I__13234 (
            .O(N__63371),
            .I(N__63320));
    Span4Mux_v I__13233 (
            .O(N__63368),
            .I(N__63320));
    LocalMux I__13232 (
            .O(N__63363),
            .I(N__63317));
    InMux I__13231 (
            .O(N__63360),
            .I(N__63306));
    InMux I__13230 (
            .O(N__63359),
            .I(N__63306));
    InMux I__13229 (
            .O(N__63356),
            .I(N__63306));
    InMux I__13228 (
            .O(N__63355),
            .I(N__63306));
    InMux I__13227 (
            .O(N__63354),
            .I(N__63306));
    Span4Mux_h I__13226 (
            .O(N__63349),
            .I(N__63299));
    Span4Mux_h I__13225 (
            .O(N__63346),
            .I(N__63299));
    LocalMux I__13224 (
            .O(N__63341),
            .I(N__63299));
    LocalMux I__13223 (
            .O(N__63338),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ));
    LocalMux I__13222 (
            .O(N__63335),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ));
    Odrv4 I__13221 (
            .O(N__63330),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ));
    LocalMux I__13220 (
            .O(N__63327),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ));
    Odrv4 I__13219 (
            .O(N__63320),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ));
    Odrv12 I__13218 (
            .O(N__63317),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ));
    LocalMux I__13217 (
            .O(N__63306),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ));
    Odrv4 I__13216 (
            .O(N__63299),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ));
    InMux I__13215 (
            .O(N__63282),
            .I(N__63279));
    LocalMux I__13214 (
            .O(N__63279),
            .I(N__63276));
    Span4Mux_h I__13213 (
            .O(N__63276),
            .I(N__63273));
    Odrv4 I__13212 (
            .O(N__63273),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_9 ));
    InMux I__13211 (
            .O(N__63270),
            .I(N__63267));
    LocalMux I__13210 (
            .O(N__63267),
            .I(N__63264));
    Span4Mux_v I__13209 (
            .O(N__63264),
            .I(N__63261));
    Odrv4 I__13208 (
            .O(N__63261),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_2 ));
    CascadeMux I__13207 (
            .O(N__63258),
            .I(N__63255));
    InMux I__13206 (
            .O(N__63255),
            .I(N__63252));
    LocalMux I__13205 (
            .O(N__63252),
            .I(N__63249));
    Span4Mux_h I__13204 (
            .O(N__63249),
            .I(N__63246));
    Sp12to4 I__13203 (
            .O(N__63246),
            .I(N__63243));
    Odrv12 I__13202 (
            .O(N__63243),
            .I(\ppm_encoder_1.pulses2count_9_i_0_2 ));
    InMux I__13201 (
            .O(N__63240),
            .I(N__63237));
    LocalMux I__13200 (
            .O(N__63237),
            .I(N__63232));
    CascadeMux I__13199 (
            .O(N__63236),
            .I(N__63228));
    InMux I__13198 (
            .O(N__63235),
            .I(N__63225));
    Span4Mux_v I__13197 (
            .O(N__63232),
            .I(N__63222));
    InMux I__13196 (
            .O(N__63231),
            .I(N__63217));
    InMux I__13195 (
            .O(N__63228),
            .I(N__63217));
    LocalMux I__13194 (
            .O(N__63225),
            .I(N__63214));
    Span4Mux_s0_v I__13193 (
            .O(N__63222),
            .I(N__63209));
    LocalMux I__13192 (
            .O(N__63217),
            .I(N__63209));
    Odrv4 I__13191 (
            .O(N__63214),
            .I(\ppm_encoder_1.init_pulsesZ0Z_2 ));
    Odrv4 I__13190 (
            .O(N__63209),
            .I(\ppm_encoder_1.init_pulsesZ0Z_2 ));
    CascadeMux I__13189 (
            .O(N__63204),
            .I(\pid_front.N_57_0_cascade_ ));
    CascadeMux I__13188 (
            .O(N__63201),
            .I(\pid_front.N_59_0_cascade_ ));
    InMux I__13187 (
            .O(N__63198),
            .I(N__63195));
    LocalMux I__13186 (
            .O(N__63195),
            .I(\pid_front.N_89_i ));
    CascadeMux I__13185 (
            .O(N__63192),
            .I(N__63189));
    InMux I__13184 (
            .O(N__63189),
            .I(N__63186));
    LocalMux I__13183 (
            .O(N__63186),
            .I(N__63183));
    Span4Mux_h I__13182 (
            .O(N__63183),
            .I(N__63180));
    Odrv4 I__13181 (
            .O(N__63180),
            .I(\pid_front.error_i_regZ0Z_24 ));
    InMux I__13180 (
            .O(N__63177),
            .I(N__63174));
    LocalMux I__13179 (
            .O(N__63174),
            .I(N__63171));
    Span4Mux_v I__13178 (
            .O(N__63171),
            .I(N__63168));
    Odrv4 I__13177 (
            .O(N__63168),
            .I(\pid_front.N_3 ));
    InMux I__13176 (
            .O(N__63165),
            .I(N__63162));
    LocalMux I__13175 (
            .O(N__63162),
            .I(N__63158));
    InMux I__13174 (
            .O(N__63161),
            .I(N__63155));
    Odrv4 I__13173 (
            .O(N__63158),
            .I(\pid_front.N_30_1 ));
    LocalMux I__13172 (
            .O(N__63155),
            .I(\pid_front.N_30_1 ));
    InMux I__13171 (
            .O(N__63150),
            .I(N__63145));
    CascadeMux I__13170 (
            .O(N__63149),
            .I(N__63142));
    InMux I__13169 (
            .O(N__63148),
            .I(N__63138));
    LocalMux I__13168 (
            .O(N__63145),
            .I(N__63135));
    InMux I__13167 (
            .O(N__63142),
            .I(N__63130));
    InMux I__13166 (
            .O(N__63141),
            .I(N__63130));
    LocalMux I__13165 (
            .O(N__63138),
            .I(\pid_front.N_15_0 ));
    Odrv4 I__13164 (
            .O(N__63135),
            .I(\pid_front.N_15_0 ));
    LocalMux I__13163 (
            .O(N__63130),
            .I(\pid_front.N_15_0 ));
    CascadeMux I__13162 (
            .O(N__63123),
            .I(\pid_front.N_15_0_cascade_ ));
    InMux I__13161 (
            .O(N__63120),
            .I(N__63116));
    InMux I__13160 (
            .O(N__63119),
            .I(N__63113));
    LocalMux I__13159 (
            .O(N__63116),
            .I(N__63110));
    LocalMux I__13158 (
            .O(N__63113),
            .I(\pid_front.N_57_0 ));
    Odrv4 I__13157 (
            .O(N__63110),
            .I(\pid_front.N_57_0 ));
    CascadeMux I__13156 (
            .O(N__63105),
            .I(\pid_front.m138_0_1_cascade_ ));
    InMux I__13155 (
            .O(N__63102),
            .I(N__63098));
    InMux I__13154 (
            .O(N__63101),
            .I(N__63093));
    LocalMux I__13153 (
            .O(N__63098),
            .I(N__63090));
    InMux I__13152 (
            .O(N__63097),
            .I(N__63085));
    InMux I__13151 (
            .O(N__63096),
            .I(N__63085));
    LocalMux I__13150 (
            .O(N__63093),
            .I(\pid_front.N_22_0 ));
    Odrv4 I__13149 (
            .O(N__63090),
            .I(\pid_front.N_22_0 ));
    LocalMux I__13148 (
            .O(N__63085),
            .I(\pid_front.N_22_0 ));
    InMux I__13147 (
            .O(N__63078),
            .I(N__63073));
    InMux I__13146 (
            .O(N__63077),
            .I(N__63068));
    InMux I__13145 (
            .O(N__63076),
            .I(N__63068));
    LocalMux I__13144 (
            .O(N__63073),
            .I(N__63063));
    LocalMux I__13143 (
            .O(N__63068),
            .I(N__63063));
    Span4Mux_v I__13142 (
            .O(N__63063),
            .I(N__63060));
    Odrv4 I__13141 (
            .O(N__63060),
            .I(\pid_front.m0_0_03 ));
    InMux I__13140 (
            .O(N__63057),
            .I(N__63054));
    LocalMux I__13139 (
            .O(N__63054),
            .I(\pid_front.m0_2_03 ));
    InMux I__13138 (
            .O(N__63051),
            .I(N__63048));
    LocalMux I__13137 (
            .O(N__63048),
            .I(\pid_front.m24_2_03_0 ));
    InMux I__13136 (
            .O(N__63045),
            .I(N__63042));
    LocalMux I__13135 (
            .O(N__63042),
            .I(N__63039));
    Odrv4 I__13134 (
            .O(N__63039),
            .I(\pid_front.m8_2_03_3_i_0 ));
    CascadeMux I__13133 (
            .O(N__63036),
            .I(N__63033));
    InMux I__13132 (
            .O(N__63033),
            .I(N__63030));
    LocalMux I__13131 (
            .O(N__63030),
            .I(N__63027));
    Odrv4 I__13130 (
            .O(N__63027),
            .I(\pid_front.error_i_regZ0Z_20 ));
    InMux I__13129 (
            .O(N__63024),
            .I(N__63020));
    InMux I__13128 (
            .O(N__63023),
            .I(N__63017));
    LocalMux I__13127 (
            .O(N__63020),
            .I(\pid_front.N_39_1 ));
    LocalMux I__13126 (
            .O(N__63017),
            .I(\pid_front.N_39_1 ));
    CascadeMux I__13125 (
            .O(N__63012),
            .I(\pid_front.m129_0_ns_1_cascade_ ));
    CascadeMux I__13124 (
            .O(N__63009),
            .I(N__63006));
    InMux I__13123 (
            .O(N__63006),
            .I(N__63003));
    LocalMux I__13122 (
            .O(N__63003),
            .I(N__63000));
    Odrv4 I__13121 (
            .O(N__63000),
            .I(\pid_front.m16_2_03_4 ));
    InMux I__13120 (
            .O(N__62997),
            .I(N__62993));
    InMux I__13119 (
            .O(N__62996),
            .I(N__62990));
    LocalMux I__13118 (
            .O(N__62993),
            .I(N__62987));
    LocalMux I__13117 (
            .O(N__62990),
            .I(N__62983));
    Span4Mux_v I__13116 (
            .O(N__62987),
            .I(N__62980));
    InMux I__13115 (
            .O(N__62986),
            .I(N__62977));
    Span4Mux_v I__13114 (
            .O(N__62983),
            .I(N__62973));
    Span4Mux_h I__13113 (
            .O(N__62980),
            .I(N__62970));
    LocalMux I__13112 (
            .O(N__62977),
            .I(N__62965));
    InMux I__13111 (
            .O(N__62976),
            .I(N__62962));
    Span4Mux_h I__13110 (
            .O(N__62973),
            .I(N__62959));
    Span4Mux_h I__13109 (
            .O(N__62970),
            .I(N__62956));
    InMux I__13108 (
            .O(N__62969),
            .I(N__62951));
    InMux I__13107 (
            .O(N__62968),
            .I(N__62951));
    Span4Mux_v I__13106 (
            .O(N__62965),
            .I(N__62948));
    LocalMux I__13105 (
            .O(N__62962),
            .I(N__62943));
    Span4Mux_h I__13104 (
            .O(N__62959),
            .I(N__62943));
    Span4Mux_h I__13103 (
            .O(N__62956),
            .I(N__62940));
    LocalMux I__13102 (
            .O(N__62951),
            .I(\pid_front.error_8 ));
    Odrv4 I__13101 (
            .O(N__62948),
            .I(\pid_front.error_8 ));
    Odrv4 I__13100 (
            .O(N__62943),
            .I(\pid_front.error_8 ));
    Odrv4 I__13099 (
            .O(N__62940),
            .I(\pid_front.error_8 ));
    CascadeMux I__13098 (
            .O(N__62931),
            .I(\pid_front.N_29_1_cascade_ ));
    CascadeMux I__13097 (
            .O(N__62928),
            .I(\pid_front.error_cry_3_0_c_RNI76FZ0Z08_cascade_ ));
    InMux I__13096 (
            .O(N__62925),
            .I(N__62921));
    InMux I__13095 (
            .O(N__62924),
            .I(N__62918));
    LocalMux I__13094 (
            .O(N__62921),
            .I(\pid_front.N_27_1 ));
    LocalMux I__13093 (
            .O(N__62918),
            .I(\pid_front.N_27_1 ));
    InMux I__13092 (
            .O(N__62913),
            .I(N__62910));
    LocalMux I__13091 (
            .O(N__62910),
            .I(\pid_front.error_cry_3_0_c_RNIJZ0Z5832 ));
    InMux I__13090 (
            .O(N__62907),
            .I(N__62904));
    LocalMux I__13089 (
            .O(N__62904),
            .I(\pid_front.error_cry_3_0_c_RNIJ5832Z0Z_0 ));
    InMux I__13088 (
            .O(N__62901),
            .I(N__62895));
    InMux I__13087 (
            .O(N__62900),
            .I(N__62888));
    InMux I__13086 (
            .O(N__62899),
            .I(N__62888));
    InMux I__13085 (
            .O(N__62898),
            .I(N__62888));
    LocalMux I__13084 (
            .O(N__62895),
            .I(\pid_front.N_28_1 ));
    LocalMux I__13083 (
            .O(N__62888),
            .I(\pid_front.N_28_1 ));
    InMux I__13082 (
            .O(N__62883),
            .I(N__62880));
    LocalMux I__13081 (
            .O(N__62880),
            .I(N__62876));
    CascadeMux I__13080 (
            .O(N__62879),
            .I(N__62873));
    Span4Mux_s3_v I__13079 (
            .O(N__62876),
            .I(N__62870));
    InMux I__13078 (
            .O(N__62873),
            .I(N__62867));
    Span4Mux_v I__13077 (
            .O(N__62870),
            .I(N__62862));
    LocalMux I__13076 (
            .O(N__62867),
            .I(N__62862));
    Odrv4 I__13075 (
            .O(N__62862),
            .I(\pid_front.error_i_regZ0Z_0 ));
    InMux I__13074 (
            .O(N__62859),
            .I(N__62855));
    InMux I__13073 (
            .O(N__62858),
            .I(N__62852));
    LocalMux I__13072 (
            .O(N__62855),
            .I(\pid_front.N_36_0 ));
    LocalMux I__13071 (
            .O(N__62852),
            .I(\pid_front.N_36_0 ));
    CascadeMux I__13070 (
            .O(N__62847),
            .I(\pid_front.N_63_cascade_ ));
    CascadeMux I__13069 (
            .O(N__62844),
            .I(\pid_front.m6_2_03_cascade_ ));
    InMux I__13068 (
            .O(N__62841),
            .I(N__62838));
    LocalMux I__13067 (
            .O(N__62838),
            .I(N__62835));
    Span4Mux_v I__13066 (
            .O(N__62835),
            .I(N__62832));
    Odrv4 I__13065 (
            .O(N__62832),
            .I(\pid_front.error_i_reg_9_rn_0_18 ));
    InMux I__13064 (
            .O(N__62829),
            .I(N__62824));
    InMux I__13063 (
            .O(N__62828),
            .I(N__62817));
    InMux I__13062 (
            .O(N__62827),
            .I(N__62817));
    LocalMux I__13061 (
            .O(N__62824),
            .I(N__62814));
    InMux I__13060 (
            .O(N__62823),
            .I(N__62809));
    InMux I__13059 (
            .O(N__62822),
            .I(N__62809));
    LocalMux I__13058 (
            .O(N__62817),
            .I(N__62806));
    Span4Mux_v I__13057 (
            .O(N__62814),
            .I(N__62801));
    LocalMux I__13056 (
            .O(N__62809),
            .I(N__62801));
    Span4Mux_v I__13055 (
            .O(N__62806),
            .I(N__62798));
    Span4Mux_h I__13054 (
            .O(N__62801),
            .I(N__62795));
    Odrv4 I__13053 (
            .O(N__62798),
            .I(\pid_front.m2_0_03_3_i_0 ));
    Odrv4 I__13052 (
            .O(N__62795),
            .I(\pid_front.m2_0_03_3_i_0 ));
    InMux I__13051 (
            .O(N__62790),
            .I(N__62787));
    LocalMux I__13050 (
            .O(N__62787),
            .I(N__62783));
    InMux I__13049 (
            .O(N__62786),
            .I(N__62779));
    Span4Mux_v I__13048 (
            .O(N__62783),
            .I(N__62776));
    InMux I__13047 (
            .O(N__62782),
            .I(N__62773));
    LocalMux I__13046 (
            .O(N__62779),
            .I(\pid_front.N_63 ));
    Odrv4 I__13045 (
            .O(N__62776),
            .I(\pid_front.N_63 ));
    LocalMux I__13044 (
            .O(N__62773),
            .I(\pid_front.N_63 ));
    InMux I__13043 (
            .O(N__62766),
            .I(N__62763));
    LocalMux I__13042 (
            .O(N__62763),
            .I(N__62760));
    Span4Mux_v I__13041 (
            .O(N__62760),
            .I(N__62757));
    Odrv4 I__13040 (
            .O(N__62757),
            .I(\pid_front.N_41_0 ));
    CascadeMux I__13039 (
            .O(N__62754),
            .I(\pid_front.N_41_0_cascade_ ));
    CascadeMux I__13038 (
            .O(N__62751),
            .I(\pid_side.g2_cascade_ ));
    InMux I__13037 (
            .O(N__62748),
            .I(N__62745));
    LocalMux I__13036 (
            .O(N__62745),
            .I(\pid_side.N_117_0 ));
    CascadeMux I__13035 (
            .O(N__62742),
            .I(N__62739));
    InMux I__13034 (
            .O(N__62739),
            .I(N__62736));
    LocalMux I__13033 (
            .O(N__62736),
            .I(N__62733));
    Span4Mux_v I__13032 (
            .O(N__62733),
            .I(N__62730));
    Odrv4 I__13031 (
            .O(N__62730),
            .I(\pid_front.error_i_regZ0Z_2 ));
    CascadeMux I__13030 (
            .O(N__62727),
            .I(N__62724));
    InMux I__13029 (
            .O(N__62724),
            .I(N__62721));
    LocalMux I__13028 (
            .O(N__62721),
            .I(N__62718));
    Span4Mux_v I__13027 (
            .O(N__62718),
            .I(N__62715));
    Odrv4 I__13026 (
            .O(N__62715),
            .I(\pid_front.error_i_regZ0Z_3 ));
    CascadeMux I__13025 (
            .O(N__62712),
            .I(\pid_side.m1_0_03_cascade_ ));
    InMux I__13024 (
            .O(N__62709),
            .I(N__62706));
    LocalMux I__13023 (
            .O(N__62706),
            .I(N__62703));
    Odrv4 I__13022 (
            .O(N__62703),
            .I(\pid_side.error_i_reg_esr_RNO_5Z0Z_17 ));
    InMux I__13021 (
            .O(N__62700),
            .I(N__62697));
    LocalMux I__13020 (
            .O(N__62697),
            .I(N__62694));
    Odrv4 I__13019 (
            .O(N__62694),
            .I(\pid_side.error_i_reg_esr_RNO_4Z0Z_17 ));
    CascadeMux I__13018 (
            .O(N__62691),
            .I(\pid_side.N_131_cascade_ ));
    InMux I__13017 (
            .O(N__62688),
            .I(N__62685));
    LocalMux I__13016 (
            .O(N__62685),
            .I(\pid_side.m5_2_03 ));
    CascadeMux I__13015 (
            .O(N__62682),
            .I(\pid_side.G_5_0_a5_0_1_cascade_ ));
    CascadeMux I__13014 (
            .O(N__62679),
            .I(\pid_side.N_9_cascade_ ));
    InMux I__13013 (
            .O(N__62676),
            .I(N__62673));
    LocalMux I__13012 (
            .O(N__62673),
            .I(\pid_side.G_5_0_1 ));
    InMux I__13011 (
            .O(N__62670),
            .I(N__62667));
    LocalMux I__13010 (
            .O(N__62667),
            .I(\pid_side.G_5_0_a5_2_0 ));
    InMux I__13009 (
            .O(N__62664),
            .I(N__62661));
    LocalMux I__13008 (
            .O(N__62661),
            .I(N__62658));
    Odrv4 I__13007 (
            .O(N__62658),
            .I(\pid_side.N_45_1 ));
    CascadeMux I__13006 (
            .O(N__62655),
            .I(N__62652));
    InMux I__13005 (
            .O(N__62652),
            .I(N__62649));
    LocalMux I__13004 (
            .O(N__62649),
            .I(\pid_side.m87_0_ns_1_0 ));
    IoInMux I__13003 (
            .O(N__62646),
            .I(N__62643));
    LocalMux I__13002 (
            .O(N__62643),
            .I(N__62640));
    Span4Mux_s3_v I__13001 (
            .O(N__62640),
            .I(N__62637));
    Span4Mux_v I__13000 (
            .O(N__62637),
            .I(N__62634));
    Span4Mux_v I__12999 (
            .O(N__62634),
            .I(N__62631));
    Odrv4 I__12998 (
            .O(N__62631),
            .I(GB_BUFFER_reset_system_g_THRU_CO));
    InMux I__12997 (
            .O(N__62628),
            .I(N__62625));
    LocalMux I__12996 (
            .O(N__62625),
            .I(\pid_side.N_6_0 ));
    CascadeMux I__12995 (
            .O(N__62622),
            .I(\pid_side.N_46_1_cascade_ ));
    InMux I__12994 (
            .O(N__62619),
            .I(N__62616));
    LocalMux I__12993 (
            .O(N__62616),
            .I(\pid_side.error_i_reg_esr_RNO_0Z0Z_23 ));
    InMux I__12992 (
            .O(N__62613),
            .I(N__62610));
    LocalMux I__12991 (
            .O(N__62610),
            .I(\pid_side.error_cry_9_c_RNIL6RZ0Z82 ));
    InMux I__12990 (
            .O(N__62607),
            .I(N__62604));
    LocalMux I__12989 (
            .O(N__62604),
            .I(N__62600));
    InMux I__12988 (
            .O(N__62603),
            .I(N__62597));
    Odrv12 I__12987 (
            .O(N__62600),
            .I(\pid_side.N_27_1 ));
    LocalMux I__12986 (
            .O(N__62597),
            .I(\pid_side.N_27_1 ));
    CascadeMux I__12985 (
            .O(N__62592),
            .I(\pid_side.error_cry_3_0_c_RNIJIPSZ0Z1_cascade_ ));
    InMux I__12984 (
            .O(N__62589),
            .I(N__62586));
    LocalMux I__12983 (
            .O(N__62586),
            .I(\pid_side.error_cry_3_0_c_RNIJIPS1Z0Z_0 ));
    CascadeMux I__12982 (
            .O(N__62583),
            .I(\pid_side.N_28_1_cascade_ ));
    CascadeMux I__12981 (
            .O(N__62580),
            .I(\pid_side.error_cry_0_c_RNI94FZ0Z58_cascade_ ));
    CascadeMux I__12980 (
            .O(N__62577),
            .I(\pid_side.m8_2_03_3_i_0_cascade_ ));
    InMux I__12979 (
            .O(N__62574),
            .I(N__62571));
    LocalMux I__12978 (
            .O(N__62571),
            .I(\pid_side.m24_2_03_0 ));
    InMux I__12977 (
            .O(N__62568),
            .I(N__62561));
    InMux I__12976 (
            .O(N__62567),
            .I(N__62561));
    InMux I__12975 (
            .O(N__62566),
            .I(N__62558));
    LocalMux I__12974 (
            .O(N__62561),
            .I(N__62555));
    LocalMux I__12973 (
            .O(N__62558),
            .I(N__62547));
    Span4Mux_h I__12972 (
            .O(N__62555),
            .I(N__62547));
    InMux I__12971 (
            .O(N__62554),
            .I(N__62540));
    InMux I__12970 (
            .O(N__62553),
            .I(N__62540));
    InMux I__12969 (
            .O(N__62552),
            .I(N__62540));
    Odrv4 I__12968 (
            .O(N__62547),
            .I(\pid_side.N_63 ));
    LocalMux I__12967 (
            .O(N__62540),
            .I(\pid_side.N_63 ));
    InMux I__12966 (
            .O(N__62535),
            .I(N__62529));
    InMux I__12965 (
            .O(N__62534),
            .I(N__62526));
    InMux I__12964 (
            .O(N__62533),
            .I(N__62521));
    InMux I__12963 (
            .O(N__62532),
            .I(N__62521));
    LocalMux I__12962 (
            .O(N__62529),
            .I(\pid_side.N_38_1 ));
    LocalMux I__12961 (
            .O(N__62526),
            .I(\pid_side.N_38_1 ));
    LocalMux I__12960 (
            .O(N__62521),
            .I(\pid_side.N_38_1 ));
    InMux I__12959 (
            .O(N__62514),
            .I(N__62511));
    LocalMux I__12958 (
            .O(N__62511),
            .I(N__62507));
    InMux I__12957 (
            .O(N__62510),
            .I(N__62504));
    Odrv4 I__12956 (
            .O(N__62507),
            .I(\pid_side.N_55_0 ));
    LocalMux I__12955 (
            .O(N__62504),
            .I(\pid_side.N_55_0 ));
    CascadeMux I__12954 (
            .O(N__62499),
            .I(\pid_side.N_110_cascade_ ));
    InMux I__12953 (
            .O(N__62496),
            .I(N__62492));
    InMux I__12952 (
            .O(N__62495),
            .I(N__62489));
    LocalMux I__12951 (
            .O(N__62492),
            .I(N__62486));
    LocalMux I__12950 (
            .O(N__62489),
            .I(N__62483));
    Odrv4 I__12949 (
            .O(N__62486),
            .I(\pid_side.N_3 ));
    Odrv4 I__12948 (
            .O(N__62483),
            .I(\pid_side.N_3 ));
    InMux I__12947 (
            .O(N__62478),
            .I(N__62474));
    InMux I__12946 (
            .O(N__62477),
            .I(N__62471));
    LocalMux I__12945 (
            .O(N__62474),
            .I(\pid_side.N_14_1 ));
    LocalMux I__12944 (
            .O(N__62471),
            .I(\pid_side.N_14_1 ));
    InMux I__12943 (
            .O(N__62466),
            .I(N__62463));
    LocalMux I__12942 (
            .O(N__62463),
            .I(\pid_side.N_104 ));
    CascadeMux I__12941 (
            .O(N__62460),
            .I(\pid_side.N_104_cascade_ ));
    InMux I__12940 (
            .O(N__62457),
            .I(N__62451));
    InMux I__12939 (
            .O(N__62456),
            .I(N__62446));
    InMux I__12938 (
            .O(N__62455),
            .I(N__62446));
    InMux I__12937 (
            .O(N__62454),
            .I(N__62443));
    LocalMux I__12936 (
            .O(N__62451),
            .I(\pid_side.N_49_0 ));
    LocalMux I__12935 (
            .O(N__62446),
            .I(\pid_side.N_49_0 ));
    LocalMux I__12934 (
            .O(N__62443),
            .I(\pid_side.N_49_0 ));
    CascadeMux I__12933 (
            .O(N__62436),
            .I(\pid_side.un4_error_i_reg_33_bm_1_cascade_ ));
    InMux I__12932 (
            .O(N__62433),
            .I(N__62426));
    InMux I__12931 (
            .O(N__62432),
            .I(N__62423));
    InMux I__12930 (
            .O(N__62431),
            .I(N__62420));
    InMux I__12929 (
            .O(N__62430),
            .I(N__62415));
    InMux I__12928 (
            .O(N__62429),
            .I(N__62415));
    LocalMux I__12927 (
            .O(N__62426),
            .I(\pid_side.N_39_0 ));
    LocalMux I__12926 (
            .O(N__62423),
            .I(\pid_side.N_39_0 ));
    LocalMux I__12925 (
            .O(N__62420),
            .I(\pid_side.N_39_0 ));
    LocalMux I__12924 (
            .O(N__62415),
            .I(\pid_side.N_39_0 ));
    CascadeMux I__12923 (
            .O(N__62406),
            .I(\pid_side.error_i_reg_esr_RNO_1Z0Z_23_cascade_ ));
    CascadeMux I__12922 (
            .O(N__62403),
            .I(\pid_side.error_cry_9_c_RNIL6R82Z0Z_0_cascade_ ));
    InMux I__12921 (
            .O(N__62400),
            .I(N__62396));
    InMux I__12920 (
            .O(N__62399),
            .I(N__62393));
    LocalMux I__12919 (
            .O(N__62396),
            .I(\pid_side.N_46_1 ));
    LocalMux I__12918 (
            .O(N__62393),
            .I(\pid_side.N_46_1 ));
    InMux I__12917 (
            .O(N__62388),
            .I(N__62382));
    InMux I__12916 (
            .O(N__62387),
            .I(N__62382));
    LocalMux I__12915 (
            .O(N__62382),
            .I(\pid_side.un1_pid_prereg_0_23 ));
    InMux I__12914 (
            .O(N__62379),
            .I(N__62375));
    InMux I__12913 (
            .O(N__62378),
            .I(N__62372));
    LocalMux I__12912 (
            .O(N__62375),
            .I(\pid_side.un1_pid_prereg_0_22 ));
    LocalMux I__12911 (
            .O(N__62372),
            .I(\pid_side.un1_pid_prereg_0_22 ));
    CascadeMux I__12910 (
            .O(N__62367),
            .I(\pid_side.un1_pid_prereg_0_24_cascade_ ));
    CascadeMux I__12909 (
            .O(N__62364),
            .I(\pid_side.N_11_0_cascade_ ));
    CascadeMux I__12908 (
            .O(N__62361),
            .I(\pid_side.N_15_1_cascade_ ));
    InMux I__12907 (
            .O(N__62358),
            .I(N__62355));
    LocalMux I__12906 (
            .O(N__62355),
            .I(\pid_side.m3_2_03 ));
    InMux I__12905 (
            .O(N__62352),
            .I(N__62347));
    InMux I__12904 (
            .O(N__62351),
            .I(N__62342));
    InMux I__12903 (
            .O(N__62350),
            .I(N__62342));
    LocalMux I__12902 (
            .O(N__62347),
            .I(\pid_side.N_15_1 ));
    LocalMux I__12901 (
            .O(N__62342),
            .I(\pid_side.N_15_1 ));
    CascadeMux I__12900 (
            .O(N__62337),
            .I(\pid_side.m4_2_03_cascade_ ));
    InMux I__12899 (
            .O(N__62334),
            .I(N__62331));
    LocalMux I__12898 (
            .O(N__62331),
            .I(\pid_side.N_30_1 ));
    CascadeMux I__12897 (
            .O(N__62328),
            .I(\pid_side.N_30_1_cascade_ ));
    CascadeMux I__12896 (
            .O(N__62325),
            .I(\pid_side.N_63_cascade_ ));
    InMux I__12895 (
            .O(N__62322),
            .I(N__62319));
    LocalMux I__12894 (
            .O(N__62319),
            .I(N__62314));
    InMux I__12893 (
            .O(N__62318),
            .I(N__62311));
    CascadeMux I__12892 (
            .O(N__62317),
            .I(N__62308));
    Span4Mux_h I__12891 (
            .O(N__62314),
            .I(N__62304));
    LocalMux I__12890 (
            .O(N__62311),
            .I(N__62301));
    InMux I__12889 (
            .O(N__62308),
            .I(N__62296));
    InMux I__12888 (
            .O(N__62307),
            .I(N__62296));
    Odrv4 I__12887 (
            .O(N__62304),
            .I(\pid_side.m2_0_03_3_i_0 ));
    Odrv4 I__12886 (
            .O(N__62301),
            .I(\pid_side.m2_0_03_3_i_0 ));
    LocalMux I__12885 (
            .O(N__62296),
            .I(\pid_side.m2_0_03_3_i_0 ));
    CascadeMux I__12884 (
            .O(N__62289),
            .I(\pid_side.un1_pid_prereg_0_23_cascade_ ));
    CascadeMux I__12883 (
            .O(N__62286),
            .I(\pid_side.un1_pid_prereg_0_22_cascade_ ));
    InMux I__12882 (
            .O(N__62283),
            .I(N__62278));
    InMux I__12881 (
            .O(N__62282),
            .I(N__62275));
    InMux I__12880 (
            .O(N__62281),
            .I(N__62272));
    LocalMux I__12879 (
            .O(N__62278),
            .I(\pid_side.error_i_acumm_preregZ0Z_7 ));
    LocalMux I__12878 (
            .O(N__62275),
            .I(\pid_side.error_i_acumm_preregZ0Z_7 ));
    LocalMux I__12877 (
            .O(N__62272),
            .I(\pid_side.error_i_acumm_preregZ0Z_7 ));
    InMux I__12876 (
            .O(N__62265),
            .I(N__62260));
    InMux I__12875 (
            .O(N__62264),
            .I(N__62257));
    InMux I__12874 (
            .O(N__62263),
            .I(N__62254));
    LocalMux I__12873 (
            .O(N__62260),
            .I(\pid_side.error_i_acumm_preregZ0Z_8 ));
    LocalMux I__12872 (
            .O(N__62257),
            .I(\pid_side.error_i_acumm_preregZ0Z_8 ));
    LocalMux I__12871 (
            .O(N__62254),
            .I(\pid_side.error_i_acumm_preregZ0Z_8 ));
    InMux I__12870 (
            .O(N__62247),
            .I(N__62243));
    InMux I__12869 (
            .O(N__62246),
            .I(N__62240));
    LocalMux I__12868 (
            .O(N__62243),
            .I(N__62235));
    LocalMux I__12867 (
            .O(N__62240),
            .I(N__62235));
    Span12Mux_v I__12866 (
            .O(N__62235),
            .I(N__62232));
    Odrv12 I__12865 (
            .O(N__62232),
            .I(\pid_side.error_i_acumm_preregZ0Z_0 ));
    InMux I__12864 (
            .O(N__62229),
            .I(N__62226));
    LocalMux I__12863 (
            .O(N__62226),
            .I(N__62222));
    InMux I__12862 (
            .O(N__62225),
            .I(N__62219));
    Odrv4 I__12861 (
            .O(N__62222),
            .I(\pid_side.error_p_reg_esr_RNISPTC1_0Z0Z_8 ));
    LocalMux I__12860 (
            .O(N__62219),
            .I(\pid_side.error_p_reg_esr_RNISPTC1_0Z0Z_8 ));
    InMux I__12859 (
            .O(N__62214),
            .I(N__62211));
    LocalMux I__12858 (
            .O(N__62211),
            .I(\pid_side.error_p_reg_esr_RNINKTC1Z0Z_7 ));
    InMux I__12857 (
            .O(N__62208),
            .I(N__62201));
    CascadeMux I__12856 (
            .O(N__62207),
            .I(N__62198));
    CascadeMux I__12855 (
            .O(N__62206),
            .I(N__62194));
    CascadeMux I__12854 (
            .O(N__62205),
            .I(N__62191));
    CascadeMux I__12853 (
            .O(N__62204),
            .I(N__62187));
    LocalMux I__12852 (
            .O(N__62201),
            .I(N__62182));
    InMux I__12851 (
            .O(N__62198),
            .I(N__62171));
    InMux I__12850 (
            .O(N__62197),
            .I(N__62171));
    InMux I__12849 (
            .O(N__62194),
            .I(N__62171));
    InMux I__12848 (
            .O(N__62191),
            .I(N__62171));
    InMux I__12847 (
            .O(N__62190),
            .I(N__62171));
    InMux I__12846 (
            .O(N__62187),
            .I(N__62166));
    InMux I__12845 (
            .O(N__62186),
            .I(N__62166));
    InMux I__12844 (
            .O(N__62185),
            .I(N__62163));
    Span4Mux_v I__12843 (
            .O(N__62182),
            .I(N__62160));
    LocalMux I__12842 (
            .O(N__62171),
            .I(N__62157));
    LocalMux I__12841 (
            .O(N__62166),
            .I(N__62154));
    LocalMux I__12840 (
            .O(N__62163),
            .I(\uart_drone.bit_CountZ0Z_2 ));
    Odrv4 I__12839 (
            .O(N__62160),
            .I(\uart_drone.bit_CountZ0Z_2 ));
    Odrv4 I__12838 (
            .O(N__62157),
            .I(\uart_drone.bit_CountZ0Z_2 ));
    Odrv4 I__12837 (
            .O(N__62154),
            .I(\uart_drone.bit_CountZ0Z_2 ));
    InMux I__12836 (
            .O(N__62145),
            .I(N__62142));
    LocalMux I__12835 (
            .O(N__62142),
            .I(N__62138));
    CascadeMux I__12834 (
            .O(N__62141),
            .I(N__62127));
    Span4Mux_v I__12833 (
            .O(N__62138),
            .I(N__62124));
    InMux I__12832 (
            .O(N__62137),
            .I(N__62113));
    InMux I__12831 (
            .O(N__62136),
            .I(N__62113));
    InMux I__12830 (
            .O(N__62135),
            .I(N__62113));
    InMux I__12829 (
            .O(N__62134),
            .I(N__62113));
    InMux I__12828 (
            .O(N__62133),
            .I(N__62113));
    InMux I__12827 (
            .O(N__62132),
            .I(N__62108));
    InMux I__12826 (
            .O(N__62131),
            .I(N__62108));
    InMux I__12825 (
            .O(N__62130),
            .I(N__62103));
    InMux I__12824 (
            .O(N__62127),
            .I(N__62103));
    Span4Mux_h I__12823 (
            .O(N__62124),
            .I(N__62100));
    LocalMux I__12822 (
            .O(N__62113),
            .I(N__62097));
    LocalMux I__12821 (
            .O(N__62108),
            .I(N__62094));
    LocalMux I__12820 (
            .O(N__62103),
            .I(\uart_drone.bit_CountZ0Z_1 ));
    Odrv4 I__12819 (
            .O(N__62100),
            .I(\uart_drone.bit_CountZ0Z_1 ));
    Odrv4 I__12818 (
            .O(N__62097),
            .I(\uart_drone.bit_CountZ0Z_1 ));
    Odrv12 I__12817 (
            .O(N__62094),
            .I(\uart_drone.bit_CountZ0Z_1 ));
    InMux I__12816 (
            .O(N__62085),
            .I(N__62081));
    InMux I__12815 (
            .O(N__62084),
            .I(N__62078));
    LocalMux I__12814 (
            .O(N__62081),
            .I(N__62075));
    LocalMux I__12813 (
            .O(N__62078),
            .I(N__62065));
    Span4Mux_h I__12812 (
            .O(N__62075),
            .I(N__62065));
    InMux I__12811 (
            .O(N__62074),
            .I(N__62054));
    InMux I__12810 (
            .O(N__62073),
            .I(N__62054));
    InMux I__12809 (
            .O(N__62072),
            .I(N__62054));
    InMux I__12808 (
            .O(N__62071),
            .I(N__62054));
    InMux I__12807 (
            .O(N__62070),
            .I(N__62054));
    Span4Mux_v I__12806 (
            .O(N__62065),
            .I(N__62048));
    LocalMux I__12805 (
            .O(N__62054),
            .I(N__62048));
    InMux I__12804 (
            .O(N__62053),
            .I(N__62042));
    Span4Mux_h I__12803 (
            .O(N__62048),
            .I(N__62039));
    InMux I__12802 (
            .O(N__62047),
            .I(N__62032));
    InMux I__12801 (
            .O(N__62046),
            .I(N__62032));
    InMux I__12800 (
            .O(N__62045),
            .I(N__62032));
    LocalMux I__12799 (
            .O(N__62042),
            .I(\uart_drone.bit_CountZ0Z_0 ));
    Odrv4 I__12798 (
            .O(N__62039),
            .I(\uart_drone.bit_CountZ0Z_0 ));
    LocalMux I__12797 (
            .O(N__62032),
            .I(\uart_drone.bit_CountZ0Z_0 ));
    InMux I__12796 (
            .O(N__62025),
            .I(N__62022));
    LocalMux I__12795 (
            .O(N__62022),
            .I(N__62019));
    Span4Mux_v I__12794 (
            .O(N__62019),
            .I(N__62016));
    Span4Mux_h I__12793 (
            .O(N__62016),
            .I(N__62013));
    Odrv4 I__12792 (
            .O(N__62013),
            .I(\uart_drone.data_Auxce_0_0_0 ));
    CascadeMux I__12791 (
            .O(N__62010),
            .I(\pid_side.N_15_0_cascade_ ));
    InMux I__12790 (
            .O(N__62007),
            .I(N__62002));
    InMux I__12789 (
            .O(N__62006),
            .I(N__61997));
    InMux I__12788 (
            .O(N__62005),
            .I(N__61997));
    LocalMux I__12787 (
            .O(N__62002),
            .I(\pid_side.error_i_acumm_preregZ0Z_10 ));
    LocalMux I__12786 (
            .O(N__61997),
            .I(\pid_side.error_i_acumm_preregZ0Z_10 ));
    CascadeMux I__12785 (
            .O(N__61992),
            .I(\pid_side.un10lt9_1_cascade_ ));
    InMux I__12784 (
            .O(N__61989),
            .I(N__61986));
    LocalMux I__12783 (
            .O(N__61986),
            .I(\pid_side.error_i_acumm16lt9_0 ));
    InMux I__12782 (
            .O(N__61983),
            .I(N__61980));
    LocalMux I__12781 (
            .O(N__61980),
            .I(\pid_side.un10lt9_1 ));
    CascadeMux I__12780 (
            .O(N__61977),
            .I(\pid_side.un10lt9_cascade_ ));
    InMux I__12779 (
            .O(N__61974),
            .I(N__61971));
    LocalMux I__12778 (
            .O(N__61971),
            .I(N__61968));
    Odrv4 I__12777 (
            .O(N__61968),
            .I(\pid_side.error_i_acumm_prereg_esr_RNIJ04NZ0Z_10 ));
    CascadeMux I__12776 (
            .O(N__61965),
            .I(\pid_side.un10lt11_0_cascade_ ));
    InMux I__12775 (
            .O(N__61962),
            .I(bfn_15_9_0_));
    InMux I__12774 (
            .O(N__61959),
            .I(N__61956));
    LocalMux I__12773 (
            .O(N__61956),
            .I(\pid_side.source_pid_1_sqmuxa_1_0_o2_sx ));
    InMux I__12772 (
            .O(N__61953),
            .I(N__61950));
    LocalMux I__12771 (
            .O(N__61950),
            .I(\pid_side.N_389 ));
    InMux I__12770 (
            .O(N__61947),
            .I(N__61944));
    LocalMux I__12769 (
            .O(N__61944),
            .I(\pid_side.source_pid_1_sqmuxa_1_0_a4_3 ));
    InMux I__12768 (
            .O(N__61941),
            .I(N__61938));
    LocalMux I__12767 (
            .O(N__61938),
            .I(\pid_side.un11lto30_i_a2_5_and ));
    InMux I__12766 (
            .O(N__61935),
            .I(N__61931));
    InMux I__12765 (
            .O(N__61934),
            .I(N__61928));
    LocalMux I__12764 (
            .O(N__61931),
            .I(N__61925));
    LocalMux I__12763 (
            .O(N__61928),
            .I(\pid_side.un11lto30_i_a2_6_and ));
    Odrv4 I__12762 (
            .O(N__61925),
            .I(\pid_side.un11lto30_i_a2_6_and ));
    CascadeMux I__12761 (
            .O(N__61920),
            .I(\pid_side.un11lto30_i_a2_5_and_cascade_ ));
    InMux I__12760 (
            .O(N__61917),
            .I(N__61913));
    InMux I__12759 (
            .O(N__61916),
            .I(N__61910));
    LocalMux I__12758 (
            .O(N__61913),
            .I(N__61907));
    LocalMux I__12757 (
            .O(N__61910),
            .I(N__61904));
    Span4Mux_v I__12756 (
            .O(N__61907),
            .I(N__61901));
    Span4Mux_h I__12755 (
            .O(N__61904),
            .I(N__61898));
    Odrv4 I__12754 (
            .O(N__61901),
            .I(\pid_side.un11lto30_i_a2_4_and ));
    Odrv4 I__12753 (
            .O(N__61898),
            .I(\pid_side.un11lto30_i_a2_4_and ));
    InMux I__12752 (
            .O(N__61893),
            .I(N__61884));
    InMux I__12751 (
            .O(N__61892),
            .I(N__61884));
    InMux I__12750 (
            .O(N__61891),
            .I(N__61879));
    InMux I__12749 (
            .O(N__61890),
            .I(N__61879));
    InMux I__12748 (
            .O(N__61889),
            .I(N__61876));
    LocalMux I__12747 (
            .O(N__61884),
            .I(\pid_side.N_98 ));
    LocalMux I__12746 (
            .O(N__61879),
            .I(\pid_side.N_98 ));
    LocalMux I__12745 (
            .O(N__61876),
            .I(\pid_side.N_98 ));
    InMux I__12744 (
            .O(N__61869),
            .I(N__61866));
    LocalMux I__12743 (
            .O(N__61866),
            .I(N__61863));
    Span4Mux_h I__12742 (
            .O(N__61863),
            .I(N__61860));
    Span4Mux_h I__12741 (
            .O(N__61860),
            .I(N__61857));
    Odrv4 I__12740 (
            .O(N__61857),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_2Z0Z_9 ));
    InMux I__12739 (
            .O(N__61854),
            .I(N__61841));
    InMux I__12738 (
            .O(N__61853),
            .I(N__61841));
    InMux I__12737 (
            .O(N__61852),
            .I(N__61841));
    CascadeMux I__12736 (
            .O(N__61851),
            .I(N__61837));
    InMux I__12735 (
            .O(N__61850),
            .I(N__61829));
    InMux I__12734 (
            .O(N__61849),
            .I(N__61829));
    InMux I__12733 (
            .O(N__61848),
            .I(N__61829));
    LocalMux I__12732 (
            .O(N__61841),
            .I(N__61826));
    InMux I__12731 (
            .O(N__61840),
            .I(N__61823));
    InMux I__12730 (
            .O(N__61837),
            .I(N__61818));
    InMux I__12729 (
            .O(N__61836),
            .I(N__61818));
    LocalMux I__12728 (
            .O(N__61829),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_3_rep2_RNIAZ0Z6041 ));
    Odrv12 I__12727 (
            .O(N__61826),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_3_rep2_RNIAZ0Z6041 ));
    LocalMux I__12726 (
            .O(N__61823),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_3_rep2_RNIAZ0Z6041 ));
    LocalMux I__12725 (
            .O(N__61818),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_3_rep2_RNIAZ0Z6041 ));
    InMux I__12724 (
            .O(N__61809),
            .I(N__61805));
    CascadeMux I__12723 (
            .O(N__61808),
            .I(N__61802));
    LocalMux I__12722 (
            .O(N__61805),
            .I(N__61799));
    InMux I__12721 (
            .O(N__61802),
            .I(N__61796));
    Span4Mux_v I__12720 (
            .O(N__61799),
            .I(N__61790));
    LocalMux I__12719 (
            .O(N__61796),
            .I(N__61790));
    InMux I__12718 (
            .O(N__61795),
            .I(N__61787));
    Span4Mux_h I__12717 (
            .O(N__61790),
            .I(N__61784));
    LocalMux I__12716 (
            .O(N__61787),
            .I(\ppm_encoder_1.rudderZ0Z_9 ));
    Odrv4 I__12715 (
            .O(N__61784),
            .I(\ppm_encoder_1.rudderZ0Z_9 ));
    InMux I__12714 (
            .O(N__61779),
            .I(N__61776));
    LocalMux I__12713 (
            .O(N__61776),
            .I(N__61773));
    Odrv4 I__12712 (
            .O(N__61773),
            .I(\ppm_encoder_1.pulses2count_9_i_2_9 ));
    CascadeMux I__12711 (
            .O(N__61770),
            .I(N__61767));
    InMux I__12710 (
            .O(N__61767),
            .I(N__61763));
    InMux I__12709 (
            .O(N__61766),
            .I(N__61759));
    LocalMux I__12708 (
            .O(N__61763),
            .I(N__61756));
    CascadeMux I__12707 (
            .O(N__61762),
            .I(N__61753));
    LocalMux I__12706 (
            .O(N__61759),
            .I(N__61750));
    Span4Mux_h I__12705 (
            .O(N__61756),
            .I(N__61747));
    InMux I__12704 (
            .O(N__61753),
            .I(N__61744));
    Span12Mux_s9_v I__12703 (
            .O(N__61750),
            .I(N__61741));
    Span4Mux_v I__12702 (
            .O(N__61747),
            .I(N__61738));
    LocalMux I__12701 (
            .O(N__61744),
            .I(\ppm_encoder_1.throttleZ0Z_6 ));
    Odrv12 I__12700 (
            .O(N__61741),
            .I(\ppm_encoder_1.throttleZ0Z_6 ));
    Odrv4 I__12699 (
            .O(N__61738),
            .I(\ppm_encoder_1.throttleZ0Z_6 ));
    InMux I__12698 (
            .O(N__61731),
            .I(N__61727));
    InMux I__12697 (
            .O(N__61730),
            .I(N__61724));
    LocalMux I__12696 (
            .O(N__61727),
            .I(N__61720));
    LocalMux I__12695 (
            .O(N__61724),
            .I(N__61717));
    InMux I__12694 (
            .O(N__61723),
            .I(N__61714));
    Span4Mux_h I__12693 (
            .O(N__61720),
            .I(N__61711));
    Span4Mux_v I__12692 (
            .O(N__61717),
            .I(N__61708));
    LocalMux I__12691 (
            .O(N__61714),
            .I(\ppm_encoder_1.aileronZ0Z_6 ));
    Odrv4 I__12690 (
            .O(N__61711),
            .I(\ppm_encoder_1.aileronZ0Z_6 ));
    Odrv4 I__12689 (
            .O(N__61708),
            .I(\ppm_encoder_1.aileronZ0Z_6 ));
    InMux I__12688 (
            .O(N__61701),
            .I(N__61698));
    LocalMux I__12687 (
            .O(N__61698),
            .I(\ppm_encoder_1.pulses2count_9_0_0_6 ));
    InMux I__12686 (
            .O(N__61695),
            .I(N__61691));
    CascadeMux I__12685 (
            .O(N__61694),
            .I(N__61686));
    LocalMux I__12684 (
            .O(N__61691),
            .I(N__61683));
    CascadeMux I__12683 (
            .O(N__61690),
            .I(N__61680));
    InMux I__12682 (
            .O(N__61689),
            .I(N__61675));
    InMux I__12681 (
            .O(N__61686),
            .I(N__61675));
    Span4Mux_v I__12680 (
            .O(N__61683),
            .I(N__61672));
    InMux I__12679 (
            .O(N__61680),
            .I(N__61669));
    LocalMux I__12678 (
            .O(N__61675),
            .I(N__61666));
    Span4Mux_h I__12677 (
            .O(N__61672),
            .I(N__61663));
    LocalMux I__12676 (
            .O(N__61669),
            .I(N__61660));
    Span4Mux_h I__12675 (
            .O(N__61666),
            .I(N__61657));
    Odrv4 I__12674 (
            .O(N__61663),
            .I(\ppm_encoder_1.init_pulsesZ0Z_6 ));
    Odrv4 I__12673 (
            .O(N__61660),
            .I(\ppm_encoder_1.init_pulsesZ0Z_6 ));
    Odrv4 I__12672 (
            .O(N__61657),
            .I(\ppm_encoder_1.init_pulsesZ0Z_6 ));
    CascadeMux I__12671 (
            .O(N__61650),
            .I(N__61647));
    InMux I__12670 (
            .O(N__61647),
            .I(N__61644));
    LocalMux I__12669 (
            .O(N__61644),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_2Z0Z_6 ));
    CascadeMux I__12668 (
            .O(N__61641),
            .I(N__61634));
    InMux I__12667 (
            .O(N__61640),
            .I(N__61620));
    InMux I__12666 (
            .O(N__61639),
            .I(N__61620));
    InMux I__12665 (
            .O(N__61638),
            .I(N__61615));
    InMux I__12664 (
            .O(N__61637),
            .I(N__61612));
    InMux I__12663 (
            .O(N__61634),
            .I(N__61605));
    InMux I__12662 (
            .O(N__61633),
            .I(N__61605));
    InMux I__12661 (
            .O(N__61632),
            .I(N__61605));
    InMux I__12660 (
            .O(N__61631),
            .I(N__61601));
    InMux I__12659 (
            .O(N__61630),
            .I(N__61596));
    InMux I__12658 (
            .O(N__61629),
            .I(N__61596));
    CascadeMux I__12657 (
            .O(N__61628),
            .I(N__61593));
    InMux I__12656 (
            .O(N__61627),
            .I(N__61590));
    InMux I__12655 (
            .O(N__61626),
            .I(N__61585));
    InMux I__12654 (
            .O(N__61625),
            .I(N__61585));
    LocalMux I__12653 (
            .O(N__61620),
            .I(N__61582));
    InMux I__12652 (
            .O(N__61619),
            .I(N__61575));
    InMux I__12651 (
            .O(N__61618),
            .I(N__61575));
    LocalMux I__12650 (
            .O(N__61615),
            .I(N__61572));
    LocalMux I__12649 (
            .O(N__61612),
            .I(N__61567));
    LocalMux I__12648 (
            .O(N__61605),
            .I(N__61567));
    InMux I__12647 (
            .O(N__61604),
            .I(N__61562));
    LocalMux I__12646 (
            .O(N__61601),
            .I(N__61559));
    LocalMux I__12645 (
            .O(N__61596),
            .I(N__61556));
    InMux I__12644 (
            .O(N__61593),
            .I(N__61553));
    LocalMux I__12643 (
            .O(N__61590),
            .I(N__61550));
    LocalMux I__12642 (
            .O(N__61585),
            .I(N__61547));
    Span4Mux_v I__12641 (
            .O(N__61582),
            .I(N__61544));
    InMux I__12640 (
            .O(N__61581),
            .I(N__61539));
    InMux I__12639 (
            .O(N__61580),
            .I(N__61539));
    LocalMux I__12638 (
            .O(N__61575),
            .I(N__61536));
    Span4Mux_v I__12637 (
            .O(N__61572),
            .I(N__61531));
    Span4Mux_v I__12636 (
            .O(N__61567),
            .I(N__61531));
    InMux I__12635 (
            .O(N__61566),
            .I(N__61528));
    InMux I__12634 (
            .O(N__61565),
            .I(N__61525));
    LocalMux I__12633 (
            .O(N__61562),
            .I(N__61518));
    Span4Mux_s3_v I__12632 (
            .O(N__61559),
            .I(N__61518));
    Span4Mux_h I__12631 (
            .O(N__61556),
            .I(N__61518));
    LocalMux I__12630 (
            .O(N__61553),
            .I(N__61509));
    Span4Mux_v I__12629 (
            .O(N__61550),
            .I(N__61509));
    Span4Mux_v I__12628 (
            .O(N__61547),
            .I(N__61509));
    Span4Mux_h I__12627 (
            .O(N__61544),
            .I(N__61509));
    LocalMux I__12626 (
            .O(N__61539),
            .I(N__61504));
    Span4Mux_v I__12625 (
            .O(N__61536),
            .I(N__61504));
    Span4Mux_h I__12624 (
            .O(N__61531),
            .I(N__61501));
    LocalMux I__12623 (
            .O(N__61528),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_0 ));
    LocalMux I__12622 (
            .O(N__61525),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_0 ));
    Odrv4 I__12621 (
            .O(N__61518),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_0 ));
    Odrv4 I__12620 (
            .O(N__61509),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_0 ));
    Odrv4 I__12619 (
            .O(N__61504),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_0 ));
    Odrv4 I__12618 (
            .O(N__61501),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_0 ));
    InMux I__12617 (
            .O(N__61488),
            .I(N__61483));
    CascadeMux I__12616 (
            .O(N__61487),
            .I(N__61480));
    CascadeMux I__12615 (
            .O(N__61486),
            .I(N__61477));
    LocalMux I__12614 (
            .O(N__61483),
            .I(N__61474));
    InMux I__12613 (
            .O(N__61480),
            .I(N__61471));
    InMux I__12612 (
            .O(N__61477),
            .I(N__61468));
    Span4Mux_h I__12611 (
            .O(N__61474),
            .I(N__61463));
    LocalMux I__12610 (
            .O(N__61471),
            .I(N__61463));
    LocalMux I__12609 (
            .O(N__61468),
            .I(\ppm_encoder_1.throttleZ0Z_13 ));
    Odrv4 I__12608 (
            .O(N__61463),
            .I(\ppm_encoder_1.throttleZ0Z_13 ));
    InMux I__12607 (
            .O(N__61458),
            .I(N__61453));
    CascadeMux I__12606 (
            .O(N__61457),
            .I(N__61444));
    CascadeMux I__12605 (
            .O(N__61456),
            .I(N__61440));
    LocalMux I__12604 (
            .O(N__61453),
            .I(N__61437));
    CascadeMux I__12603 (
            .O(N__61452),
            .I(N__61434));
    CascadeMux I__12602 (
            .O(N__61451),
            .I(N__61431));
    CascadeMux I__12601 (
            .O(N__61450),
            .I(N__61427));
    CascadeMux I__12600 (
            .O(N__61449),
            .I(N__61424));
    CascadeMux I__12599 (
            .O(N__61448),
            .I(N__61421));
    CascadeMux I__12598 (
            .O(N__61447),
            .I(N__61414));
    InMux I__12597 (
            .O(N__61444),
            .I(N__61407));
    InMux I__12596 (
            .O(N__61443),
            .I(N__61407));
    InMux I__12595 (
            .O(N__61440),
            .I(N__61407));
    Span4Mux_v I__12594 (
            .O(N__61437),
            .I(N__61404));
    InMux I__12593 (
            .O(N__61434),
            .I(N__61397));
    InMux I__12592 (
            .O(N__61431),
            .I(N__61397));
    InMux I__12591 (
            .O(N__61430),
            .I(N__61397));
    InMux I__12590 (
            .O(N__61427),
            .I(N__61389));
    InMux I__12589 (
            .O(N__61424),
            .I(N__61389));
    InMux I__12588 (
            .O(N__61421),
            .I(N__61384));
    InMux I__12587 (
            .O(N__61420),
            .I(N__61384));
    InMux I__12586 (
            .O(N__61419),
            .I(N__61379));
    InMux I__12585 (
            .O(N__61418),
            .I(N__61379));
    InMux I__12584 (
            .O(N__61417),
            .I(N__61376));
    InMux I__12583 (
            .O(N__61414),
            .I(N__61373));
    LocalMux I__12582 (
            .O(N__61407),
            .I(N__61370));
    Span4Mux_h I__12581 (
            .O(N__61404),
            .I(N__61365));
    LocalMux I__12580 (
            .O(N__61397),
            .I(N__61365));
    CascadeMux I__12579 (
            .O(N__61396),
            .I(N__61362));
    InMux I__12578 (
            .O(N__61395),
            .I(N__61357));
    InMux I__12577 (
            .O(N__61394),
            .I(N__61357));
    LocalMux I__12576 (
            .O(N__61389),
            .I(N__61352));
    LocalMux I__12575 (
            .O(N__61384),
            .I(N__61352));
    LocalMux I__12574 (
            .O(N__61379),
            .I(N__61349));
    LocalMux I__12573 (
            .O(N__61376),
            .I(N__61346));
    LocalMux I__12572 (
            .O(N__61373),
            .I(N__61341));
    Span4Mux_v I__12571 (
            .O(N__61370),
            .I(N__61341));
    Span4Mux_v I__12570 (
            .O(N__61365),
            .I(N__61338));
    InMux I__12569 (
            .O(N__61362),
            .I(N__61335));
    LocalMux I__12568 (
            .O(N__61357),
            .I(N__61332));
    Span4Mux_v I__12567 (
            .O(N__61352),
            .I(N__61329));
    Span4Mux_v I__12566 (
            .O(N__61349),
            .I(N__61326));
    Span4Mux_s2_v I__12565 (
            .O(N__61346),
            .I(N__61319));
    Span4Mux_s2_v I__12564 (
            .O(N__61341),
            .I(N__61319));
    Span4Mux_s2_v I__12563 (
            .O(N__61338),
            .I(N__61319));
    LocalMux I__12562 (
            .O(N__61335),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_1 ));
    Odrv12 I__12561 (
            .O(N__61332),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_1 ));
    Odrv4 I__12560 (
            .O(N__61329),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_1 ));
    Odrv4 I__12559 (
            .O(N__61326),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_1 ));
    Odrv4 I__12558 (
            .O(N__61319),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_1 ));
    InMux I__12557 (
            .O(N__61308),
            .I(N__61304));
    CascadeMux I__12556 (
            .O(N__61307),
            .I(N__61300));
    LocalMux I__12555 (
            .O(N__61304),
            .I(N__61297));
    InMux I__12554 (
            .O(N__61303),
            .I(N__61294));
    InMux I__12553 (
            .O(N__61300),
            .I(N__61291));
    Span4Mux_h I__12552 (
            .O(N__61297),
            .I(N__61286));
    LocalMux I__12551 (
            .O(N__61294),
            .I(N__61286));
    LocalMux I__12550 (
            .O(N__61291),
            .I(\ppm_encoder_1.aileronZ0Z_13 ));
    Odrv4 I__12549 (
            .O(N__61286),
            .I(\ppm_encoder_1.aileronZ0Z_13 ));
    InMux I__12548 (
            .O(N__61281),
            .I(N__61278));
    LocalMux I__12547 (
            .O(N__61278),
            .I(\ppm_encoder_1.pulses2count_9_0_0_13 ));
    InMux I__12546 (
            .O(N__61275),
            .I(N__61272));
    LocalMux I__12545 (
            .O(N__61272),
            .I(\pid_side.source_pid10lt4_0 ));
    InMux I__12544 (
            .O(N__61269),
            .I(N__61266));
    LocalMux I__12543 (
            .O(N__61266),
            .I(\pid_side.un11lto30_i_a2_0_and ));
    InMux I__12542 (
            .O(N__61263),
            .I(N__61260));
    LocalMux I__12541 (
            .O(N__61260),
            .I(N__61257));
    Span4Mux_h I__12540 (
            .O(N__61257),
            .I(N__61254));
    Odrv4 I__12539 (
            .O(N__61254),
            .I(\pid_side.N_11_i ));
    InMux I__12538 (
            .O(N__61251),
            .I(N__61248));
    LocalMux I__12537 (
            .O(N__61248),
            .I(N__61245));
    Odrv4 I__12536 (
            .O(N__61245),
            .I(\pid_side.un11lto30_i_a2_2_and ));
    CascadeMux I__12535 (
            .O(N__61242),
            .I(N__61239));
    InMux I__12534 (
            .O(N__61239),
            .I(N__61233));
    InMux I__12533 (
            .O(N__61238),
            .I(N__61233));
    LocalMux I__12532 (
            .O(N__61233),
            .I(N__61230));
    Span4Mux_h I__12531 (
            .O(N__61230),
            .I(N__61227));
    Span4Mux_v I__12530 (
            .O(N__61227),
            .I(N__61224));
    Odrv4 I__12529 (
            .O(N__61224),
            .I(\ppm_encoder_1.N_486_9 ));
    CascadeMux I__12528 (
            .O(N__61221),
            .I(\ppm_encoder_1.N_486_18_cascade_ ));
    InMux I__12527 (
            .O(N__61218),
            .I(N__61214));
    InMux I__12526 (
            .O(N__61217),
            .I(N__61211));
    LocalMux I__12525 (
            .O(N__61214),
            .I(N__61208));
    LocalMux I__12524 (
            .O(N__61211),
            .I(N__61205));
    Span4Mux_v I__12523 (
            .O(N__61208),
            .I(N__61199));
    Span4Mux_h I__12522 (
            .O(N__61205),
            .I(N__61196));
    InMux I__12521 (
            .O(N__61204),
            .I(N__61193));
    InMux I__12520 (
            .O(N__61203),
            .I(N__61188));
    InMux I__12519 (
            .O(N__61202),
            .I(N__61188));
    Odrv4 I__12518 (
            .O(N__61199),
            .I(\ppm_encoder_1.PPM_STATEZ0Z_1 ));
    Odrv4 I__12517 (
            .O(N__61196),
            .I(\ppm_encoder_1.PPM_STATEZ0Z_1 ));
    LocalMux I__12516 (
            .O(N__61193),
            .I(\ppm_encoder_1.PPM_STATEZ0Z_1 ));
    LocalMux I__12515 (
            .O(N__61188),
            .I(\ppm_encoder_1.PPM_STATEZ0Z_1 ));
    InMux I__12514 (
            .O(N__61179),
            .I(N__61173));
    InMux I__12513 (
            .O(N__61178),
            .I(N__61173));
    LocalMux I__12512 (
            .O(N__61173),
            .I(N__61170));
    Span4Mux_h I__12511 (
            .O(N__61170),
            .I(N__61167));
    Odrv4 I__12510 (
            .O(N__61167),
            .I(\ppm_encoder_1.counter_RNI09RH2Z0Z_18 ));
    InMux I__12509 (
            .O(N__61164),
            .I(N__61156));
    InMux I__12508 (
            .O(N__61163),
            .I(N__61156));
    InMux I__12507 (
            .O(N__61162),
            .I(N__61153));
    InMux I__12506 (
            .O(N__61161),
            .I(N__61150));
    LocalMux I__12505 (
            .O(N__61156),
            .I(N__61147));
    LocalMux I__12504 (
            .O(N__61153),
            .I(N__61144));
    LocalMux I__12503 (
            .O(N__61150),
            .I(N__61141));
    Span4Mux_h I__12502 (
            .O(N__61147),
            .I(N__61138));
    Span4Mux_h I__12501 (
            .O(N__61144),
            .I(N__61130));
    Span4Mux_h I__12500 (
            .O(N__61141),
            .I(N__61130));
    Span4Mux_h I__12499 (
            .O(N__61138),
            .I(N__61127));
    InMux I__12498 (
            .O(N__61137),
            .I(N__61124));
    InMux I__12497 (
            .O(N__61136),
            .I(N__61119));
    InMux I__12496 (
            .O(N__61135),
            .I(N__61119));
    Odrv4 I__12495 (
            .O(N__61130),
            .I(\ppm_encoder_1.PPM_STATEZ0Z_0 ));
    Odrv4 I__12494 (
            .O(N__61127),
            .I(\ppm_encoder_1.PPM_STATEZ0Z_0 ));
    LocalMux I__12493 (
            .O(N__61124),
            .I(\ppm_encoder_1.PPM_STATEZ0Z_0 ));
    LocalMux I__12492 (
            .O(N__61119),
            .I(\ppm_encoder_1.PPM_STATEZ0Z_0 ));
    InMux I__12491 (
            .O(N__61110),
            .I(N__61106));
    InMux I__12490 (
            .O(N__61109),
            .I(N__61102));
    LocalMux I__12489 (
            .O(N__61106),
            .I(N__61099));
    InMux I__12488 (
            .O(N__61105),
            .I(N__61096));
    LocalMux I__12487 (
            .O(N__61102),
            .I(N__61093));
    Span4Mux_v I__12486 (
            .O(N__61099),
            .I(N__61086));
    LocalMux I__12485 (
            .O(N__61096),
            .I(N__61086));
    Span4Mux_v I__12484 (
            .O(N__61093),
            .I(N__61086));
    Odrv4 I__12483 (
            .O(N__61086),
            .I(\ppm_encoder_1.counter24_0_N_2_THRU_CO ));
    CascadeMux I__12482 (
            .O(N__61083),
            .I(\ppm_encoder_1.counter_RNI09RH2Z0Z_18_cascade_ ));
    InMux I__12481 (
            .O(N__61080),
            .I(N__61077));
    LocalMux I__12480 (
            .O(N__61077),
            .I(N__61074));
    Span4Mux_h I__12479 (
            .O(N__61074),
            .I(N__61071));
    Span4Mux_s2_v I__12478 (
            .O(N__61071),
            .I(N__61068));
    Odrv4 I__12477 (
            .O(N__61068),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_17 ));
    CascadeMux I__12476 (
            .O(N__61065),
            .I(N__61061));
    CascadeMux I__12475 (
            .O(N__61064),
            .I(N__61058));
    InMux I__12474 (
            .O(N__61061),
            .I(N__61047));
    InMux I__12473 (
            .O(N__61058),
            .I(N__61047));
    CascadeMux I__12472 (
            .O(N__61057),
            .I(N__61044));
    InMux I__12471 (
            .O(N__61056),
            .I(N__61034));
    InMux I__12470 (
            .O(N__61055),
            .I(N__61034));
    InMux I__12469 (
            .O(N__61054),
            .I(N__61034));
    InMux I__12468 (
            .O(N__61053),
            .I(N__61029));
    InMux I__12467 (
            .O(N__61052),
            .I(N__61029));
    LocalMux I__12466 (
            .O(N__61047),
            .I(N__61026));
    InMux I__12465 (
            .O(N__61044),
            .I(N__61023));
    CascadeMux I__12464 (
            .O(N__61043),
            .I(N__61020));
    CascadeMux I__12463 (
            .O(N__61042),
            .I(N__61016));
    InMux I__12462 (
            .O(N__61041),
            .I(N__61011));
    LocalMux I__12461 (
            .O(N__61034),
            .I(N__61008));
    LocalMux I__12460 (
            .O(N__61029),
            .I(N__61001));
    Span4Mux_h I__12459 (
            .O(N__61026),
            .I(N__61001));
    LocalMux I__12458 (
            .O(N__61023),
            .I(N__61001));
    InMux I__12457 (
            .O(N__61020),
            .I(N__60996));
    InMux I__12456 (
            .O(N__61019),
            .I(N__60996));
    InMux I__12455 (
            .O(N__61016),
            .I(N__60991));
    InMux I__12454 (
            .O(N__61015),
            .I(N__60991));
    InMux I__12453 (
            .O(N__61014),
            .I(N__60988));
    LocalMux I__12452 (
            .O(N__61011),
            .I(N__60978));
    Span4Mux_v I__12451 (
            .O(N__61008),
            .I(N__60978));
    Span4Mux_v I__12450 (
            .O(N__61001),
            .I(N__60978));
    LocalMux I__12449 (
            .O(N__60996),
            .I(N__60975));
    LocalMux I__12448 (
            .O(N__60991),
            .I(N__60972));
    LocalMux I__12447 (
            .O(N__60988),
            .I(N__60969));
    InMux I__12446 (
            .O(N__60987),
            .I(N__60964));
    InMux I__12445 (
            .O(N__60986),
            .I(N__60964));
    InMux I__12444 (
            .O(N__60985),
            .I(N__60961));
    Span4Mux_h I__12443 (
            .O(N__60978),
            .I(N__60958));
    Span12Mux_s0_v I__12442 (
            .O(N__60975),
            .I(N__60953));
    Span12Mux_h I__12441 (
            .O(N__60972),
            .I(N__60953));
    Odrv12 I__12440 (
            .O(N__60969),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_3_repZ0Z2 ));
    LocalMux I__12439 (
            .O(N__60964),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_3_repZ0Z2 ));
    LocalMux I__12438 (
            .O(N__60961),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_3_repZ0Z2 ));
    Odrv4 I__12437 (
            .O(N__60958),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_3_repZ0Z2 ));
    Odrv12 I__12436 (
            .O(N__60953),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_3_repZ0Z2 ));
    CascadeMux I__12435 (
            .O(N__60942),
            .I(N__60935));
    InMux I__12434 (
            .O(N__60941),
            .I(N__60926));
    InMux I__12433 (
            .O(N__60940),
            .I(N__60926));
    InMux I__12432 (
            .O(N__60939),
            .I(N__60918));
    InMux I__12431 (
            .O(N__60938),
            .I(N__60918));
    InMux I__12430 (
            .O(N__60935),
            .I(N__60909));
    InMux I__12429 (
            .O(N__60934),
            .I(N__60909));
    InMux I__12428 (
            .O(N__60933),
            .I(N__60909));
    InMux I__12427 (
            .O(N__60932),
            .I(N__60909));
    InMux I__12426 (
            .O(N__60931),
            .I(N__60901));
    LocalMux I__12425 (
            .O(N__60926),
            .I(N__60898));
    InMux I__12424 (
            .O(N__60925),
            .I(N__60894));
    InMux I__12423 (
            .O(N__60924),
            .I(N__60891));
    InMux I__12422 (
            .O(N__60923),
            .I(N__60888));
    LocalMux I__12421 (
            .O(N__60918),
            .I(N__60885));
    LocalMux I__12420 (
            .O(N__60909),
            .I(N__60882));
    InMux I__12419 (
            .O(N__60908),
            .I(N__60876));
    InMux I__12418 (
            .O(N__60907),
            .I(N__60869));
    InMux I__12417 (
            .O(N__60906),
            .I(N__60869));
    InMux I__12416 (
            .O(N__60905),
            .I(N__60869));
    InMux I__12415 (
            .O(N__60904),
            .I(N__60866));
    LocalMux I__12414 (
            .O(N__60901),
            .I(N__60861));
    Span4Mux_s1_v I__12413 (
            .O(N__60898),
            .I(N__60861));
    InMux I__12412 (
            .O(N__60897),
            .I(N__60856));
    LocalMux I__12411 (
            .O(N__60894),
            .I(N__60853));
    LocalMux I__12410 (
            .O(N__60891),
            .I(N__60848));
    LocalMux I__12409 (
            .O(N__60888),
            .I(N__60848));
    Span4Mux_s2_v I__12408 (
            .O(N__60885),
            .I(N__60843));
    Span4Mux_h I__12407 (
            .O(N__60882),
            .I(N__60843));
    InMux I__12406 (
            .O(N__60881),
            .I(N__60836));
    InMux I__12405 (
            .O(N__60880),
            .I(N__60836));
    InMux I__12404 (
            .O(N__60879),
            .I(N__60836));
    LocalMux I__12403 (
            .O(N__60876),
            .I(N__60833));
    LocalMux I__12402 (
            .O(N__60869),
            .I(N__60830));
    LocalMux I__12401 (
            .O(N__60866),
            .I(N__60825));
    Span4Mux_v I__12400 (
            .O(N__60861),
            .I(N__60825));
    InMux I__12399 (
            .O(N__60860),
            .I(N__60820));
    InMux I__12398 (
            .O(N__60859),
            .I(N__60820));
    LocalMux I__12397 (
            .O(N__60856),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z2 ));
    Odrv4 I__12396 (
            .O(N__60853),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z2 ));
    Odrv4 I__12395 (
            .O(N__60848),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z2 ));
    Odrv4 I__12394 (
            .O(N__60843),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z2 ));
    LocalMux I__12393 (
            .O(N__60836),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z2 ));
    Odrv4 I__12392 (
            .O(N__60833),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z2 ));
    Odrv12 I__12391 (
            .O(N__60830),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z2 ));
    Odrv4 I__12390 (
            .O(N__60825),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z2 ));
    LocalMux I__12389 (
            .O(N__60820),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z2 ));
    CascadeMux I__12388 (
            .O(N__60801),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_3_rep2_RNIAZ0Z6041_cascade_ ));
    CascadeMux I__12387 (
            .O(N__60798),
            .I(N__60795));
    InMux I__12386 (
            .O(N__60795),
            .I(N__60791));
    InMux I__12385 (
            .O(N__60794),
            .I(N__60787));
    LocalMux I__12384 (
            .O(N__60791),
            .I(N__60784));
    InMux I__12383 (
            .O(N__60790),
            .I(N__60781));
    LocalMux I__12382 (
            .O(N__60787),
            .I(N__60778));
    Span4Mux_h I__12381 (
            .O(N__60784),
            .I(N__60775));
    LocalMux I__12380 (
            .O(N__60781),
            .I(\ppm_encoder_1.rudderZ0Z_10 ));
    Odrv12 I__12379 (
            .O(N__60778),
            .I(\ppm_encoder_1.rudderZ0Z_10 ));
    Odrv4 I__12378 (
            .O(N__60775),
            .I(\ppm_encoder_1.rudderZ0Z_10 ));
    InMux I__12377 (
            .O(N__60768),
            .I(N__60765));
    LocalMux I__12376 (
            .O(N__60765),
            .I(N__60762));
    Odrv4 I__12375 (
            .O(N__60762),
            .I(\ppm_encoder_1.pulses2count_9_i_0_2_10 ));
    InMux I__12374 (
            .O(N__60759),
            .I(N__60754));
    InMux I__12373 (
            .O(N__60758),
            .I(N__60751));
    CascadeMux I__12372 (
            .O(N__60757),
            .I(N__60748));
    LocalMux I__12371 (
            .O(N__60754),
            .I(N__60745));
    LocalMux I__12370 (
            .O(N__60751),
            .I(N__60742));
    InMux I__12369 (
            .O(N__60748),
            .I(N__60739));
    Span4Mux_v I__12368 (
            .O(N__60745),
            .I(N__60736));
    Span12Mux_s6_v I__12367 (
            .O(N__60742),
            .I(N__60733));
    LocalMux I__12366 (
            .O(N__60739),
            .I(N__60728));
    Span4Mux_h I__12365 (
            .O(N__60736),
            .I(N__60728));
    Odrv12 I__12364 (
            .O(N__60733),
            .I(\ppm_encoder_1.throttleZ0Z_10 ));
    Odrv4 I__12363 (
            .O(N__60728),
            .I(\ppm_encoder_1.throttleZ0Z_10 ));
    InMux I__12362 (
            .O(N__60723),
            .I(N__60720));
    LocalMux I__12361 (
            .O(N__60720),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_2Z0Z_10 ));
    InMux I__12360 (
            .O(N__60717),
            .I(N__60713));
    CascadeMux I__12359 (
            .O(N__60716),
            .I(N__60710));
    LocalMux I__12358 (
            .O(N__60713),
            .I(N__60707));
    InMux I__12357 (
            .O(N__60710),
            .I(N__60704));
    Span4Mux_h I__12356 (
            .O(N__60707),
            .I(N__60700));
    LocalMux I__12355 (
            .O(N__60704),
            .I(N__60697));
    InMux I__12354 (
            .O(N__60703),
            .I(N__60694));
    Span4Mux_h I__12353 (
            .O(N__60700),
            .I(N__60689));
    Span4Mux_v I__12352 (
            .O(N__60697),
            .I(N__60689));
    LocalMux I__12351 (
            .O(N__60694),
            .I(\ppm_encoder_1.throttleZ0Z_8 ));
    Odrv4 I__12350 (
            .O(N__60689),
            .I(\ppm_encoder_1.throttleZ0Z_8 ));
    InMux I__12349 (
            .O(N__60684),
            .I(N__60679));
    InMux I__12348 (
            .O(N__60683),
            .I(N__60676));
    CascadeMux I__12347 (
            .O(N__60682),
            .I(N__60673));
    LocalMux I__12346 (
            .O(N__60679),
            .I(N__60670));
    LocalMux I__12345 (
            .O(N__60676),
            .I(N__60667));
    InMux I__12344 (
            .O(N__60673),
            .I(N__60664));
    Span4Mux_h I__12343 (
            .O(N__60670),
            .I(N__60661));
    Span4Mux_s2_v I__12342 (
            .O(N__60667),
            .I(N__60658));
    LocalMux I__12341 (
            .O(N__60664),
            .I(\ppm_encoder_1.rudderZ0Z_8 ));
    Odrv4 I__12340 (
            .O(N__60661),
            .I(\ppm_encoder_1.rudderZ0Z_8 ));
    Odrv4 I__12339 (
            .O(N__60658),
            .I(\ppm_encoder_1.rudderZ0Z_8 ));
    CascadeMux I__12338 (
            .O(N__60651),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_2Z0Z_8_cascade_ ));
    InMux I__12337 (
            .O(N__60648),
            .I(N__60645));
    LocalMux I__12336 (
            .O(N__60645),
            .I(N__60642));
    Span4Mux_h I__12335 (
            .O(N__60642),
            .I(N__60639));
    Odrv4 I__12334 (
            .O(N__60639),
            .I(\ppm_encoder_1.pulses2count_9_i_2_8 ));
    CascadeMux I__12333 (
            .O(N__60636),
            .I(N__60633));
    InMux I__12332 (
            .O(N__60633),
            .I(N__60630));
    LocalMux I__12331 (
            .O(N__60630),
            .I(N__60627));
    Span4Mux_v I__12330 (
            .O(N__60627),
            .I(N__60624));
    Span4Mux_h I__12329 (
            .O(N__60624),
            .I(N__60621));
    Odrv4 I__12328 (
            .O(N__60621),
            .I(\ppm_encoder_1.pulses2count_9_i_1_9 ));
    CascadeMux I__12327 (
            .O(N__60618),
            .I(N__60615));
    InMux I__12326 (
            .O(N__60615),
            .I(N__60612));
    LocalMux I__12325 (
            .O(N__60612),
            .I(\ppm_encoder_1.pulses2countZ0Z_9 ));
    InMux I__12324 (
            .O(N__60609),
            .I(N__60605));
    InMux I__12323 (
            .O(N__60608),
            .I(N__60602));
    LocalMux I__12322 (
            .O(N__60605),
            .I(N__60598));
    LocalMux I__12321 (
            .O(N__60602),
            .I(N__60595));
    InMux I__12320 (
            .O(N__60601),
            .I(N__60592));
    Odrv12 I__12319 (
            .O(N__60598),
            .I(\ppm_encoder_1.init_pulsesZ0Z_18 ));
    Odrv4 I__12318 (
            .O(N__60595),
            .I(\ppm_encoder_1.init_pulsesZ0Z_18 ));
    LocalMux I__12317 (
            .O(N__60592),
            .I(\ppm_encoder_1.init_pulsesZ0Z_18 ));
    InMux I__12316 (
            .O(N__60585),
            .I(N__60582));
    LocalMux I__12315 (
            .O(N__60582),
            .I(\ppm_encoder_1.pulses2countZ0Z_18 ));
    InMux I__12314 (
            .O(N__60579),
            .I(N__60573));
    CascadeMux I__12313 (
            .O(N__60578),
            .I(N__60570));
    CascadeMux I__12312 (
            .O(N__60577),
            .I(N__60567));
    InMux I__12311 (
            .O(N__60576),
            .I(N__60564));
    LocalMux I__12310 (
            .O(N__60573),
            .I(N__60561));
    InMux I__12309 (
            .O(N__60570),
            .I(N__60556));
    InMux I__12308 (
            .O(N__60567),
            .I(N__60556));
    LocalMux I__12307 (
            .O(N__60564),
            .I(N__60553));
    Span4Mux_s2_v I__12306 (
            .O(N__60561),
            .I(N__60548));
    LocalMux I__12305 (
            .O(N__60556),
            .I(N__60548));
    Odrv12 I__12304 (
            .O(N__60553),
            .I(\ppm_encoder_1.init_pulsesZ0Z_10 ));
    Odrv4 I__12303 (
            .O(N__60548),
            .I(\ppm_encoder_1.init_pulsesZ0Z_10 ));
    InMux I__12302 (
            .O(N__60543),
            .I(N__60540));
    LocalMux I__12301 (
            .O(N__60540),
            .I(\ppm_encoder_1.pulses2count_9_i_0_1_10 ));
    InMux I__12300 (
            .O(N__60537),
            .I(N__60534));
    LocalMux I__12299 (
            .O(N__60534),
            .I(\ppm_encoder_1.pulses2countZ0Z_10 ));
    InMux I__12298 (
            .O(N__60531),
            .I(N__60528));
    LocalMux I__12297 (
            .O(N__60528),
            .I(\ppm_encoder_1.pulses2countZ0Z_11 ));
    InMux I__12296 (
            .O(N__60525),
            .I(N__60522));
    LocalMux I__12295 (
            .O(N__60522),
            .I(N__60519));
    Span4Mux_s1_v I__12294 (
            .O(N__60519),
            .I(N__60516));
    Odrv4 I__12293 (
            .O(N__60516),
            .I(\ppm_encoder_1.counter24_0_I_33_c_RNOZ0 ));
    InMux I__12292 (
            .O(N__60513),
            .I(N__60510));
    LocalMux I__12291 (
            .O(N__60510),
            .I(N__60507));
    Span12Mux_v I__12290 (
            .O(N__60507),
            .I(N__60504));
    Odrv12 I__12289 (
            .O(N__60504),
            .I(\ppm_encoder_1.ppm_output_reg_RNOZ0Z_0 ));
    InMux I__12288 (
            .O(N__60501),
            .I(N__60498));
    LocalMux I__12287 (
            .O(N__60498),
            .I(N__60495));
    Span4Mux_h I__12286 (
            .O(N__60495),
            .I(N__60492));
    Odrv4 I__12285 (
            .O(N__60492),
            .I(\ppm_encoder_1.un1_PPM_STATE_0_sqmuxa_0_i_a2_18_10 ));
    CascadeMux I__12284 (
            .O(N__60489),
            .I(\ppm_encoder_1.un1_PPM_STATE_0_sqmuxa_0_i_a2_18_11_cascade_ ));
    InMux I__12283 (
            .O(N__60486),
            .I(N__60483));
    LocalMux I__12282 (
            .O(N__60483),
            .I(\ppm_encoder_1.un1_PPM_STATE_0_sqmuxa_0_i_a2_18_8 ));
    InMux I__12281 (
            .O(N__60480),
            .I(N__60477));
    LocalMux I__12280 (
            .O(N__60477),
            .I(\ppm_encoder_1.N_486_18 ));
    InMux I__12279 (
            .O(N__60474),
            .I(N__60471));
    LocalMux I__12278 (
            .O(N__60471),
            .I(N__60468));
    Span4Mux_h I__12277 (
            .O(N__60468),
            .I(N__60465));
    Odrv4 I__12276 (
            .O(N__60465),
            .I(\ppm_encoder_1.elevator_RNIC96OZ0Z_5 ));
    CascadeMux I__12275 (
            .O(N__60462),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_2Z0Z_5_cascade_ ));
    InMux I__12274 (
            .O(N__60459),
            .I(N__60456));
    LocalMux I__12273 (
            .O(N__60456),
            .I(N__60452));
    InMux I__12272 (
            .O(N__60455),
            .I(N__60449));
    Span4Mux_h I__12271 (
            .O(N__60452),
            .I(N__60444));
    LocalMux I__12270 (
            .O(N__60449),
            .I(N__60444));
    Span4Mux_h I__12269 (
            .O(N__60444),
            .I(N__60441));
    Odrv4 I__12268 (
            .O(N__60441),
            .I(\ppm_encoder_1.rudderZ0Z_5 ));
    InMux I__12267 (
            .O(N__60438),
            .I(N__60435));
    LocalMux I__12266 (
            .O(N__60435),
            .I(N__60432));
    Span12Mux_h I__12265 (
            .O(N__60432),
            .I(N__60429));
    Odrv12 I__12264 (
            .O(N__60429),
            .I(\ppm_encoder_1.pulses2count_9_i_0_5 ));
    CascadeMux I__12263 (
            .O(N__60426),
            .I(\ppm_encoder_1.pulses2count_9_i_2_5_cascade_ ));
    CascadeMux I__12262 (
            .O(N__60423),
            .I(N__60420));
    InMux I__12261 (
            .O(N__60420),
            .I(N__60417));
    LocalMux I__12260 (
            .O(N__60417),
            .I(\ppm_encoder_1.pulses2countZ0Z_5 ));
    InMux I__12259 (
            .O(N__60414),
            .I(N__60411));
    LocalMux I__12258 (
            .O(N__60411),
            .I(N__60408));
    Span4Mux_h I__12257 (
            .O(N__60408),
            .I(N__60405));
    IoSpan4Mux I__12256 (
            .O(N__60405),
            .I(N__60402));
    Odrv4 I__12255 (
            .O(N__60402),
            .I(\ppm_encoder_1.pulses2count_9_0_0_0 ));
    CascadeMux I__12254 (
            .O(N__60399),
            .I(N__60396));
    InMux I__12253 (
            .O(N__60396),
            .I(N__60393));
    LocalMux I__12252 (
            .O(N__60393),
            .I(N__60390));
    Span4Mux_s3_v I__12251 (
            .O(N__60390),
            .I(N__60387));
    Odrv4 I__12250 (
            .O(N__60387),
            .I(\ppm_encoder_1.pulses2countZ0Z_13 ));
    InMux I__12249 (
            .O(N__60384),
            .I(N__60381));
    LocalMux I__12248 (
            .O(N__60381),
            .I(N__60378));
    Odrv4 I__12247 (
            .O(N__60378),
            .I(\ppm_encoder_1.counter24_0_I_39_c_RNOZ0 ));
    InMux I__12246 (
            .O(N__60375),
            .I(N__60372));
    LocalMux I__12245 (
            .O(N__60372),
            .I(N__60368));
    CascadeMux I__12244 (
            .O(N__60371),
            .I(N__60364));
    Span4Mux_v I__12243 (
            .O(N__60368),
            .I(N__60361));
    InMux I__12242 (
            .O(N__60367),
            .I(N__60358));
    InMux I__12241 (
            .O(N__60364),
            .I(N__60355));
    Span4Mux_h I__12240 (
            .O(N__60361),
            .I(N__60350));
    LocalMux I__12239 (
            .O(N__60358),
            .I(N__60350));
    LocalMux I__12238 (
            .O(N__60355),
            .I(\ppm_encoder_1.aileronZ0Z_12 ));
    Odrv4 I__12237 (
            .O(N__60350),
            .I(\ppm_encoder_1.aileronZ0Z_12 ));
    InMux I__12236 (
            .O(N__60345),
            .I(N__60342));
    LocalMux I__12235 (
            .O(N__60342),
            .I(N__60339));
    Span4Mux_s2_v I__12234 (
            .O(N__60339),
            .I(N__60336));
    Span4Mux_v I__12233 (
            .O(N__60336),
            .I(N__60333));
    Span4Mux_h I__12232 (
            .O(N__60333),
            .I(N__60330));
    Odrv4 I__12231 (
            .O(N__60330),
            .I(\ppm_encoder_1.pulses2count_9_0_3_12 ));
    InMux I__12230 (
            .O(N__60327),
            .I(N__60324));
    LocalMux I__12229 (
            .O(N__60324),
            .I(\ppm_encoder_1.pulses2countZ0Z_12 ));
    InMux I__12228 (
            .O(N__60321),
            .I(N__60318));
    LocalMux I__12227 (
            .O(N__60318),
            .I(N__60315));
    Span4Mux_h I__12226 (
            .O(N__60315),
            .I(N__60312));
    Span4Mux_v I__12225 (
            .O(N__60312),
            .I(N__60309));
    Odrv4 I__12224 (
            .O(N__60309),
            .I(\ppm_encoder_1.pulses2count_9_0_3_11 ));
    CascadeMux I__12223 (
            .O(N__60306),
            .I(N__60303));
    InMux I__12222 (
            .O(N__60303),
            .I(N__60300));
    LocalMux I__12221 (
            .O(N__60300),
            .I(N__60296));
    InMux I__12220 (
            .O(N__60299),
            .I(N__60293));
    Span4Mux_s2_v I__12219 (
            .O(N__60296),
            .I(N__60287));
    LocalMux I__12218 (
            .O(N__60293),
            .I(N__60287));
    InMux I__12217 (
            .O(N__60292),
            .I(N__60284));
    Span4Mux_v I__12216 (
            .O(N__60287),
            .I(N__60281));
    LocalMux I__12215 (
            .O(N__60284),
            .I(\ppm_encoder_1.aileronZ0Z_11 ));
    Odrv4 I__12214 (
            .O(N__60281),
            .I(\ppm_encoder_1.aileronZ0Z_11 ));
    InMux I__12213 (
            .O(N__60276),
            .I(N__60273));
    LocalMux I__12212 (
            .O(N__60273),
            .I(\ppm_encoder_1.counter24_0_I_9_c_RNOZ0 ));
    InMux I__12211 (
            .O(N__60270),
            .I(N__60267));
    LocalMux I__12210 (
            .O(N__60267),
            .I(N__60264));
    Odrv4 I__12209 (
            .O(N__60264),
            .I(\ppm_encoder_1.counter24_0_I_27_c_RNOZ0 ));
    CascadeMux I__12208 (
            .O(N__60261),
            .I(N__60258));
    InMux I__12207 (
            .O(N__60258),
            .I(N__60255));
    LocalMux I__12206 (
            .O(N__60255),
            .I(N__60252));
    Span4Mux_h I__12205 (
            .O(N__60252),
            .I(N__60249));
    Span4Mux_h I__12204 (
            .O(N__60249),
            .I(N__60246));
    Odrv4 I__12203 (
            .O(N__60246),
            .I(\ppm_encoder_1.pulses2count_9_i_1_8 ));
    InMux I__12202 (
            .O(N__60243),
            .I(N__60240));
    LocalMux I__12201 (
            .O(N__60240),
            .I(N__60236));
    CascadeMux I__12200 (
            .O(N__60239),
            .I(N__60232));
    Span4Mux_h I__12199 (
            .O(N__60236),
            .I(N__60228));
    InMux I__12198 (
            .O(N__60235),
            .I(N__60223));
    InMux I__12197 (
            .O(N__60232),
            .I(N__60223));
    InMux I__12196 (
            .O(N__60231),
            .I(N__60220));
    Span4Mux_h I__12195 (
            .O(N__60228),
            .I(N__60215));
    LocalMux I__12194 (
            .O(N__60223),
            .I(N__60215));
    LocalMux I__12193 (
            .O(N__60220),
            .I(\ppm_encoder_1.init_pulsesZ0Z_8 ));
    Odrv4 I__12192 (
            .O(N__60215),
            .I(\ppm_encoder_1.init_pulsesZ0Z_8 ));
    InMux I__12191 (
            .O(N__60210),
            .I(N__60207));
    LocalMux I__12190 (
            .O(N__60207),
            .I(\ppm_encoder_1.pulses2countZ0Z_8 ));
    InMux I__12189 (
            .O(N__60204),
            .I(N__60198));
    InMux I__12188 (
            .O(N__60203),
            .I(N__60198));
    LocalMux I__12187 (
            .O(N__60198),
            .I(N__60192));
    InMux I__12186 (
            .O(N__60197),
            .I(N__60189));
    CascadeMux I__12185 (
            .O(N__60196),
            .I(N__60186));
    InMux I__12184 (
            .O(N__60195),
            .I(N__60181));
    Span4Mux_v I__12183 (
            .O(N__60192),
            .I(N__60178));
    LocalMux I__12182 (
            .O(N__60189),
            .I(N__60175));
    InMux I__12181 (
            .O(N__60186),
            .I(N__60172));
    InMux I__12180 (
            .O(N__60185),
            .I(N__60169));
    CascadeMux I__12179 (
            .O(N__60184),
            .I(N__60166));
    LocalMux I__12178 (
            .O(N__60181),
            .I(N__60162));
    Span4Mux_v I__12177 (
            .O(N__60178),
            .I(N__60157));
    Span4Mux_h I__12176 (
            .O(N__60175),
            .I(N__60157));
    LocalMux I__12175 (
            .O(N__60172),
            .I(N__60154));
    LocalMux I__12174 (
            .O(N__60169),
            .I(N__60151));
    InMux I__12173 (
            .O(N__60166),
            .I(N__60146));
    InMux I__12172 (
            .O(N__60165),
            .I(N__60146));
    Span4Mux_h I__12171 (
            .O(N__60162),
            .I(N__60141));
    Span4Mux_v I__12170 (
            .O(N__60157),
            .I(N__60141));
    Span12Mux_s10_h I__12169 (
            .O(N__60154),
            .I(N__60136));
    Span12Mux_v I__12168 (
            .O(N__60151),
            .I(N__60136));
    LocalMux I__12167 (
            .O(N__60146),
            .I(\pid_front.stateZ0Z_0 ));
    Odrv4 I__12166 (
            .O(N__60141),
            .I(\pid_front.stateZ0Z_0 ));
    Odrv12 I__12165 (
            .O(N__60136),
            .I(\pid_front.stateZ0Z_0 ));
    CascadeMux I__12164 (
            .O(N__60129),
            .I(N__60125));
    CascadeMux I__12163 (
            .O(N__60128),
            .I(N__60122));
    InMux I__12162 (
            .O(N__60125),
            .I(N__60109));
    InMux I__12161 (
            .O(N__60122),
            .I(N__60094));
    InMux I__12160 (
            .O(N__60121),
            .I(N__60094));
    InMux I__12159 (
            .O(N__60120),
            .I(N__60094));
    InMux I__12158 (
            .O(N__60119),
            .I(N__60094));
    InMux I__12157 (
            .O(N__60118),
            .I(N__60094));
    InMux I__12156 (
            .O(N__60117),
            .I(N__60094));
    InMux I__12155 (
            .O(N__60116),
            .I(N__60094));
    InMux I__12154 (
            .O(N__60115),
            .I(N__60090));
    InMux I__12153 (
            .O(N__60114),
            .I(N__60087));
    InMux I__12152 (
            .O(N__60113),
            .I(N__60082));
    InMux I__12151 (
            .O(N__60112),
            .I(N__60082));
    LocalMux I__12150 (
            .O(N__60109),
            .I(N__60076));
    LocalMux I__12149 (
            .O(N__60094),
            .I(N__60076));
    CascadeMux I__12148 (
            .O(N__60093),
            .I(N__60073));
    LocalMux I__12147 (
            .O(N__60090),
            .I(N__60070));
    LocalMux I__12146 (
            .O(N__60087),
            .I(N__60067));
    LocalMux I__12145 (
            .O(N__60082),
            .I(N__60064));
    InMux I__12144 (
            .O(N__60081),
            .I(N__60061));
    Span4Mux_v I__12143 (
            .O(N__60076),
            .I(N__60057));
    InMux I__12142 (
            .O(N__60073),
            .I(N__60054));
    Span4Mux_h I__12141 (
            .O(N__60070),
            .I(N__60051));
    Span4Mux_v I__12140 (
            .O(N__60067),
            .I(N__60048));
    Span4Mux_v I__12139 (
            .O(N__60064),
            .I(N__60045));
    LocalMux I__12138 (
            .O(N__60061),
            .I(N__60042));
    InMux I__12137 (
            .O(N__60060),
            .I(N__60039));
    Span4Mux_h I__12136 (
            .O(N__60057),
            .I(N__60036));
    LocalMux I__12135 (
            .O(N__60054),
            .I(N__60033));
    Span4Mux_h I__12134 (
            .O(N__60051),
            .I(N__60024));
    Span4Mux_v I__12133 (
            .O(N__60048),
            .I(N__60024));
    Span4Mux_h I__12132 (
            .O(N__60045),
            .I(N__60024));
    Span4Mux_h I__12131 (
            .O(N__60042),
            .I(N__60024));
    LocalMux I__12130 (
            .O(N__60039),
            .I(N__60019));
    Span4Mux_v I__12129 (
            .O(N__60036),
            .I(N__60019));
    Span4Mux_h I__12128 (
            .O(N__60033),
            .I(N__60014));
    Span4Mux_v I__12127 (
            .O(N__60024),
            .I(N__60014));
    Odrv4 I__12126 (
            .O(N__60019),
            .I(\pid_front.stateZ0Z_1 ));
    Odrv4 I__12125 (
            .O(N__60014),
            .I(\pid_front.stateZ0Z_1 ));
    CascadeMux I__12124 (
            .O(N__60009),
            .I(\pid_front.N_196_mux_cascade_ ));
    CEMux I__12123 (
            .O(N__60006),
            .I(N__60002));
    CEMux I__12122 (
            .O(N__60005),
            .I(N__59999));
    LocalMux I__12121 (
            .O(N__60002),
            .I(N__59996));
    LocalMux I__12120 (
            .O(N__59999),
            .I(N__59993));
    Span4Mux_v I__12119 (
            .O(N__59996),
            .I(N__59990));
    Span4Mux_h I__12118 (
            .O(N__59993),
            .I(N__59987));
    Sp12to4 I__12117 (
            .O(N__59990),
            .I(N__59984));
    Span4Mux_h I__12116 (
            .O(N__59987),
            .I(N__59981));
    Span12Mux_h I__12115 (
            .O(N__59984),
            .I(N__59978));
    Odrv4 I__12114 (
            .O(N__59981),
            .I(\pid_front.error_i_acumm_1_sqmuxa_1_i ));
    Odrv12 I__12113 (
            .O(N__59978),
            .I(\pid_front.error_i_acumm_1_sqmuxa_1_i ));
    CascadeMux I__12112 (
            .O(N__59973),
            .I(N__59970));
    InMux I__12111 (
            .O(N__59970),
            .I(N__59967));
    LocalMux I__12110 (
            .O(N__59967),
            .I(pid_side_m153_e_5));
    IoInMux I__12109 (
            .O(N__59964),
            .I(N__59961));
    LocalMux I__12108 (
            .O(N__59961),
            .I(N__59958));
    Span4Mux_s0_v I__12107 (
            .O(N__59958),
            .I(N__59955));
    Sp12to4 I__12106 (
            .O(N__59955),
            .I(N__59946));
    InMux I__12105 (
            .O(N__59954),
            .I(N__59941));
    InMux I__12104 (
            .O(N__59953),
            .I(N__59941));
    InMux I__12103 (
            .O(N__59952),
            .I(N__59936));
    InMux I__12102 (
            .O(N__59951),
            .I(N__59936));
    InMux I__12101 (
            .O(N__59950),
            .I(N__59933));
    InMux I__12100 (
            .O(N__59949),
            .I(N__59930));
    Span12Mux_h I__12099 (
            .O(N__59946),
            .I(N__59925));
    LocalMux I__12098 (
            .O(N__59941),
            .I(N__59925));
    LocalMux I__12097 (
            .O(N__59936),
            .I(N__59922));
    LocalMux I__12096 (
            .O(N__59933),
            .I(N__59917));
    LocalMux I__12095 (
            .O(N__59930),
            .I(N__59909));
    Span12Mux_v I__12094 (
            .O(N__59925),
            .I(N__59909));
    Span12Mux_s5_v I__12093 (
            .O(N__59922),
            .I(N__59909));
    InMux I__12092 (
            .O(N__59921),
            .I(N__59904));
    InMux I__12091 (
            .O(N__59920),
            .I(N__59901));
    Span12Mux_s11_v I__12090 (
            .O(N__59917),
            .I(N__59898));
    InMux I__12089 (
            .O(N__59916),
            .I(N__59895));
    Span12Mux_v I__12088 (
            .O(N__59909),
            .I(N__59892));
    InMux I__12087 (
            .O(N__59908),
            .I(N__59887));
    InMux I__12086 (
            .O(N__59907),
            .I(N__59887));
    LocalMux I__12085 (
            .O(N__59904),
            .I(debug_CH1_0A_c));
    LocalMux I__12084 (
            .O(N__59901),
            .I(debug_CH1_0A_c));
    Odrv12 I__12083 (
            .O(N__59898),
            .I(debug_CH1_0A_c));
    LocalMux I__12082 (
            .O(N__59895),
            .I(debug_CH1_0A_c));
    Odrv12 I__12081 (
            .O(N__59892),
            .I(debug_CH1_0A_c));
    LocalMux I__12080 (
            .O(N__59887),
            .I(debug_CH1_0A_c));
    CascadeMux I__12079 (
            .O(N__59874),
            .I(pid_side_m153_e_5_cascade_));
    InMux I__12078 (
            .O(N__59871),
            .I(N__59868));
    LocalMux I__12077 (
            .O(N__59868),
            .I(N__59865));
    Span4Mux_v I__12076 (
            .O(N__59865),
            .I(N__59860));
    CascadeMux I__12075 (
            .O(N__59864),
            .I(N__59856));
    CascadeMux I__12074 (
            .O(N__59863),
            .I(N__59853));
    Span4Mux_v I__12073 (
            .O(N__59860),
            .I(N__59850));
    CascadeMux I__12072 (
            .O(N__59859),
            .I(N__59845));
    InMux I__12071 (
            .O(N__59856),
            .I(N__59839));
    InMux I__12070 (
            .O(N__59853),
            .I(N__59839));
    Span4Mux_v I__12069 (
            .O(N__59850),
            .I(N__59836));
    InMux I__12068 (
            .O(N__59849),
            .I(N__59832));
    InMux I__12067 (
            .O(N__59848),
            .I(N__59827));
    InMux I__12066 (
            .O(N__59845),
            .I(N__59827));
    InMux I__12065 (
            .O(N__59844),
            .I(N__59824));
    LocalMux I__12064 (
            .O(N__59839),
            .I(N__59821));
    Span4Mux_v I__12063 (
            .O(N__59836),
            .I(N__59818));
    InMux I__12062 (
            .O(N__59835),
            .I(N__59815));
    LocalMux I__12061 (
            .O(N__59832),
            .I(\pid_side.stateZ0Z_0 ));
    LocalMux I__12060 (
            .O(N__59827),
            .I(\pid_side.stateZ0Z_0 ));
    LocalMux I__12059 (
            .O(N__59824),
            .I(\pid_side.stateZ0Z_0 ));
    Odrv4 I__12058 (
            .O(N__59821),
            .I(\pid_side.stateZ0Z_0 ));
    Odrv4 I__12057 (
            .O(N__59818),
            .I(\pid_side.stateZ0Z_0 ));
    LocalMux I__12056 (
            .O(N__59815),
            .I(\pid_side.stateZ0Z_0 ));
    InMux I__12055 (
            .O(N__59802),
            .I(N__59799));
    LocalMux I__12054 (
            .O(N__59799),
            .I(N__59796));
    Span4Mux_h I__12053 (
            .O(N__59796),
            .I(N__59793));
    Span4Mux_v I__12052 (
            .O(N__59793),
            .I(N__59790));
    Sp12to4 I__12051 (
            .O(N__59790),
            .I(N__59787));
    Odrv12 I__12050 (
            .O(N__59787),
            .I(\pid_side.N_196_mux ));
    CascadeMux I__12049 (
            .O(N__59784),
            .I(N__59781));
    InMux I__12048 (
            .O(N__59781),
            .I(N__59778));
    LocalMux I__12047 (
            .O(N__59778),
            .I(\ppm_encoder_1.counter24_0_I_15_c_RNOZ0 ));
    CascadeMux I__12046 (
            .O(N__59775),
            .I(N__59772));
    InMux I__12045 (
            .O(N__59772),
            .I(N__59769));
    LocalMux I__12044 (
            .O(N__59769),
            .I(N__59766));
    Span4Mux_v I__12043 (
            .O(N__59766),
            .I(N__59763));
    Span4Mux_h I__12042 (
            .O(N__59763),
            .I(N__59760));
    Odrv4 I__12041 (
            .O(N__59760),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_2Z0Z_4 ));
    InMux I__12040 (
            .O(N__59757),
            .I(N__59754));
    LocalMux I__12039 (
            .O(N__59754),
            .I(N__59750));
    CascadeMux I__12038 (
            .O(N__59753),
            .I(N__59747));
    Span4Mux_h I__12037 (
            .O(N__59750),
            .I(N__59744));
    InMux I__12036 (
            .O(N__59747),
            .I(N__59741));
    Odrv4 I__12035 (
            .O(N__59744),
            .I(\ppm_encoder_1.rudderZ0Z_4 ));
    LocalMux I__12034 (
            .O(N__59741),
            .I(\ppm_encoder_1.rudderZ0Z_4 ));
    InMux I__12033 (
            .O(N__59736),
            .I(N__59733));
    LocalMux I__12032 (
            .O(N__59733),
            .I(N__59730));
    Span4Mux_v I__12031 (
            .O(N__59730),
            .I(N__59727));
    Span4Mux_h I__12030 (
            .O(N__59727),
            .I(N__59724));
    Odrv4 I__12029 (
            .O(N__59724),
            .I(\ppm_encoder_1.pulses2count_9_i_1_4 ));
    CascadeMux I__12028 (
            .O(N__59721),
            .I(\ppm_encoder_1.pulses2count_9_i_2_4_cascade_ ));
    CascadeMux I__12027 (
            .O(N__59718),
            .I(N__59712));
    InMux I__12026 (
            .O(N__59717),
            .I(N__59709));
    InMux I__12025 (
            .O(N__59716),
            .I(N__59706));
    InMux I__12024 (
            .O(N__59715),
            .I(N__59701));
    InMux I__12023 (
            .O(N__59712),
            .I(N__59701));
    LocalMux I__12022 (
            .O(N__59709),
            .I(N__59698));
    LocalMux I__12021 (
            .O(N__59706),
            .I(N__59695));
    LocalMux I__12020 (
            .O(N__59701),
            .I(N__59692));
    Span4Mux_h I__12019 (
            .O(N__59698),
            .I(N__59687));
    Span4Mux_s1_v I__12018 (
            .O(N__59695),
            .I(N__59687));
    Span4Mux_h I__12017 (
            .O(N__59692),
            .I(N__59684));
    Odrv4 I__12016 (
            .O(N__59687),
            .I(\ppm_encoder_1.init_pulsesZ0Z_4 ));
    Odrv4 I__12015 (
            .O(N__59684),
            .I(\ppm_encoder_1.init_pulsesZ0Z_4 ));
    InMux I__12014 (
            .O(N__59679),
            .I(N__59676));
    LocalMux I__12013 (
            .O(N__59676),
            .I(\ppm_encoder_1.pulses2countZ0Z_4 ));
    InMux I__12012 (
            .O(N__59673),
            .I(N__59670));
    LocalMux I__12011 (
            .O(N__59670),
            .I(N__59667));
    Span4Mux_s1_v I__12010 (
            .O(N__59667),
            .I(N__59663));
    CascadeMux I__12009 (
            .O(N__59666),
            .I(N__59658));
    Span4Mux_h I__12008 (
            .O(N__59663),
            .I(N__59655));
    InMux I__12007 (
            .O(N__59662),
            .I(N__59652));
    InMux I__12006 (
            .O(N__59661),
            .I(N__59647));
    InMux I__12005 (
            .O(N__59658),
            .I(N__59647));
    Odrv4 I__12004 (
            .O(N__59655),
            .I(\ppm_encoder_1.init_pulsesZ0Z_5 ));
    LocalMux I__12003 (
            .O(N__59652),
            .I(\ppm_encoder_1.init_pulsesZ0Z_5 ));
    LocalMux I__12002 (
            .O(N__59647),
            .I(\ppm_encoder_1.init_pulsesZ0Z_5 ));
    InMux I__12001 (
            .O(N__59640),
            .I(N__59637));
    LocalMux I__12000 (
            .O(N__59637),
            .I(\pid_front.N_25_0 ));
    CascadeMux I__11999 (
            .O(N__59634),
            .I(\pid_front.error_cry_4_c_RNI81RMZ0Z1_cascade_ ));
    InMux I__11998 (
            .O(N__59631),
            .I(N__59628));
    LocalMux I__11997 (
            .O(N__59628),
            .I(N__59625));
    Odrv4 I__11996 (
            .O(N__59625),
            .I(\pid_front.error_cry_4_c_RNI81RM1Z0Z_0 ));
    CascadeMux I__11995 (
            .O(N__59622),
            .I(\pid_front.N_38_1_cascade_ ));
    InMux I__11994 (
            .O(N__59619),
            .I(N__59615));
    InMux I__11993 (
            .O(N__59618),
            .I(N__59612));
    LocalMux I__11992 (
            .O(N__59615),
            .I(N__59609));
    LocalMux I__11991 (
            .O(N__59612),
            .I(\pid_front.N_37_1 ));
    Odrv4 I__11990 (
            .O(N__59609),
            .I(\pid_front.N_37_1 ));
    CascadeMux I__11989 (
            .O(N__59604),
            .I(\pid_front.N_39_1_cascade_ ));
    CascadeMux I__11988 (
            .O(N__59601),
            .I(N__59598));
    InMux I__11987 (
            .O(N__59598),
            .I(N__59595));
    LocalMux I__11986 (
            .O(N__59595),
            .I(\pid_front.error_i_regZ0Z_10 ));
    InMux I__11985 (
            .O(N__59592),
            .I(N__59589));
    LocalMux I__11984 (
            .O(N__59589),
            .I(\pid_front.N_38_1 ));
    CascadeMux I__11983 (
            .O(N__59586),
            .I(\pid_front.N_110_cascade_ ));
    InMux I__11982 (
            .O(N__59583),
            .I(N__59580));
    LocalMux I__11981 (
            .O(N__59580),
            .I(\pid_front.m2_2_03 ));
    CascadeMux I__11980 (
            .O(N__59577),
            .I(\pid_front.error_i_reg_9_rn_1_14_cascade_ ));
    InMux I__11979 (
            .O(N__59574),
            .I(N__59571));
    LocalMux I__11978 (
            .O(N__59571),
            .I(N__59568));
    Odrv4 I__11977 (
            .O(N__59568),
            .I(\pid_front.N_136 ));
    InMux I__11976 (
            .O(N__59565),
            .I(N__59562));
    LocalMux I__11975 (
            .O(N__59562),
            .I(N__59559));
    Odrv4 I__11974 (
            .O(N__59559),
            .I(\pid_front.error_i_regZ0Z_14 ));
    CascadeMux I__11973 (
            .O(N__59556),
            .I(\pid_front.m10_2_03_3_i_0_cascade_ ));
    InMux I__11972 (
            .O(N__59553),
            .I(N__59550));
    LocalMux I__11971 (
            .O(N__59550),
            .I(N__59547));
    Odrv4 I__11970 (
            .O(N__59547),
            .I(\pid_front.m26_2_03_0 ));
    CascadeMux I__11969 (
            .O(N__59544),
            .I(N__59541));
    InMux I__11968 (
            .O(N__59541),
            .I(N__59538));
    LocalMux I__11967 (
            .O(N__59538),
            .I(\pid_front.error_i_regZ0Z_22 ));
    CascadeMux I__11966 (
            .O(N__59535),
            .I(\pid_front.error_i_reg_esr_RNO_4Z0Z_21_cascade_ ));
    InMux I__11965 (
            .O(N__59532),
            .I(N__59529));
    LocalMux I__11964 (
            .O(N__59529),
            .I(\pid_front.g0_5_1 ));
    CascadeMux I__11963 (
            .O(N__59526),
            .I(\pid_front.N_126_0_cascade_ ));
    InMux I__11962 (
            .O(N__59523),
            .I(N__59520));
    LocalMux I__11961 (
            .O(N__59520),
            .I(\pid_front.N_88_0_0 ));
    CascadeMux I__11960 (
            .O(N__59517),
            .I(\pid_front.m25_2_03_0_cascade_ ));
    InMux I__11959 (
            .O(N__59514),
            .I(N__59510));
    InMux I__11958 (
            .O(N__59513),
            .I(N__59507));
    LocalMux I__11957 (
            .O(N__59510),
            .I(N__59504));
    LocalMux I__11956 (
            .O(N__59507),
            .I(N__59501));
    Odrv4 I__11955 (
            .O(N__59504),
            .I(\pid_front.m9_2_03_3_i_0 ));
    Odrv12 I__11954 (
            .O(N__59501),
            .I(\pid_front.m9_2_03_3_i_0 ));
    InMux I__11953 (
            .O(N__59496),
            .I(N__59493));
    LocalMux I__11952 (
            .O(N__59493),
            .I(\pid_front.error_i_regZ0Z_21 ));
    CascadeMux I__11951 (
            .O(N__59490),
            .I(N__59487));
    InMux I__11950 (
            .O(N__59487),
            .I(N__59484));
    LocalMux I__11949 (
            .O(N__59484),
            .I(\pid_front.error_i_regZ0Z_12 ));
    CascadeMux I__11948 (
            .O(N__59481),
            .I(N__59478));
    InMux I__11947 (
            .O(N__59478),
            .I(N__59475));
    LocalMux I__11946 (
            .O(N__59475),
            .I(\pid_front.error_i_regZ0Z_18 ));
    InMux I__11945 (
            .O(N__59472),
            .I(N__59469));
    LocalMux I__11944 (
            .O(N__59469),
            .I(N__59466));
    Span4Mux_v I__11943 (
            .O(N__59466),
            .I(N__59463));
    Span4Mux_v I__11942 (
            .O(N__59463),
            .I(N__59459));
    InMux I__11941 (
            .O(N__59462),
            .I(N__59456));
    Sp12to4 I__11940 (
            .O(N__59459),
            .I(N__59452));
    LocalMux I__11939 (
            .O(N__59456),
            .I(N__59449));
    InMux I__11938 (
            .O(N__59455),
            .I(N__59446));
    Span12Mux_h I__11937 (
            .O(N__59452),
            .I(N__59441));
    Span12Mux_s7_v I__11936 (
            .O(N__59449),
            .I(N__59441));
    LocalMux I__11935 (
            .O(N__59446),
            .I(N__59438));
    Span12Mux_h I__11934 (
            .O(N__59441),
            .I(N__59432));
    Span4Mux_v I__11933 (
            .O(N__59438),
            .I(N__59429));
    InMux I__11932 (
            .O(N__59437),
            .I(N__59426));
    InMux I__11931 (
            .O(N__59436),
            .I(N__59423));
    InMux I__11930 (
            .O(N__59435),
            .I(N__59420));
    Odrv12 I__11929 (
            .O(N__59432),
            .I(\pid_front.error_9 ));
    Odrv4 I__11928 (
            .O(N__59429),
            .I(\pid_front.error_9 ));
    LocalMux I__11927 (
            .O(N__59426),
            .I(\pid_front.error_9 ));
    LocalMux I__11926 (
            .O(N__59423),
            .I(\pid_front.error_9 ));
    LocalMux I__11925 (
            .O(N__59420),
            .I(\pid_front.error_9 ));
    CascadeMux I__11924 (
            .O(N__59409),
            .I(\pid_front.N_36_0_cascade_ ));
    CascadeMux I__11923 (
            .O(N__59406),
            .I(\pid_front.N_37_1_cascade_ ));
    InMux I__11922 (
            .O(N__59403),
            .I(N__59400));
    LocalMux I__11921 (
            .O(N__59400),
            .I(\pid_front.N_18_1 ));
    InMux I__11920 (
            .O(N__59397),
            .I(N__59394));
    LocalMux I__11919 (
            .O(N__59394),
            .I(\pid_front.error_i_reg_esr_RNO_2_0_16 ));
    CascadeMux I__11918 (
            .O(N__59391),
            .I(\pid_front.error_cry_1_0_c_RNIOOIF3Z0Z_0_cascade_ ));
    CascadeMux I__11917 (
            .O(N__59388),
            .I(\pid_front.N_116_0_cascade_ ));
    InMux I__11916 (
            .O(N__59385),
            .I(N__59382));
    LocalMux I__11915 (
            .O(N__59382),
            .I(\pid_front.error_cry_1_0_c_RNIOOIFZ0Z3 ));
    InMux I__11914 (
            .O(N__59379),
            .I(N__59376));
    LocalMux I__11913 (
            .O(N__59376),
            .I(\pid_front.N_21_1 ));
    CascadeMux I__11912 (
            .O(N__59373),
            .I(\pid_front.error_cry_6_c_RNI1ADU1Z0Z_0_cascade_ ));
    InMux I__11911 (
            .O(N__59370),
            .I(N__59367));
    LocalMux I__11910 (
            .O(N__59367),
            .I(\pid_front.error_cry_6_c_RNI1ADUZ0Z1 ));
    InMux I__11909 (
            .O(N__59364),
            .I(N__59361));
    LocalMux I__11908 (
            .O(N__59361),
            .I(N__59358));
    Odrv4 I__11907 (
            .O(N__59358),
            .I(\pid_front.m4_2_03 ));
    CascadeMux I__11906 (
            .O(N__59355),
            .I(\pid_front.error_i_reg_9_rn_0_16_cascade_ ));
    CascadeMux I__11905 (
            .O(N__59352),
            .I(N__59349));
    InMux I__11904 (
            .O(N__59349),
            .I(N__59346));
    LocalMux I__11903 (
            .O(N__59346),
            .I(N__59343));
    Odrv4 I__11902 (
            .O(N__59343),
            .I(\pid_front.error_i_regZ0Z_16 ));
    InMux I__11901 (
            .O(N__59340),
            .I(N__59337));
    LocalMux I__11900 (
            .O(N__59337),
            .I(\pid_front.error_i_reg_esr_RNO_0Z0Z_16 ));
    InMux I__11899 (
            .O(N__59334),
            .I(N__59329));
    InMux I__11898 (
            .O(N__59333),
            .I(N__59326));
    InMux I__11897 (
            .O(N__59332),
            .I(N__59323));
    LocalMux I__11896 (
            .O(N__59329),
            .I(N__59320));
    LocalMux I__11895 (
            .O(N__59326),
            .I(N__59315));
    LocalMux I__11894 (
            .O(N__59323),
            .I(N__59312));
    Span4Mux_h I__11893 (
            .O(N__59320),
            .I(N__59309));
    InMux I__11892 (
            .O(N__59319),
            .I(N__59304));
    InMux I__11891 (
            .O(N__59318),
            .I(N__59304));
    Span4Mux_v I__11890 (
            .O(N__59315),
            .I(N__59297));
    Span4Mux_h I__11889 (
            .O(N__59312),
            .I(N__59297));
    Span4Mux_v I__11888 (
            .O(N__59309),
            .I(N__59292));
    LocalMux I__11887 (
            .O(N__59304),
            .I(N__59292));
    InMux I__11886 (
            .O(N__59303),
            .I(N__59287));
    InMux I__11885 (
            .O(N__59302),
            .I(N__59287));
    Span4Mux_h I__11884 (
            .O(N__59297),
            .I(N__59281));
    Span4Mux_h I__11883 (
            .O(N__59292),
            .I(N__59281));
    LocalMux I__11882 (
            .O(N__59287),
            .I(N__59278));
    InMux I__11881 (
            .O(N__59286),
            .I(N__59275));
    Span4Mux_v I__11880 (
            .O(N__59281),
            .I(N__59271));
    Span12Mux_h I__11879 (
            .O(N__59278),
            .I(N__59266));
    LocalMux I__11878 (
            .O(N__59275),
            .I(N__59266));
    InMux I__11877 (
            .O(N__59274),
            .I(N__59263));
    Odrv4 I__11876 (
            .O(N__59271),
            .I(uart_drone_data_0));
    Odrv12 I__11875 (
            .O(N__59266),
            .I(uart_drone_data_0));
    LocalMux I__11874 (
            .O(N__59263),
            .I(uart_drone_data_0));
    InMux I__11873 (
            .O(N__59256),
            .I(N__59253));
    LocalMux I__11872 (
            .O(N__59253),
            .I(dron_frame_decoder_1_source_H_disp_front_fast_0));
    CEMux I__11871 (
            .O(N__59250),
            .I(N__59247));
    LocalMux I__11870 (
            .O(N__59247),
            .I(N__59243));
    CEMux I__11869 (
            .O(N__59246),
            .I(N__59240));
    Span4Mux_v I__11868 (
            .O(N__59243),
            .I(N__59235));
    LocalMux I__11867 (
            .O(N__59240),
            .I(N__59235));
    Span4Mux_v I__11866 (
            .O(N__59235),
            .I(N__59232));
    Odrv4 I__11865 (
            .O(N__59232),
            .I(\dron_frame_decoder_1.N_708_0 ));
    InMux I__11864 (
            .O(N__59229),
            .I(N__59226));
    LocalMux I__11863 (
            .O(N__59226),
            .I(N__59223));
    Span4Mux_h I__11862 (
            .O(N__59223),
            .I(N__59220));
    Span4Mux_v I__11861 (
            .O(N__59220),
            .I(N__59217));
    Odrv4 I__11860 (
            .O(N__59217),
            .I(\pid_side.un4_error_i_reg_31_ns_1_0 ));
    InMux I__11859 (
            .O(N__59214),
            .I(N__59211));
    LocalMux I__11858 (
            .O(N__59211),
            .I(\pid_front.m11_0_ns_1 ));
    CascadeMux I__11857 (
            .O(N__59208),
            .I(\pid_front.N_48_1_cascade_ ));
    InMux I__11856 (
            .O(N__59205),
            .I(N__59201));
    InMux I__11855 (
            .O(N__59204),
            .I(N__59198));
    LocalMux I__11854 (
            .O(N__59201),
            .I(N__59192));
    LocalMux I__11853 (
            .O(N__59198),
            .I(N__59189));
    InMux I__11852 (
            .O(N__59197),
            .I(N__59186));
    InMux I__11851 (
            .O(N__59196),
            .I(N__59183));
    InMux I__11850 (
            .O(N__59195),
            .I(N__59179));
    Span4Mux_v I__11849 (
            .O(N__59192),
            .I(N__59176));
    Span4Mux_v I__11848 (
            .O(N__59189),
            .I(N__59173));
    LocalMux I__11847 (
            .O(N__59186),
            .I(N__59168));
    LocalMux I__11846 (
            .O(N__59183),
            .I(N__59168));
    InMux I__11845 (
            .O(N__59182),
            .I(N__59163));
    LocalMux I__11844 (
            .O(N__59179),
            .I(N__59160));
    Span4Mux_h I__11843 (
            .O(N__59176),
            .I(N__59157));
    Span4Mux_v I__11842 (
            .O(N__59173),
            .I(N__59154));
    Span4Mux_v I__11841 (
            .O(N__59168),
            .I(N__59151));
    CascadeMux I__11840 (
            .O(N__59167),
            .I(N__59148));
    InMux I__11839 (
            .O(N__59166),
            .I(N__59144));
    LocalMux I__11838 (
            .O(N__59163),
            .I(N__59139));
    Span12Mux_h I__11837 (
            .O(N__59160),
            .I(N__59139));
    Span4Mux_v I__11836 (
            .O(N__59157),
            .I(N__59136));
    Span4Mux_h I__11835 (
            .O(N__59154),
            .I(N__59131));
    Span4Mux_v I__11834 (
            .O(N__59151),
            .I(N__59131));
    InMux I__11833 (
            .O(N__59148),
            .I(N__59128));
    InMux I__11832 (
            .O(N__59147),
            .I(N__59125));
    LocalMux I__11831 (
            .O(N__59144),
            .I(uart_drone_data_1));
    Odrv12 I__11830 (
            .O(N__59139),
            .I(uart_drone_data_1));
    Odrv4 I__11829 (
            .O(N__59136),
            .I(uart_drone_data_1));
    Odrv4 I__11828 (
            .O(N__59131),
            .I(uart_drone_data_1));
    LocalMux I__11827 (
            .O(N__59128),
            .I(uart_drone_data_1));
    LocalMux I__11826 (
            .O(N__59125),
            .I(uart_drone_data_1));
    InMux I__11825 (
            .O(N__59112),
            .I(N__59109));
    LocalMux I__11824 (
            .O(N__59109),
            .I(drone_H_disp_front_1));
    InMux I__11823 (
            .O(N__59106),
            .I(N__59101));
    InMux I__11822 (
            .O(N__59105),
            .I(N__59098));
    InMux I__11821 (
            .O(N__59104),
            .I(N__59095));
    LocalMux I__11820 (
            .O(N__59101),
            .I(N__59090));
    LocalMux I__11819 (
            .O(N__59098),
            .I(N__59087));
    LocalMux I__11818 (
            .O(N__59095),
            .I(N__59084));
    InMux I__11817 (
            .O(N__59094),
            .I(N__59081));
    InMux I__11816 (
            .O(N__59093),
            .I(N__59078));
    Span4Mux_v I__11815 (
            .O(N__59090),
            .I(N__59075));
    Span4Mux_h I__11814 (
            .O(N__59087),
            .I(N__59072));
    Span4Mux_v I__11813 (
            .O(N__59084),
            .I(N__59067));
    LocalMux I__11812 (
            .O(N__59081),
            .I(N__59067));
    LocalMux I__11811 (
            .O(N__59078),
            .I(N__59064));
    Span4Mux_h I__11810 (
            .O(N__59075),
            .I(N__59056));
    Span4Mux_v I__11809 (
            .O(N__59072),
            .I(N__59056));
    Span4Mux_h I__11808 (
            .O(N__59067),
            .I(N__59056));
    Span4Mux_h I__11807 (
            .O(N__59064),
            .I(N__59053));
    InMux I__11806 (
            .O(N__59063),
            .I(N__59050));
    Span4Mux_v I__11805 (
            .O(N__59056),
            .I(N__59046));
    Sp12to4 I__11804 (
            .O(N__59053),
            .I(N__59041));
    LocalMux I__11803 (
            .O(N__59050),
            .I(N__59041));
    InMux I__11802 (
            .O(N__59049),
            .I(N__59038));
    Odrv4 I__11801 (
            .O(N__59046),
            .I(uart_drone_data_2));
    Odrv12 I__11800 (
            .O(N__59041),
            .I(uart_drone_data_2));
    LocalMux I__11799 (
            .O(N__59038),
            .I(uart_drone_data_2));
    InMux I__11798 (
            .O(N__59031),
            .I(N__59028));
    LocalMux I__11797 (
            .O(N__59028),
            .I(drone_H_disp_front_2));
    InMux I__11796 (
            .O(N__59025),
            .I(N__59020));
    InMux I__11795 (
            .O(N__59024),
            .I(N__59017));
    InMux I__11794 (
            .O(N__59023),
            .I(N__59013));
    LocalMux I__11793 (
            .O(N__59020),
            .I(N__59009));
    LocalMux I__11792 (
            .O(N__59017),
            .I(N__59006));
    InMux I__11791 (
            .O(N__59016),
            .I(N__59003));
    LocalMux I__11790 (
            .O(N__59013),
            .I(N__59000));
    InMux I__11789 (
            .O(N__59012),
            .I(N__58997));
    Span4Mux_v I__11788 (
            .O(N__59009),
            .I(N__58994));
    Span4Mux_h I__11787 (
            .O(N__59006),
            .I(N__58991));
    LocalMux I__11786 (
            .O(N__59003),
            .I(N__58988));
    Span4Mux_v I__11785 (
            .O(N__59000),
            .I(N__58983));
    LocalMux I__11784 (
            .O(N__58997),
            .I(N__58983));
    Span4Mux_h I__11783 (
            .O(N__58994),
            .I(N__58975));
    Span4Mux_v I__11782 (
            .O(N__58991),
            .I(N__58975));
    Span4Mux_h I__11781 (
            .O(N__58988),
            .I(N__58975));
    Span4Mux_h I__11780 (
            .O(N__58983),
            .I(N__58972));
    InMux I__11779 (
            .O(N__58982),
            .I(N__58969));
    Span4Mux_v I__11778 (
            .O(N__58975),
            .I(N__58963));
    Sp12to4 I__11777 (
            .O(N__58972),
            .I(N__58958));
    LocalMux I__11776 (
            .O(N__58969),
            .I(N__58958));
    InMux I__11775 (
            .O(N__58968),
            .I(N__58955));
    InMux I__11774 (
            .O(N__58967),
            .I(N__58950));
    InMux I__11773 (
            .O(N__58966),
            .I(N__58950));
    Odrv4 I__11772 (
            .O(N__58963),
            .I(uart_drone_data_3));
    Odrv12 I__11771 (
            .O(N__58958),
            .I(uart_drone_data_3));
    LocalMux I__11770 (
            .O(N__58955),
            .I(uart_drone_data_3));
    LocalMux I__11769 (
            .O(N__58950),
            .I(uart_drone_data_3));
    InMux I__11768 (
            .O(N__58941),
            .I(N__58938));
    LocalMux I__11767 (
            .O(N__58938),
            .I(drone_H_disp_front_3));
    InMux I__11766 (
            .O(N__58935),
            .I(N__58931));
    InMux I__11765 (
            .O(N__58934),
            .I(N__58925));
    LocalMux I__11764 (
            .O(N__58931),
            .I(N__58922));
    InMux I__11763 (
            .O(N__58930),
            .I(N__58919));
    InMux I__11762 (
            .O(N__58929),
            .I(N__58915));
    InMux I__11761 (
            .O(N__58928),
            .I(N__58912));
    LocalMux I__11760 (
            .O(N__58925),
            .I(N__58909));
    Span4Mux_v I__11759 (
            .O(N__58922),
            .I(N__58906));
    LocalMux I__11758 (
            .O(N__58919),
            .I(N__58903));
    InMux I__11757 (
            .O(N__58918),
            .I(N__58900));
    LocalMux I__11756 (
            .O(N__58915),
            .I(N__58897));
    LocalMux I__11755 (
            .O(N__58912),
            .I(N__58894));
    Span4Mux_v I__11754 (
            .O(N__58909),
            .I(N__58891));
    Span4Mux_h I__11753 (
            .O(N__58906),
            .I(N__58888));
    Span4Mux_v I__11752 (
            .O(N__58903),
            .I(N__58885));
    LocalMux I__11751 (
            .O(N__58900),
            .I(N__58878));
    Span4Mux_h I__11750 (
            .O(N__58897),
            .I(N__58878));
    Span4Mux_v I__11749 (
            .O(N__58894),
            .I(N__58878));
    Span4Mux_v I__11748 (
            .O(N__58891),
            .I(N__58870));
    Span4Mux_v I__11747 (
            .O(N__58888),
            .I(N__58870));
    Span4Mux_h I__11746 (
            .O(N__58885),
            .I(N__58865));
    Span4Mux_v I__11745 (
            .O(N__58878),
            .I(N__58865));
    InMux I__11744 (
            .O(N__58877),
            .I(N__58862));
    InMux I__11743 (
            .O(N__58876),
            .I(N__58857));
    InMux I__11742 (
            .O(N__58875),
            .I(N__58857));
    Odrv4 I__11741 (
            .O(N__58870),
            .I(uart_drone_data_4));
    Odrv4 I__11740 (
            .O(N__58865),
            .I(uart_drone_data_4));
    LocalMux I__11739 (
            .O(N__58862),
            .I(uart_drone_data_4));
    LocalMux I__11738 (
            .O(N__58857),
            .I(uart_drone_data_4));
    InMux I__11737 (
            .O(N__58848),
            .I(N__58845));
    LocalMux I__11736 (
            .O(N__58845),
            .I(\dron_frame_decoder_1.drone_H_disp_front_4 ));
    InMux I__11735 (
            .O(N__58842),
            .I(N__58838));
    InMux I__11734 (
            .O(N__58841),
            .I(N__58835));
    LocalMux I__11733 (
            .O(N__58838),
            .I(N__58830));
    LocalMux I__11732 (
            .O(N__58835),
            .I(N__58826));
    InMux I__11731 (
            .O(N__58834),
            .I(N__58822));
    InMux I__11730 (
            .O(N__58833),
            .I(N__58819));
    Span4Mux_v I__11729 (
            .O(N__58830),
            .I(N__58816));
    InMux I__11728 (
            .O(N__58829),
            .I(N__58813));
    Span4Mux_v I__11727 (
            .O(N__58826),
            .I(N__58810));
    InMux I__11726 (
            .O(N__58825),
            .I(N__58807));
    LocalMux I__11725 (
            .O(N__58822),
            .I(N__58804));
    LocalMux I__11724 (
            .O(N__58819),
            .I(N__58801));
    Span4Mux_v I__11723 (
            .O(N__58816),
            .I(N__58796));
    LocalMux I__11722 (
            .O(N__58813),
            .I(N__58796));
    Span4Mux_h I__11721 (
            .O(N__58810),
            .I(N__58791));
    LocalMux I__11720 (
            .O(N__58807),
            .I(N__58791));
    Span12Mux_s11_h I__11719 (
            .O(N__58804),
            .I(N__58787));
    Span12Mux_v I__11718 (
            .O(N__58801),
            .I(N__58784));
    Span4Mux_v I__11717 (
            .O(N__58796),
            .I(N__58781));
    Span4Mux_v I__11716 (
            .O(N__58791),
            .I(N__58778));
    InMux I__11715 (
            .O(N__58790),
            .I(N__58775));
    Odrv12 I__11714 (
            .O(N__58787),
            .I(uart_drone_data_5));
    Odrv12 I__11713 (
            .O(N__58784),
            .I(uart_drone_data_5));
    Odrv4 I__11712 (
            .O(N__58781),
            .I(uart_drone_data_5));
    Odrv4 I__11711 (
            .O(N__58778),
            .I(uart_drone_data_5));
    LocalMux I__11710 (
            .O(N__58775),
            .I(uart_drone_data_5));
    InMux I__11709 (
            .O(N__58764),
            .I(N__58761));
    LocalMux I__11708 (
            .O(N__58761),
            .I(\dron_frame_decoder_1.drone_H_disp_front_5 ));
    InMux I__11707 (
            .O(N__58758),
            .I(N__58754));
    InMux I__11706 (
            .O(N__58757),
            .I(N__58749));
    LocalMux I__11705 (
            .O(N__58754),
            .I(N__58746));
    InMux I__11704 (
            .O(N__58753),
            .I(N__58743));
    InMux I__11703 (
            .O(N__58752),
            .I(N__58739));
    LocalMux I__11702 (
            .O(N__58749),
            .I(N__58735));
    Span4Mux_v I__11701 (
            .O(N__58746),
            .I(N__58732));
    LocalMux I__11700 (
            .O(N__58743),
            .I(N__58729));
    InMux I__11699 (
            .O(N__58742),
            .I(N__58726));
    LocalMux I__11698 (
            .O(N__58739),
            .I(N__58722));
    CascadeMux I__11697 (
            .O(N__58738),
            .I(N__58719));
    Span4Mux_v I__11696 (
            .O(N__58735),
            .I(N__58716));
    Span4Mux_h I__11695 (
            .O(N__58732),
            .I(N__58713));
    Span4Mux_v I__11694 (
            .O(N__58729),
            .I(N__58708));
    LocalMux I__11693 (
            .O(N__58726),
            .I(N__58708));
    InMux I__11692 (
            .O(N__58725),
            .I(N__58705));
    Span4Mux_v I__11691 (
            .O(N__58722),
            .I(N__58702));
    InMux I__11690 (
            .O(N__58719),
            .I(N__58699));
    Span4Mux_h I__11689 (
            .O(N__58716),
            .I(N__58694));
    Span4Mux_v I__11688 (
            .O(N__58713),
            .I(N__58689));
    Span4Mux_v I__11687 (
            .O(N__58708),
            .I(N__58689));
    LocalMux I__11686 (
            .O(N__58705),
            .I(N__58686));
    Span4Mux_v I__11685 (
            .O(N__58702),
            .I(N__58681));
    LocalMux I__11684 (
            .O(N__58699),
            .I(N__58681));
    InMux I__11683 (
            .O(N__58698),
            .I(N__58676));
    InMux I__11682 (
            .O(N__58697),
            .I(N__58676));
    Odrv4 I__11681 (
            .O(N__58694),
            .I(uart_drone_data_6));
    Odrv4 I__11680 (
            .O(N__58689),
            .I(uart_drone_data_6));
    Odrv12 I__11679 (
            .O(N__58686),
            .I(uart_drone_data_6));
    Odrv4 I__11678 (
            .O(N__58681),
            .I(uart_drone_data_6));
    LocalMux I__11677 (
            .O(N__58676),
            .I(uart_drone_data_6));
    InMux I__11676 (
            .O(N__58665),
            .I(N__58662));
    LocalMux I__11675 (
            .O(N__58662),
            .I(\dron_frame_decoder_1.drone_H_disp_front_6 ));
    InMux I__11674 (
            .O(N__58659),
            .I(N__58655));
    InMux I__11673 (
            .O(N__58658),
            .I(N__58652));
    LocalMux I__11672 (
            .O(N__58655),
            .I(N__58648));
    LocalMux I__11671 (
            .O(N__58652),
            .I(N__58645));
    InMux I__11670 (
            .O(N__58651),
            .I(N__58640));
    Span4Mux_v I__11669 (
            .O(N__58648),
            .I(N__58635));
    Span4Mux_h I__11668 (
            .O(N__58645),
            .I(N__58635));
    InMux I__11667 (
            .O(N__58644),
            .I(N__58631));
    InMux I__11666 (
            .O(N__58643),
            .I(N__58628));
    LocalMux I__11665 (
            .O(N__58640),
            .I(N__58624));
    Span4Mux_h I__11664 (
            .O(N__58635),
            .I(N__58621));
    InMux I__11663 (
            .O(N__58634),
            .I(N__58618));
    LocalMux I__11662 (
            .O(N__58631),
            .I(N__58615));
    LocalMux I__11661 (
            .O(N__58628),
            .I(N__58612));
    CascadeMux I__11660 (
            .O(N__58627),
            .I(N__58609));
    Span4Mux_v I__11659 (
            .O(N__58624),
            .I(N__58606));
    Span4Mux_v I__11658 (
            .O(N__58621),
            .I(N__58603));
    LocalMux I__11657 (
            .O(N__58618),
            .I(N__58596));
    Span12Mux_h I__11656 (
            .O(N__58615),
            .I(N__58596));
    Span12Mux_s11_h I__11655 (
            .O(N__58612),
            .I(N__58596));
    InMux I__11654 (
            .O(N__58609),
            .I(N__58593));
    Odrv4 I__11653 (
            .O(N__58606),
            .I(uart_drone_data_7));
    Odrv4 I__11652 (
            .O(N__58603),
            .I(uart_drone_data_7));
    Odrv12 I__11651 (
            .O(N__58596),
            .I(uart_drone_data_7));
    LocalMux I__11650 (
            .O(N__58593),
            .I(uart_drone_data_7));
    InMux I__11649 (
            .O(N__58584),
            .I(N__58581));
    LocalMux I__11648 (
            .O(N__58581),
            .I(\dron_frame_decoder_1.drone_H_disp_front_7 ));
    CascadeMux I__11647 (
            .O(N__58578),
            .I(\pid_front.m0_0_03_cascade_ ));
    InMux I__11646 (
            .O(N__58575),
            .I(N__58572));
    LocalMux I__11645 (
            .O(N__58572),
            .I(\dron_frame_decoder_1.drone_H_disp_side_5 ));
    InMux I__11644 (
            .O(N__58569),
            .I(N__58566));
    LocalMux I__11643 (
            .O(N__58566),
            .I(\dron_frame_decoder_1.drone_H_disp_side_6 ));
    InMux I__11642 (
            .O(N__58563),
            .I(N__58560));
    LocalMux I__11641 (
            .O(N__58560),
            .I(\dron_frame_decoder_1.drone_H_disp_side_7 ));
    InMux I__11640 (
            .O(N__58557),
            .I(N__58554));
    LocalMux I__11639 (
            .O(N__58554),
            .I(N__58551));
    Span4Mux_h I__11638 (
            .O(N__58551),
            .I(N__58548));
    Odrv4 I__11637 (
            .O(N__58548),
            .I(\pid_side.N_88_0_0 ));
    CascadeMux I__11636 (
            .O(N__58545),
            .I(\pid_side.error_cry_5_c_RNIN1DBZ0Z2_cascade_ ));
    InMux I__11635 (
            .O(N__58542),
            .I(N__58539));
    LocalMux I__11634 (
            .O(N__58539),
            .I(\pid_side.error_cry_5_c_RNIN1DB2Z0Z_0 ));
    CascadeMux I__11633 (
            .O(N__58536),
            .I(\pid_side.N_103_0_cascade_ ));
    InMux I__11632 (
            .O(N__58533),
            .I(N__58529));
    InMux I__11631 (
            .O(N__58532),
            .I(N__58526));
    LocalMux I__11630 (
            .O(N__58529),
            .I(N__58523));
    LocalMux I__11629 (
            .O(N__58526),
            .I(\pid_side.N_53_0 ));
    Odrv4 I__11628 (
            .O(N__58523),
            .I(\pid_side.N_53_0 ));
    CascadeMux I__11627 (
            .O(N__58518),
            .I(\pid_side.N_50_1_cascade_ ));
    InMux I__11626 (
            .O(N__58515),
            .I(N__58512));
    LocalMux I__11625 (
            .O(N__58512),
            .I(N__58508));
    InMux I__11624 (
            .O(N__58511),
            .I(N__58505));
    Odrv4 I__11623 (
            .O(N__58508),
            .I(\pid_side.N_50_1 ));
    LocalMux I__11622 (
            .O(N__58505),
            .I(\pid_side.N_50_1 ));
    InMux I__11621 (
            .O(N__58500),
            .I(N__58497));
    LocalMux I__11620 (
            .O(N__58497),
            .I(N__58494));
    Odrv4 I__11619 (
            .O(N__58494),
            .I(\pid_side.error_i_reg_9_rn_0_27 ));
    InMux I__11618 (
            .O(N__58491),
            .I(N__58488));
    LocalMux I__11617 (
            .O(N__58488),
            .I(\dron_frame_decoder_1.drone_H_disp_side_4 ));
    InMux I__11616 (
            .O(N__58485),
            .I(N__58482));
    LocalMux I__11615 (
            .O(N__58482),
            .I(\pid_side.error_cry_1_0_c_RNIEAJZ0Z82 ));
    CascadeMux I__11614 (
            .O(N__58479),
            .I(\pid_side.error_cry_1_0_c_RNIEAJ82Z0Z_0_cascade_ ));
    CascadeMux I__11613 (
            .O(N__58476),
            .I(\pid_side.N_39_0_cascade_ ));
    InMux I__11612 (
            .O(N__58473),
            .I(N__58470));
    LocalMux I__11611 (
            .O(N__58470),
            .I(N__58467));
    Odrv4 I__11610 (
            .O(N__58467),
            .I(\pid_side.m7_2_03 ));
    CascadeMux I__11609 (
            .O(N__58464),
            .I(\pid_side.m134_0_ns_1_cascade_ ));
    CascadeMux I__11608 (
            .O(N__58461),
            .I(\pid_side.m19_2_03_0_cascade_ ));
    InMux I__11607 (
            .O(N__58458),
            .I(N__58455));
    LocalMux I__11606 (
            .O(N__58455),
            .I(\pid_side.g1 ));
    CascadeMux I__11605 (
            .O(N__58452),
            .I(\pid_side.g3_cascade_ ));
    CascadeMux I__11604 (
            .O(N__58449),
            .I(\pid_side.m37_1_ns_1_cascade_ ));
    CascadeMux I__11603 (
            .O(N__58446),
            .I(\pid_side.N_38_1_cascade_ ));
    CascadeMux I__11602 (
            .O(N__58443),
            .I(\pid_side.error_i_reg_esr_RNO_3Z0Z_22_cascade_ ));
    InMux I__11601 (
            .O(N__58440),
            .I(N__58437));
    LocalMux I__11600 (
            .O(N__58437),
            .I(\pid_side.error_i_reg_esr_RNO_2Z0Z_22 ));
    InMux I__11599 (
            .O(N__58434),
            .I(N__58431));
    LocalMux I__11598 (
            .O(N__58431),
            .I(\pid_side.error_i_reg_esr_RNO_1Z0Z_22 ));
    InMux I__11597 (
            .O(N__58428),
            .I(N__58425));
    LocalMux I__11596 (
            .O(N__58425),
            .I(N__58421));
    InMux I__11595 (
            .O(N__58424),
            .I(N__58418));
    Odrv4 I__11594 (
            .O(N__58421),
            .I(\pid_side.N_37_1 ));
    LocalMux I__11593 (
            .O(N__58418),
            .I(\pid_side.N_37_1 ));
    CascadeMux I__11592 (
            .O(N__58413),
            .I(\pid_side.m136_ns_1_cascade_ ));
    InMux I__11591 (
            .O(N__58410),
            .I(N__58407));
    LocalMux I__11590 (
            .O(N__58407),
            .I(\pid_side.m18_2_03_4 ));
    CascadeMux I__11589 (
            .O(N__58404),
            .I(\pid_side.error_p_reg_esr_RNIIFTC1Z0Z_6_cascade_ ));
    InMux I__11588 (
            .O(N__58401),
            .I(N__58398));
    LocalMux I__11587 (
            .O(N__58398),
            .I(\pid_side.error_p_reg_esr_RNINKTC1_0Z0Z_7 ));
    InMux I__11586 (
            .O(N__58395),
            .I(N__58389));
    InMux I__11585 (
            .O(N__58394),
            .I(N__58389));
    LocalMux I__11584 (
            .O(N__58389),
            .I(N__58386));
    Span12Mux_v I__11583 (
            .O(N__58386),
            .I(N__58383));
    Odrv12 I__11582 (
            .O(N__58383),
            .I(\pid_side.N_2368_i ));
    InMux I__11581 (
            .O(N__58380),
            .I(N__58371));
    InMux I__11580 (
            .O(N__58379),
            .I(N__58371));
    InMux I__11579 (
            .O(N__58378),
            .I(N__58371));
    LocalMux I__11578 (
            .O(N__58371),
            .I(\pid_side.error_d_reg_prevZ0Z_6 ));
    CascadeMux I__11577 (
            .O(N__58368),
            .I(\pid_side.error_p_reg_esr_RNINKTC1Z0Z_7_cascade_ ));
    CascadeMux I__11576 (
            .O(N__58365),
            .I(\pid_side.error_i_reg_9_rn_0_19_cascade_ ));
    CascadeMux I__11575 (
            .O(N__58362),
            .I(\pid_side.m2_2_03_cascade_ ));
    CascadeMux I__11574 (
            .O(N__58359),
            .I(\pid_side.error_i_acumm_prereg_esr_RNIGSJVZ0Z_7_cascade_ ));
    InMux I__11573 (
            .O(N__58356),
            .I(N__58353));
    LocalMux I__11572 (
            .O(N__58353),
            .I(\pid_side.error_i_acumm_prereg_esr_RNIJ04N_0Z0Z_10 ));
    CascadeMux I__11571 (
            .O(N__58350),
            .I(\pid_side.error_p_reg_esr_RNINKTC1_0Z0Z_7_cascade_ ));
    CascadeMux I__11570 (
            .O(N__58347),
            .I(\pid_side.N_2362_i_cascade_ ));
    InMux I__11569 (
            .O(N__58344),
            .I(N__58341));
    LocalMux I__11568 (
            .O(N__58341),
            .I(\pid_side.error_p_reg_esr_RNIIFTC1Z0Z_6 ));
    InMux I__11567 (
            .O(N__58338),
            .I(N__58335));
    LocalMux I__11566 (
            .O(N__58335),
            .I(N__58332));
    Span4Mux_v I__11565 (
            .O(N__58332),
            .I(N__58329));
    Span4Mux_h I__11564 (
            .O(N__58329),
            .I(N__58325));
    InMux I__11563 (
            .O(N__58328),
            .I(N__58322));
    Sp12to4 I__11562 (
            .O(N__58325),
            .I(N__58317));
    LocalMux I__11561 (
            .O(N__58322),
            .I(N__58317));
    Odrv12 I__11560 (
            .O(N__58317),
            .I(side_order_12));
    InMux I__11559 (
            .O(N__58314),
            .I(N__58311));
    LocalMux I__11558 (
            .O(N__58311),
            .I(N__58307));
    InMux I__11557 (
            .O(N__58310),
            .I(N__58304));
    Span4Mux_h I__11556 (
            .O(N__58307),
            .I(N__58301));
    LocalMux I__11555 (
            .O(N__58304),
            .I(N__58298));
    Odrv4 I__11554 (
            .O(N__58301),
            .I(side_order_13));
    Odrv12 I__11553 (
            .O(N__58298),
            .I(side_order_13));
    CEMux I__11552 (
            .O(N__58293),
            .I(N__58288));
    CEMux I__11551 (
            .O(N__58292),
            .I(N__58285));
    CEMux I__11550 (
            .O(N__58291),
            .I(N__58282));
    LocalMux I__11549 (
            .O(N__58288),
            .I(N__58278));
    LocalMux I__11548 (
            .O(N__58285),
            .I(N__58275));
    LocalMux I__11547 (
            .O(N__58282),
            .I(N__58272));
    CEMux I__11546 (
            .O(N__58281),
            .I(N__58269));
    Span4Mux_v I__11545 (
            .O(N__58278),
            .I(N__58266));
    Span4Mux_h I__11544 (
            .O(N__58275),
            .I(N__58261));
    Span4Mux_h I__11543 (
            .O(N__58272),
            .I(N__58261));
    LocalMux I__11542 (
            .O(N__58269),
            .I(N__58258));
    Odrv4 I__11541 (
            .O(N__58266),
            .I(\pid_side.state_0_1 ));
    Odrv4 I__11540 (
            .O(N__58261),
            .I(\pid_side.state_0_1 ));
    Odrv4 I__11539 (
            .O(N__58258),
            .I(\pid_side.state_0_1 ));
    SRMux I__11538 (
            .O(N__58251),
            .I(N__58248));
    LocalMux I__11537 (
            .O(N__58248),
            .I(N__58242));
    SRMux I__11536 (
            .O(N__58247),
            .I(N__58239));
    SRMux I__11535 (
            .O(N__58246),
            .I(N__58236));
    SRMux I__11534 (
            .O(N__58245),
            .I(N__58233));
    Span4Mux_h I__11533 (
            .O(N__58242),
            .I(N__58230));
    LocalMux I__11532 (
            .O(N__58239),
            .I(N__58227));
    LocalMux I__11531 (
            .O(N__58236),
            .I(N__58224));
    LocalMux I__11530 (
            .O(N__58233),
            .I(N__58221));
    Span4Mux_h I__11529 (
            .O(N__58230),
            .I(N__58218));
    Span4Mux_h I__11528 (
            .O(N__58227),
            .I(N__58215));
    Odrv4 I__11527 (
            .O(N__58224),
            .I(\pid_side.un1_reset_0_i ));
    Odrv4 I__11526 (
            .O(N__58221),
            .I(\pid_side.un1_reset_0_i ));
    Odrv4 I__11525 (
            .O(N__58218),
            .I(\pid_side.un1_reset_0_i ));
    Odrv4 I__11524 (
            .O(N__58215),
            .I(\pid_side.un1_reset_0_i ));
    CascadeMux I__11523 (
            .O(N__58206),
            .I(\pid_side.state_ns_0_cascade_ ));
    CascadeMux I__11522 (
            .O(N__58203),
            .I(N__58199));
    InMux I__11521 (
            .O(N__58202),
            .I(N__58196));
    InMux I__11520 (
            .O(N__58199),
            .I(N__58193));
    LocalMux I__11519 (
            .O(N__58196),
            .I(N__58188));
    LocalMux I__11518 (
            .O(N__58193),
            .I(N__58188));
    Span4Mux_h I__11517 (
            .O(N__58188),
            .I(N__58185));
    Odrv4 I__11516 (
            .O(N__58185),
            .I(side_order_6));
    InMux I__11515 (
            .O(N__58182),
            .I(N__58178));
    InMux I__11514 (
            .O(N__58181),
            .I(N__58175));
    LocalMux I__11513 (
            .O(N__58178),
            .I(N__58172));
    LocalMux I__11512 (
            .O(N__58175),
            .I(N__58169));
    Span4Mux_h I__11511 (
            .O(N__58172),
            .I(N__58166));
    Odrv12 I__11510 (
            .O(N__58169),
            .I(side_order_2));
    Odrv4 I__11509 (
            .O(N__58166),
            .I(side_order_2));
    CascadeMux I__11508 (
            .O(N__58161),
            .I(\pid_side.un1_reset_0_i_cascade_ ));
    CascadeMux I__11507 (
            .O(N__58158),
            .I(N__58153));
    CascadeMux I__11506 (
            .O(N__58157),
            .I(N__58148));
    InMux I__11505 (
            .O(N__58156),
            .I(N__58145));
    InMux I__11504 (
            .O(N__58153),
            .I(N__58136));
    InMux I__11503 (
            .O(N__58152),
            .I(N__58136));
    InMux I__11502 (
            .O(N__58151),
            .I(N__58136));
    InMux I__11501 (
            .O(N__58148),
            .I(N__58136));
    LocalMux I__11500 (
            .O(N__58145),
            .I(\pid_side.N_75 ));
    LocalMux I__11499 (
            .O(N__58136),
            .I(\pid_side.N_75 ));
    CascadeMux I__11498 (
            .O(N__58131),
            .I(\pid_side.N_75_cascade_ ));
    InMux I__11497 (
            .O(N__58128),
            .I(N__58125));
    LocalMux I__11496 (
            .O(N__58125),
            .I(\pid_side.N_102 ));
    CascadeMux I__11495 (
            .O(N__58122),
            .I(N__58115));
    CascadeMux I__11494 (
            .O(N__58121),
            .I(N__58112));
    CascadeMux I__11493 (
            .O(N__58120),
            .I(N__58104));
    InMux I__11492 (
            .O(N__58119),
            .I(N__58097));
    InMux I__11491 (
            .O(N__58118),
            .I(N__58097));
    InMux I__11490 (
            .O(N__58115),
            .I(N__58092));
    InMux I__11489 (
            .O(N__58112),
            .I(N__58092));
    InMux I__11488 (
            .O(N__58111),
            .I(N__58075));
    InMux I__11487 (
            .O(N__58110),
            .I(N__58075));
    InMux I__11486 (
            .O(N__58109),
            .I(N__58075));
    InMux I__11485 (
            .O(N__58108),
            .I(N__58075));
    InMux I__11484 (
            .O(N__58107),
            .I(N__58075));
    InMux I__11483 (
            .O(N__58104),
            .I(N__58075));
    InMux I__11482 (
            .O(N__58103),
            .I(N__58075));
    InMux I__11481 (
            .O(N__58102),
            .I(N__58075));
    LocalMux I__11480 (
            .O(N__58097),
            .I(\pid_side.N_76 ));
    LocalMux I__11479 (
            .O(N__58092),
            .I(\pid_side.N_76 ));
    LocalMux I__11478 (
            .O(N__58075),
            .I(\pid_side.N_76 ));
    InMux I__11477 (
            .O(N__58068),
            .I(N__58064));
    CascadeMux I__11476 (
            .O(N__58067),
            .I(N__58061));
    LocalMux I__11475 (
            .O(N__58064),
            .I(N__58057));
    InMux I__11474 (
            .O(N__58061),
            .I(N__58054));
    CascadeMux I__11473 (
            .O(N__58060),
            .I(N__58051));
    Span4Mux_v I__11472 (
            .O(N__58057),
            .I(N__58046));
    LocalMux I__11471 (
            .O(N__58054),
            .I(N__58046));
    InMux I__11470 (
            .O(N__58051),
            .I(N__58043));
    Span4Mux_h I__11469 (
            .O(N__58046),
            .I(N__58040));
    LocalMux I__11468 (
            .O(N__58043),
            .I(\ppm_encoder_1.elevatorZ0Z_2 ));
    Odrv4 I__11467 (
            .O(N__58040),
            .I(\ppm_encoder_1.elevatorZ0Z_2 ));
    InMux I__11466 (
            .O(N__58035),
            .I(N__58029));
    InMux I__11465 (
            .O(N__58034),
            .I(N__58029));
    LocalMux I__11464 (
            .O(N__58029),
            .I(N__58025));
    InMux I__11463 (
            .O(N__58028),
            .I(N__58022));
    Span4Mux_v I__11462 (
            .O(N__58025),
            .I(N__58019));
    LocalMux I__11461 (
            .O(N__58022),
            .I(\ppm_encoder_1.elevatorZ0Z_1 ));
    Odrv4 I__11460 (
            .O(N__58019),
            .I(\ppm_encoder_1.elevatorZ0Z_1 ));
    InMux I__11459 (
            .O(N__58014),
            .I(N__58006));
    InMux I__11458 (
            .O(N__58013),
            .I(N__58001));
    InMux I__11457 (
            .O(N__58012),
            .I(N__57998));
    InMux I__11456 (
            .O(N__58011),
            .I(N__57995));
    InMux I__11455 (
            .O(N__58010),
            .I(N__57991));
    InMux I__11454 (
            .O(N__58009),
            .I(N__57987));
    LocalMux I__11453 (
            .O(N__58006),
            .I(N__57984));
    InMux I__11452 (
            .O(N__58005),
            .I(N__57979));
    InMux I__11451 (
            .O(N__58004),
            .I(N__57975));
    LocalMux I__11450 (
            .O(N__58001),
            .I(N__57970));
    LocalMux I__11449 (
            .O(N__57998),
            .I(N__57970));
    LocalMux I__11448 (
            .O(N__57995),
            .I(N__57967));
    InMux I__11447 (
            .O(N__57994),
            .I(N__57964));
    LocalMux I__11446 (
            .O(N__57991),
            .I(N__57960));
    InMux I__11445 (
            .O(N__57990),
            .I(N__57957));
    LocalMux I__11444 (
            .O(N__57987),
            .I(N__57952));
    Span4Mux_h I__11443 (
            .O(N__57984),
            .I(N__57952));
    InMux I__11442 (
            .O(N__57983),
            .I(N__57949));
    InMux I__11441 (
            .O(N__57982),
            .I(N__57946));
    LocalMux I__11440 (
            .O(N__57979),
            .I(N__57943));
    InMux I__11439 (
            .O(N__57978),
            .I(N__57940));
    LocalMux I__11438 (
            .O(N__57975),
            .I(N__57931));
    Span4Mux_v I__11437 (
            .O(N__57970),
            .I(N__57931));
    Span4Mux_h I__11436 (
            .O(N__57967),
            .I(N__57931));
    LocalMux I__11435 (
            .O(N__57964),
            .I(N__57931));
    InMux I__11434 (
            .O(N__57963),
            .I(N__57928));
    Odrv4 I__11433 (
            .O(N__57960),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIJQ7DZ0Z_1 ));
    LocalMux I__11432 (
            .O(N__57957),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIJQ7DZ0Z_1 ));
    Odrv4 I__11431 (
            .O(N__57952),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIJQ7DZ0Z_1 ));
    LocalMux I__11430 (
            .O(N__57949),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIJQ7DZ0Z_1 ));
    LocalMux I__11429 (
            .O(N__57946),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIJQ7DZ0Z_1 ));
    Odrv4 I__11428 (
            .O(N__57943),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIJQ7DZ0Z_1 ));
    LocalMux I__11427 (
            .O(N__57940),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIJQ7DZ0Z_1 ));
    Odrv4 I__11426 (
            .O(N__57931),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIJQ7DZ0Z_1 ));
    LocalMux I__11425 (
            .O(N__57928),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIJQ7DZ0Z_1 ));
    CascadeMux I__11424 (
            .O(N__57909),
            .I(N__57906));
    InMux I__11423 (
            .O(N__57906),
            .I(N__57901));
    InMux I__11422 (
            .O(N__57905),
            .I(N__57896));
    InMux I__11421 (
            .O(N__57904),
            .I(N__57896));
    LocalMux I__11420 (
            .O(N__57901),
            .I(N__57893));
    LocalMux I__11419 (
            .O(N__57896),
            .I(\ppm_encoder_1.throttleZ0Z_1 ));
    Odrv4 I__11418 (
            .O(N__57893),
            .I(\ppm_encoder_1.throttleZ0Z_1 ));
    InMux I__11417 (
            .O(N__57888),
            .I(N__57885));
    LocalMux I__11416 (
            .O(N__57885),
            .I(N__57882));
    Odrv4 I__11415 (
            .O(N__57882),
            .I(\ppm_encoder_1.throttle_RNI2JJC1Z0Z_1 ));
    InMux I__11414 (
            .O(N__57879),
            .I(N__57876));
    LocalMux I__11413 (
            .O(N__57876),
            .I(N__57873));
    Odrv12 I__11412 (
            .O(N__57873),
            .I(\ppm_encoder_1.counter24_0_I_21_c_RNOZ0 ));
    InMux I__11411 (
            .O(N__57870),
            .I(N__57866));
    CascadeMux I__11410 (
            .O(N__57869),
            .I(N__57863));
    LocalMux I__11409 (
            .O(N__57866),
            .I(N__57859));
    InMux I__11408 (
            .O(N__57863),
            .I(N__57856));
    InMux I__11407 (
            .O(N__57862),
            .I(N__57853));
    Span4Mux_v I__11406 (
            .O(N__57859),
            .I(N__57848));
    LocalMux I__11405 (
            .O(N__57856),
            .I(N__57848));
    LocalMux I__11404 (
            .O(N__57853),
            .I(\ppm_encoder_1.rudderZ0Z_7 ));
    Odrv4 I__11403 (
            .O(N__57848),
            .I(\ppm_encoder_1.rudderZ0Z_7 ));
    InMux I__11402 (
            .O(N__57843),
            .I(N__57840));
    LocalMux I__11401 (
            .O(N__57840),
            .I(N__57837));
    Span4Mux_v I__11400 (
            .O(N__57837),
            .I(N__57834));
    Odrv4 I__11399 (
            .O(N__57834),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_2Z0Z_7 ));
    InMux I__11398 (
            .O(N__57831),
            .I(N__57828));
    LocalMux I__11397 (
            .O(N__57828),
            .I(N__57825));
    Span4Mux_h I__11396 (
            .O(N__57825),
            .I(N__57821));
    InMux I__11395 (
            .O(N__57824),
            .I(N__57818));
    Odrv4 I__11394 (
            .O(N__57821),
            .I(\ppm_encoder_1.elevator_RNIEB6OZ0Z_7 ));
    LocalMux I__11393 (
            .O(N__57818),
            .I(\ppm_encoder_1.elevator_RNIEB6OZ0Z_7 ));
    InMux I__11392 (
            .O(N__57813),
            .I(N__57810));
    LocalMux I__11391 (
            .O(N__57810),
            .I(\ppm_encoder_1.pulses2count_9_i_0_7 ));
    CascadeMux I__11390 (
            .O(N__57807),
            .I(\ppm_encoder_1.pulses2count_9_i_2_7_cascade_ ));
    CascadeMux I__11389 (
            .O(N__57804),
            .I(N__57801));
    InMux I__11388 (
            .O(N__57801),
            .I(N__57798));
    LocalMux I__11387 (
            .O(N__57798),
            .I(\ppm_encoder_1.pulses2countZ0Z_7 ));
    InMux I__11386 (
            .O(N__57795),
            .I(N__57791));
    CascadeMux I__11385 (
            .O(N__57794),
            .I(N__57788));
    LocalMux I__11384 (
            .O(N__57791),
            .I(N__57785));
    InMux I__11383 (
            .O(N__57788),
            .I(N__57782));
    Span4Mux_h I__11382 (
            .O(N__57785),
            .I(N__57778));
    LocalMux I__11381 (
            .O(N__57782),
            .I(N__57775));
    InMux I__11380 (
            .O(N__57781),
            .I(N__57772));
    Span4Mux_h I__11379 (
            .O(N__57778),
            .I(N__57767));
    Span4Mux_h I__11378 (
            .O(N__57775),
            .I(N__57767));
    LocalMux I__11377 (
            .O(N__57772),
            .I(\ppm_encoder_1.rudderZ0Z_6 ));
    Odrv4 I__11376 (
            .O(N__57767),
            .I(\ppm_encoder_1.rudderZ0Z_6 ));
    InMux I__11375 (
            .O(N__57762),
            .I(N__57759));
    LocalMux I__11374 (
            .O(N__57759),
            .I(N__57755));
    InMux I__11373 (
            .O(N__57758),
            .I(N__57752));
    Span4Mux_h I__11372 (
            .O(N__57755),
            .I(N__57749));
    LocalMux I__11371 (
            .O(N__57752),
            .I(N__57746));
    Odrv4 I__11370 (
            .O(N__57749),
            .I(\ppm_encoder_1.elevator_RNIDA6OZ0Z_6 ));
    Odrv4 I__11369 (
            .O(N__57746),
            .I(\ppm_encoder_1.elevator_RNIDA6OZ0Z_6 ));
    CascadeMux I__11368 (
            .O(N__57741),
            .I(\ppm_encoder_1.pulses2count_9_0_2_6_cascade_ ));
    InMux I__11367 (
            .O(N__57738),
            .I(N__57735));
    LocalMux I__11366 (
            .O(N__57735),
            .I(\ppm_encoder_1.pulses2countZ0Z_6 ));
    InMux I__11365 (
            .O(N__57732),
            .I(N__57729));
    LocalMux I__11364 (
            .O(N__57729),
            .I(\ppm_encoder_1.pulses2count_9_0_2_13 ));
    CascadeMux I__11363 (
            .O(N__57726),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_2_cascade_ ));
    InMux I__11362 (
            .O(N__57723),
            .I(N__57720));
    LocalMux I__11361 (
            .O(N__57720),
            .I(N__57717));
    Span4Mux_h I__11360 (
            .O(N__57717),
            .I(N__57714));
    Odrv4 I__11359 (
            .O(N__57714),
            .I(\ppm_encoder_1.init_pulses_RNI5GAI5Z0Z_2 ));
    InMux I__11358 (
            .O(N__57711),
            .I(N__57707));
    InMux I__11357 (
            .O(N__57710),
            .I(N__57704));
    LocalMux I__11356 (
            .O(N__57707),
            .I(N__57699));
    LocalMux I__11355 (
            .O(N__57704),
            .I(N__57696));
    InMux I__11354 (
            .O(N__57703),
            .I(N__57691));
    InMux I__11353 (
            .O(N__57702),
            .I(N__57691));
    Span4Mux_s3_v I__11352 (
            .O(N__57699),
            .I(N__57682));
    Span4Mux_s3_v I__11351 (
            .O(N__57696),
            .I(N__57682));
    LocalMux I__11350 (
            .O(N__57691),
            .I(N__57682));
    CascadeMux I__11349 (
            .O(N__57690),
            .I(N__57676));
    CascadeMux I__11348 (
            .O(N__57689),
            .I(N__57673));
    Span4Mux_h I__11347 (
            .O(N__57682),
            .I(N__57670));
    InMux I__11346 (
            .O(N__57681),
            .I(N__57667));
    InMux I__11345 (
            .O(N__57680),
            .I(N__57662));
    InMux I__11344 (
            .O(N__57679),
            .I(N__57662));
    InMux I__11343 (
            .O(N__57676),
            .I(N__57657));
    InMux I__11342 (
            .O(N__57673),
            .I(N__57657));
    Odrv4 I__11341 (
            .O(N__57670),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_3_repZ0Z1 ));
    LocalMux I__11340 (
            .O(N__57667),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_3_repZ0Z1 ));
    LocalMux I__11339 (
            .O(N__57662),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_3_repZ0Z1 ));
    LocalMux I__11338 (
            .O(N__57657),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_3_repZ0Z1 ));
    CascadeMux I__11337 (
            .O(N__57648),
            .I(N__57644));
    InMux I__11336 (
            .O(N__57647),
            .I(N__57641));
    InMux I__11335 (
            .O(N__57644),
            .I(N__57638));
    LocalMux I__11334 (
            .O(N__57641),
            .I(N__57635));
    LocalMux I__11333 (
            .O(N__57638),
            .I(N__57632));
    Span4Mux_s1_v I__11332 (
            .O(N__57635),
            .I(N__57629));
    Span4Mux_s2_v I__11331 (
            .O(N__57632),
            .I(N__57626));
    Span4Mux_h I__11330 (
            .O(N__57629),
            .I(N__57621));
    Span4Mux_h I__11329 (
            .O(N__57626),
            .I(N__57618));
    InMux I__11328 (
            .O(N__57625),
            .I(N__57613));
    InMux I__11327 (
            .O(N__57624),
            .I(N__57613));
    Odrv4 I__11326 (
            .O(N__57621),
            .I(\ppm_encoder_1.N_259_i_i ));
    Odrv4 I__11325 (
            .O(N__57618),
            .I(\ppm_encoder_1.N_259_i_i ));
    LocalMux I__11324 (
            .O(N__57613),
            .I(\ppm_encoder_1.N_259_i_i ));
    InMux I__11323 (
            .O(N__57606),
            .I(N__57603));
    LocalMux I__11322 (
            .O(N__57603),
            .I(N__57598));
    CascadeMux I__11321 (
            .O(N__57602),
            .I(N__57594));
    InMux I__11320 (
            .O(N__57601),
            .I(N__57590));
    Span4Mux_s2_v I__11319 (
            .O(N__57598),
            .I(N__57587));
    InMux I__11318 (
            .O(N__57597),
            .I(N__57580));
    InMux I__11317 (
            .O(N__57594),
            .I(N__57580));
    InMux I__11316 (
            .O(N__57593),
            .I(N__57580));
    LocalMux I__11315 (
            .O(N__57590),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_1 ));
    Odrv4 I__11314 (
            .O(N__57587),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_1 ));
    LocalMux I__11313 (
            .O(N__57580),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_1 ));
    CascadeMux I__11312 (
            .O(N__57573),
            .I(N__57569));
    InMux I__11311 (
            .O(N__57572),
            .I(N__57566));
    InMux I__11310 (
            .O(N__57569),
            .I(N__57563));
    LocalMux I__11309 (
            .O(N__57566),
            .I(N__57560));
    LocalMux I__11308 (
            .O(N__57563),
            .I(N__57557));
    Span4Mux_h I__11307 (
            .O(N__57560),
            .I(N__57554));
    Span4Mux_v I__11306 (
            .O(N__57557),
            .I(N__57551));
    Span4Mux_h I__11305 (
            .O(N__57554),
            .I(N__57548));
    Span4Mux_h I__11304 (
            .O(N__57551),
            .I(N__57545));
    Odrv4 I__11303 (
            .O(N__57548),
            .I(\ppm_encoder_1.throttleZ0Z_14 ));
    Odrv4 I__11302 (
            .O(N__57545),
            .I(\ppm_encoder_1.throttleZ0Z_14 ));
    InMux I__11301 (
            .O(N__57540),
            .I(N__57537));
    LocalMux I__11300 (
            .O(N__57537),
            .I(N__57533));
    InMux I__11299 (
            .O(N__57536),
            .I(N__57530));
    Span4Mux_h I__11298 (
            .O(N__57533),
            .I(N__57527));
    LocalMux I__11297 (
            .O(N__57530),
            .I(N__57524));
    Span4Mux_v I__11296 (
            .O(N__57527),
            .I(N__57521));
    Span12Mux_s9_v I__11295 (
            .O(N__57524),
            .I(N__57518));
    Odrv4 I__11294 (
            .O(N__57521),
            .I(\ppm_encoder_1.aileronZ0Z_14 ));
    Odrv12 I__11293 (
            .O(N__57518),
            .I(\ppm_encoder_1.aileronZ0Z_14 ));
    CascadeMux I__11292 (
            .O(N__57513),
            .I(\ppm_encoder_1.pulses2count_9_i_0_14_cascade_ ));
    InMux I__11291 (
            .O(N__57510),
            .I(N__57506));
    CascadeMux I__11290 (
            .O(N__57509),
            .I(N__57502));
    LocalMux I__11289 (
            .O(N__57506),
            .I(N__57499));
    InMux I__11288 (
            .O(N__57505),
            .I(N__57494));
    InMux I__11287 (
            .O(N__57502),
            .I(N__57494));
    Span4Mux_v I__11286 (
            .O(N__57499),
            .I(N__57488));
    LocalMux I__11285 (
            .O(N__57494),
            .I(N__57488));
    InMux I__11284 (
            .O(N__57493),
            .I(N__57485));
    Span4Mux_h I__11283 (
            .O(N__57488),
            .I(N__57482));
    LocalMux I__11282 (
            .O(N__57485),
            .I(\ppm_encoder_1.init_pulsesZ0Z_14 ));
    Odrv4 I__11281 (
            .O(N__57482),
            .I(\ppm_encoder_1.init_pulsesZ0Z_14 ));
    CascadeMux I__11280 (
            .O(N__57477),
            .I(\ppm_encoder_1.pulses2count_9_i_1_14_cascade_ ));
    InMux I__11279 (
            .O(N__57474),
            .I(N__57471));
    LocalMux I__11278 (
            .O(N__57471),
            .I(N__57467));
    InMux I__11277 (
            .O(N__57470),
            .I(N__57464));
    Span4Mux_v I__11276 (
            .O(N__57467),
            .I(N__57461));
    LocalMux I__11275 (
            .O(N__57464),
            .I(N__57458));
    Odrv4 I__11274 (
            .O(N__57461),
            .I(\ppm_encoder_1.elevator_esr_RNI6C0M1Z0Z_14 ));
    Odrv4 I__11273 (
            .O(N__57458),
            .I(\ppm_encoder_1.elevator_esr_RNI6C0M1Z0Z_14 ));
    CascadeMux I__11272 (
            .O(N__57453),
            .I(N__57450));
    InMux I__11271 (
            .O(N__57450),
            .I(N__57446));
    CascadeMux I__11270 (
            .O(N__57449),
            .I(N__57443));
    LocalMux I__11269 (
            .O(N__57446),
            .I(N__57440));
    InMux I__11268 (
            .O(N__57443),
            .I(N__57437));
    Span4Mux_v I__11267 (
            .O(N__57440),
            .I(N__57431));
    LocalMux I__11266 (
            .O(N__57437),
            .I(N__57431));
    InMux I__11265 (
            .O(N__57436),
            .I(N__57428));
    Span4Mux_h I__11264 (
            .O(N__57431),
            .I(N__57425));
    LocalMux I__11263 (
            .O(N__57428),
            .I(N__57422));
    Odrv4 I__11262 (
            .O(N__57425),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_ns_0 ));
    Odrv12 I__11261 (
            .O(N__57422),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_ns_0 ));
    CascadeMux I__11260 (
            .O(N__57417),
            .I(N__57413));
    InMux I__11259 (
            .O(N__57416),
            .I(N__57410));
    InMux I__11258 (
            .O(N__57413),
            .I(N__57407));
    LocalMux I__11257 (
            .O(N__57410),
            .I(N__57403));
    LocalMux I__11256 (
            .O(N__57407),
            .I(N__57400));
    InMux I__11255 (
            .O(N__57406),
            .I(N__57397));
    Span4Mux_v I__11254 (
            .O(N__57403),
            .I(N__57392));
    Span4Mux_h I__11253 (
            .O(N__57400),
            .I(N__57392));
    LocalMux I__11252 (
            .O(N__57397),
            .I(N__57389));
    Span4Mux_v I__11251 (
            .O(N__57392),
            .I(N__57386));
    Span4Mux_h I__11250 (
            .O(N__57389),
            .I(N__57383));
    Odrv4 I__11249 (
            .O(N__57386),
            .I(\ppm_encoder_1.N_56 ));
    Odrv4 I__11248 (
            .O(N__57383),
            .I(\ppm_encoder_1.N_56 ));
    CascadeMux I__11247 (
            .O(N__57378),
            .I(N__57374));
    InMux I__11246 (
            .O(N__57377),
            .I(N__57371));
    InMux I__11245 (
            .O(N__57374),
            .I(N__57368));
    LocalMux I__11244 (
            .O(N__57371),
            .I(N__57365));
    LocalMux I__11243 (
            .O(N__57368),
            .I(N__57362));
    Span4Mux_v I__11242 (
            .O(N__57365),
            .I(N__57356));
    Span4Mux_h I__11241 (
            .O(N__57362),
            .I(N__57356));
    InMux I__11240 (
            .O(N__57361),
            .I(N__57353));
    Span4Mux_h I__11239 (
            .O(N__57356),
            .I(N__57350));
    LocalMux I__11238 (
            .O(N__57353),
            .I(\ppm_encoder_1.throttleZ0Z_11 ));
    Odrv4 I__11237 (
            .O(N__57350),
            .I(\ppm_encoder_1.throttleZ0Z_11 ));
    InMux I__11236 (
            .O(N__57345),
            .I(N__57342));
    LocalMux I__11235 (
            .O(N__57342),
            .I(N__57339));
    Span4Mux_s2_v I__11234 (
            .O(N__57339),
            .I(N__57336));
    Odrv4 I__11233 (
            .O(N__57336),
            .I(\ppm_encoder_1.un2_throttle_iv_0_1_11 ));
    InMux I__11232 (
            .O(N__57333),
            .I(N__57327));
    InMux I__11231 (
            .O(N__57332),
            .I(N__57324));
    InMux I__11230 (
            .O(N__57331),
            .I(N__57321));
    InMux I__11229 (
            .O(N__57330),
            .I(N__57318));
    LocalMux I__11228 (
            .O(N__57327),
            .I(N__57315));
    LocalMux I__11227 (
            .O(N__57324),
            .I(N__57312));
    LocalMux I__11226 (
            .O(N__57321),
            .I(N__57309));
    LocalMux I__11225 (
            .O(N__57318),
            .I(N__57306));
    Span4Mux_v I__11224 (
            .O(N__57315),
            .I(N__57301));
    Span4Mux_h I__11223 (
            .O(N__57312),
            .I(N__57301));
    Span4Mux_h I__11222 (
            .O(N__57309),
            .I(N__57298));
    Span4Mux_h I__11221 (
            .O(N__57306),
            .I(N__57295));
    Odrv4 I__11220 (
            .O(N__57301),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIM4C21Z0Z_2 ));
    Odrv4 I__11219 (
            .O(N__57298),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIM4C21Z0Z_2 ));
    Odrv4 I__11218 (
            .O(N__57295),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIM4C21Z0Z_2 ));
    CascadeMux I__11217 (
            .O(N__57288),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIM4C21Z0Z_2_cascade_ ));
    CascadeMux I__11216 (
            .O(N__57285),
            .I(N__57282));
    InMux I__11215 (
            .O(N__57282),
            .I(N__57279));
    LocalMux I__11214 (
            .O(N__57279),
            .I(N__57276));
    Span4Mux_h I__11213 (
            .O(N__57276),
            .I(N__57273));
    Odrv4 I__11212 (
            .O(N__57273),
            .I(\ppm_encoder_1.init_pulses_RNIN1203Z0Z_2 ));
    InMux I__11211 (
            .O(N__57270),
            .I(N__57267));
    LocalMux I__11210 (
            .O(N__57267),
            .I(N__57263));
    CascadeMux I__11209 (
            .O(N__57266),
            .I(N__57258));
    Span4Mux_s3_v I__11208 (
            .O(N__57263),
            .I(N__57250));
    InMux I__11207 (
            .O(N__57262),
            .I(N__57247));
    InMux I__11206 (
            .O(N__57261),
            .I(N__57244));
    InMux I__11205 (
            .O(N__57258),
            .I(N__57239));
    InMux I__11204 (
            .O(N__57257),
            .I(N__57239));
    InMux I__11203 (
            .O(N__57256),
            .I(N__57234));
    InMux I__11202 (
            .O(N__57255),
            .I(N__57234));
    InMux I__11201 (
            .O(N__57254),
            .I(N__57229));
    InMux I__11200 (
            .O(N__57253),
            .I(N__57229));
    Odrv4 I__11199 (
            .O(N__57250),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2 ));
    LocalMux I__11198 (
            .O(N__57247),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2 ));
    LocalMux I__11197 (
            .O(N__57244),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2 ));
    LocalMux I__11196 (
            .O(N__57239),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2 ));
    LocalMux I__11195 (
            .O(N__57234),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2 ));
    LocalMux I__11194 (
            .O(N__57229),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2 ));
    CascadeMux I__11193 (
            .O(N__57216),
            .I(N__57213));
    InMux I__11192 (
            .O(N__57213),
            .I(N__57206));
    InMux I__11191 (
            .O(N__57212),
            .I(N__57203));
    InMux I__11190 (
            .O(N__57211),
            .I(N__57200));
    InMux I__11189 (
            .O(N__57210),
            .I(N__57195));
    InMux I__11188 (
            .O(N__57209),
            .I(N__57195));
    LocalMux I__11187 (
            .O(N__57206),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0 ));
    LocalMux I__11186 (
            .O(N__57203),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0 ));
    LocalMux I__11185 (
            .O(N__57200),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0 ));
    LocalMux I__11184 (
            .O(N__57195),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0 ));
    InMux I__11183 (
            .O(N__57186),
            .I(N__57179));
    InMux I__11182 (
            .O(N__57185),
            .I(N__57176));
    InMux I__11181 (
            .O(N__57184),
            .I(N__57173));
    InMux I__11180 (
            .O(N__57183),
            .I(N__57170));
    InMux I__11179 (
            .O(N__57182),
            .I(N__57167));
    LocalMux I__11178 (
            .O(N__57179),
            .I(N__57163));
    LocalMux I__11177 (
            .O(N__57176),
            .I(N__57160));
    LocalMux I__11176 (
            .O(N__57173),
            .I(N__57152));
    LocalMux I__11175 (
            .O(N__57170),
            .I(N__57148));
    LocalMux I__11174 (
            .O(N__57167),
            .I(N__57145));
    InMux I__11173 (
            .O(N__57166),
            .I(N__57141));
    Span4Mux_v I__11172 (
            .O(N__57163),
            .I(N__57136));
    Span4Mux_s1_v I__11171 (
            .O(N__57160),
            .I(N__57136));
    InMux I__11170 (
            .O(N__57159),
            .I(N__57133));
    InMux I__11169 (
            .O(N__57158),
            .I(N__57128));
    InMux I__11168 (
            .O(N__57157),
            .I(N__57128));
    InMux I__11167 (
            .O(N__57156),
            .I(N__57125));
    InMux I__11166 (
            .O(N__57155),
            .I(N__57119));
    Span4Mux_v I__11165 (
            .O(N__57152),
            .I(N__57116));
    InMux I__11164 (
            .O(N__57151),
            .I(N__57113));
    Span4Mux_v I__11163 (
            .O(N__57148),
            .I(N__57108));
    Span4Mux_v I__11162 (
            .O(N__57145),
            .I(N__57108));
    InMux I__11161 (
            .O(N__57144),
            .I(N__57105));
    LocalMux I__11160 (
            .O(N__57141),
            .I(N__57100));
    Span4Mux_h I__11159 (
            .O(N__57136),
            .I(N__57100));
    LocalMux I__11158 (
            .O(N__57133),
            .I(N__57093));
    LocalMux I__11157 (
            .O(N__57128),
            .I(N__57093));
    LocalMux I__11156 (
            .O(N__57125),
            .I(N__57093));
    InMux I__11155 (
            .O(N__57124),
            .I(N__57086));
    InMux I__11154 (
            .O(N__57123),
            .I(N__57086));
    InMux I__11153 (
            .O(N__57122),
            .I(N__57086));
    LocalMux I__11152 (
            .O(N__57119),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIIP7DZ0Z_0 ));
    Odrv4 I__11151 (
            .O(N__57116),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIIP7DZ0Z_0 ));
    LocalMux I__11150 (
            .O(N__57113),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIIP7DZ0Z_0 ));
    Odrv4 I__11149 (
            .O(N__57108),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIIP7DZ0Z_0 ));
    LocalMux I__11148 (
            .O(N__57105),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIIP7DZ0Z_0 ));
    Odrv4 I__11147 (
            .O(N__57100),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIIP7DZ0Z_0 ));
    Odrv12 I__11146 (
            .O(N__57093),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIIP7DZ0Z_0 ));
    LocalMux I__11145 (
            .O(N__57086),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIIP7DZ0Z_0 ));
    InMux I__11144 (
            .O(N__57069),
            .I(N__57063));
    InMux I__11143 (
            .O(N__57068),
            .I(N__57060));
    InMux I__11142 (
            .O(N__57067),
            .I(N__57053));
    InMux I__11141 (
            .O(N__57066),
            .I(N__57048));
    LocalMux I__11140 (
            .O(N__57063),
            .I(N__57043));
    LocalMux I__11139 (
            .O(N__57060),
            .I(N__57043));
    InMux I__11138 (
            .O(N__57059),
            .I(N__57040));
    InMux I__11137 (
            .O(N__57058),
            .I(N__57034));
    InMux I__11136 (
            .O(N__57057),
            .I(N__57034));
    InMux I__11135 (
            .O(N__57056),
            .I(N__57031));
    LocalMux I__11134 (
            .O(N__57053),
            .I(N__57028));
    InMux I__11133 (
            .O(N__57052),
            .I(N__57022));
    InMux I__11132 (
            .O(N__57051),
            .I(N__57019));
    LocalMux I__11131 (
            .O(N__57048),
            .I(N__57016));
    Span4Mux_s3_v I__11130 (
            .O(N__57043),
            .I(N__57011));
    LocalMux I__11129 (
            .O(N__57040),
            .I(N__57011));
    InMux I__11128 (
            .O(N__57039),
            .I(N__57006));
    LocalMux I__11127 (
            .O(N__57034),
            .I(N__56999));
    LocalMux I__11126 (
            .O(N__57031),
            .I(N__56999));
    Span4Mux_h I__11125 (
            .O(N__57028),
            .I(N__56999));
    InMux I__11124 (
            .O(N__57027),
            .I(N__56994));
    InMux I__11123 (
            .O(N__57026),
            .I(N__56994));
    InMux I__11122 (
            .O(N__57025),
            .I(N__56991));
    LocalMux I__11121 (
            .O(N__57022),
            .I(N__56988));
    LocalMux I__11120 (
            .O(N__57019),
            .I(N__56981));
    Span4Mux_s3_v I__11119 (
            .O(N__57016),
            .I(N__56981));
    Span4Mux_h I__11118 (
            .O(N__57011),
            .I(N__56981));
    InMux I__11117 (
            .O(N__57010),
            .I(N__56978));
    InMux I__11116 (
            .O(N__57009),
            .I(N__56975));
    LocalMux I__11115 (
            .O(N__57006),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI5QE01Z0Z_3 ));
    Odrv4 I__11114 (
            .O(N__56999),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI5QE01Z0Z_3 ));
    LocalMux I__11113 (
            .O(N__56994),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI5QE01Z0Z_3 ));
    LocalMux I__11112 (
            .O(N__56991),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI5QE01Z0Z_3 ));
    Odrv4 I__11111 (
            .O(N__56988),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI5QE01Z0Z_3 ));
    Odrv4 I__11110 (
            .O(N__56981),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI5QE01Z0Z_3 ));
    LocalMux I__11109 (
            .O(N__56978),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI5QE01Z0Z_3 ));
    LocalMux I__11108 (
            .O(N__56975),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI5QE01Z0Z_3 ));
    InMux I__11107 (
            .O(N__56958),
            .I(N__56955));
    LocalMux I__11106 (
            .O(N__56955),
            .I(\ppm_encoder_1.un2_throttle_iv_0_1_2 ));
    CascadeMux I__11105 (
            .O(N__56952),
            .I(\ppm_encoder_1.un2_throttle_iv_0_2_2_cascade_ ));
    InMux I__11104 (
            .O(N__56949),
            .I(N__56941));
    InMux I__11103 (
            .O(N__56948),
            .I(N__56932));
    InMux I__11102 (
            .O(N__56947),
            .I(N__56929));
    InMux I__11101 (
            .O(N__56946),
            .I(N__56925));
    InMux I__11100 (
            .O(N__56945),
            .I(N__56921));
    InMux I__11099 (
            .O(N__56944),
            .I(N__56918));
    LocalMux I__11098 (
            .O(N__56941),
            .I(N__56915));
    InMux I__11097 (
            .O(N__56940),
            .I(N__56912));
    InMux I__11096 (
            .O(N__56939),
            .I(N__56909));
    InMux I__11095 (
            .O(N__56938),
            .I(N__56904));
    InMux I__11094 (
            .O(N__56937),
            .I(N__56904));
    InMux I__11093 (
            .O(N__56936),
            .I(N__56899));
    InMux I__11092 (
            .O(N__56935),
            .I(N__56899));
    LocalMux I__11091 (
            .O(N__56932),
            .I(N__56894));
    LocalMux I__11090 (
            .O(N__56929),
            .I(N__56894));
    InMux I__11089 (
            .O(N__56928),
            .I(N__56891));
    LocalMux I__11088 (
            .O(N__56925),
            .I(N__56888));
    InMux I__11087 (
            .O(N__56924),
            .I(N__56885));
    LocalMux I__11086 (
            .O(N__56921),
            .I(N__56882));
    LocalMux I__11085 (
            .O(N__56918),
            .I(N__56879));
    Span4Mux_s3_v I__11084 (
            .O(N__56915),
            .I(N__56876));
    LocalMux I__11083 (
            .O(N__56912),
            .I(N__56871));
    LocalMux I__11082 (
            .O(N__56909),
            .I(N__56871));
    LocalMux I__11081 (
            .O(N__56904),
            .I(N__56868));
    LocalMux I__11080 (
            .O(N__56899),
            .I(N__56865));
    Span4Mux_v I__11079 (
            .O(N__56894),
            .I(N__56856));
    LocalMux I__11078 (
            .O(N__56891),
            .I(N__56856));
    Span4Mux_h I__11077 (
            .O(N__56888),
            .I(N__56856));
    LocalMux I__11076 (
            .O(N__56885),
            .I(N__56853));
    Span4Mux_v I__11075 (
            .O(N__56882),
            .I(N__56846));
    Span4Mux_s3_v I__11074 (
            .O(N__56879),
            .I(N__56846));
    Span4Mux_h I__11073 (
            .O(N__56876),
            .I(N__56846));
    Span4Mux_v I__11072 (
            .O(N__56871),
            .I(N__56839));
    Span4Mux_s3_v I__11071 (
            .O(N__56868),
            .I(N__56839));
    Span4Mux_h I__11070 (
            .O(N__56865),
            .I(N__56839));
    InMux I__11069 (
            .O(N__56864),
            .I(N__56834));
    InMux I__11068 (
            .O(N__56863),
            .I(N__56834));
    Span4Mux_h I__11067 (
            .O(N__56856),
            .I(N__56829));
    Span4Mux_h I__11066 (
            .O(N__56853),
            .I(N__56829));
    Odrv4 I__11065 (
            .O(N__56846),
            .I(\ppm_encoder_1.PPM_STATE_RNI5C4LZ0Z_1 ));
    Odrv4 I__11064 (
            .O(N__56839),
            .I(\ppm_encoder_1.PPM_STATE_RNI5C4LZ0Z_1 ));
    LocalMux I__11063 (
            .O(N__56834),
            .I(\ppm_encoder_1.PPM_STATE_RNI5C4LZ0Z_1 ));
    Odrv4 I__11062 (
            .O(N__56829),
            .I(\ppm_encoder_1.PPM_STATE_RNI5C4LZ0Z_1 ));
    InMux I__11061 (
            .O(N__56820),
            .I(\ppm_encoder_1.counter24_0_N_2 ));
    InMux I__11060 (
            .O(N__56817),
            .I(N__56813));
    CascadeMux I__11059 (
            .O(N__56816),
            .I(N__56810));
    LocalMux I__11058 (
            .O(N__56813),
            .I(N__56807));
    InMux I__11057 (
            .O(N__56810),
            .I(N__56804));
    Span4Mux_v I__11056 (
            .O(N__56807),
            .I(N__56798));
    LocalMux I__11055 (
            .O(N__56804),
            .I(N__56798));
    InMux I__11054 (
            .O(N__56803),
            .I(N__56795));
    Span4Mux_h I__11053 (
            .O(N__56798),
            .I(N__56792));
    LocalMux I__11052 (
            .O(N__56795),
            .I(\ppm_encoder_1.aileronZ0Z_10 ));
    Odrv4 I__11051 (
            .O(N__56792),
            .I(\ppm_encoder_1.aileronZ0Z_10 ));
    InMux I__11050 (
            .O(N__56787),
            .I(N__56784));
    LocalMux I__11049 (
            .O(N__56784),
            .I(N__56781));
    Span4Mux_s3_v I__11048 (
            .O(N__56781),
            .I(N__56776));
    InMux I__11047 (
            .O(N__56780),
            .I(N__56773));
    CascadeMux I__11046 (
            .O(N__56779),
            .I(N__56770));
    Span4Mux_h I__11045 (
            .O(N__56776),
            .I(N__56765));
    LocalMux I__11044 (
            .O(N__56773),
            .I(N__56765));
    InMux I__11043 (
            .O(N__56770),
            .I(N__56762));
    Span4Mux_v I__11042 (
            .O(N__56765),
            .I(N__56759));
    LocalMux I__11041 (
            .O(N__56762),
            .I(\ppm_encoder_1.elevatorZ0Z_10 ));
    Odrv4 I__11040 (
            .O(N__56759),
            .I(\ppm_encoder_1.elevatorZ0Z_10 ));
    CascadeMux I__11039 (
            .O(N__56754),
            .I(N__56751));
    InMux I__11038 (
            .O(N__56751),
            .I(N__56748));
    LocalMux I__11037 (
            .O(N__56748),
            .I(\ppm_encoder_1.counter24_0_I_57_c_RNOZ0 ));
    CascadeMux I__11036 (
            .O(N__56745),
            .I(N__56742));
    InMux I__11035 (
            .O(N__56742),
            .I(N__56739));
    LocalMux I__11034 (
            .O(N__56739),
            .I(N__56736));
    Odrv12 I__11033 (
            .O(N__56736),
            .I(\ppm_encoder_1.N_258_i_i ));
    CascadeMux I__11032 (
            .O(N__56733),
            .I(\ppm_encoder_1.N_258_i_i_cascade_ ));
    InMux I__11031 (
            .O(N__56730),
            .I(N__56727));
    LocalMux I__11030 (
            .O(N__56727),
            .I(N__56724));
    Odrv12 I__11029 (
            .O(N__56724),
            .I(\ppm_encoder_1.init_pulses_RNI40GS4Z0Z_1 ));
    InMux I__11028 (
            .O(N__56721),
            .I(N__56716));
    InMux I__11027 (
            .O(N__56720),
            .I(N__56710));
    InMux I__11026 (
            .O(N__56719),
            .I(N__56710));
    LocalMux I__11025 (
            .O(N__56716),
            .I(N__56707));
    CascadeMux I__11024 (
            .O(N__56715),
            .I(N__56704));
    LocalMux I__11023 (
            .O(N__56710),
            .I(N__56701));
    Span4Mux_h I__11022 (
            .O(N__56707),
            .I(N__56698));
    InMux I__11021 (
            .O(N__56704),
            .I(N__56695));
    Span4Mux_v I__11020 (
            .O(N__56701),
            .I(N__56692));
    Odrv4 I__11019 (
            .O(N__56698),
            .I(\ppm_encoder_1.init_pulsesZ0Z_7 ));
    LocalMux I__11018 (
            .O(N__56695),
            .I(\ppm_encoder_1.init_pulsesZ0Z_7 ));
    Odrv4 I__11017 (
            .O(N__56692),
            .I(\ppm_encoder_1.init_pulsesZ0Z_7 ));
    CascadeMux I__11016 (
            .O(N__56685),
            .I(\ppm_encoder_1.PPM_STATE_RNI5C4LZ0Z_1_cascade_ ));
    InMux I__11015 (
            .O(N__56682),
            .I(N__56679));
    LocalMux I__11014 (
            .O(N__56679),
            .I(\ppm_encoder_1.aileron_RNIFUAPZ0Z_1 ));
    CascadeMux I__11013 (
            .O(N__56676),
            .I(\ppm_encoder_1.init_pulses_RNI7A1R_0Z0Z_1_cascade_ ));
    InMux I__11012 (
            .O(N__56673),
            .I(N__56670));
    LocalMux I__11011 (
            .O(N__56670),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_1 ));
    InMux I__11010 (
            .O(N__56667),
            .I(N__56663));
    InMux I__11009 (
            .O(N__56666),
            .I(N__56660));
    LocalMux I__11008 (
            .O(N__56663),
            .I(N__56657));
    LocalMux I__11007 (
            .O(N__56660),
            .I(N__56654));
    Span4Mux_v I__11006 (
            .O(N__56657),
            .I(N__56647));
    Span4Mux_v I__11005 (
            .O(N__56654),
            .I(N__56647));
    InMux I__11004 (
            .O(N__56653),
            .I(N__56644));
    InMux I__11003 (
            .O(N__56652),
            .I(N__56641));
    Span4Mux_v I__11002 (
            .O(N__56647),
            .I(N__56623));
    LocalMux I__11001 (
            .O(N__56644),
            .I(N__56623));
    LocalMux I__11000 (
            .O(N__56641),
            .I(N__56623));
    InMux I__10999 (
            .O(N__56640),
            .I(N__56620));
    InMux I__10998 (
            .O(N__56639),
            .I(N__56617));
    InMux I__10997 (
            .O(N__56638),
            .I(N__56614));
    CascadeMux I__10996 (
            .O(N__56637),
            .I(N__56611));
    CascadeMux I__10995 (
            .O(N__56636),
            .I(N__56608));
    CascadeMux I__10994 (
            .O(N__56635),
            .I(N__56605));
    CascadeMux I__10993 (
            .O(N__56634),
            .I(N__56602));
    CascadeMux I__10992 (
            .O(N__56633),
            .I(N__56599));
    CascadeMux I__10991 (
            .O(N__56632),
            .I(N__56596));
    CascadeMux I__10990 (
            .O(N__56631),
            .I(N__56591));
    InMux I__10989 (
            .O(N__56630),
            .I(N__56588));
    Span4Mux_v I__10988 (
            .O(N__56623),
            .I(N__56581));
    LocalMux I__10987 (
            .O(N__56620),
            .I(N__56581));
    LocalMux I__10986 (
            .O(N__56617),
            .I(N__56581));
    LocalMux I__10985 (
            .O(N__56614),
            .I(N__56577));
    InMux I__10984 (
            .O(N__56611),
            .I(N__56570));
    InMux I__10983 (
            .O(N__56608),
            .I(N__56570));
    InMux I__10982 (
            .O(N__56605),
            .I(N__56559));
    InMux I__10981 (
            .O(N__56602),
            .I(N__56559));
    InMux I__10980 (
            .O(N__56599),
            .I(N__56559));
    InMux I__10979 (
            .O(N__56596),
            .I(N__56559));
    InMux I__10978 (
            .O(N__56595),
            .I(N__56559));
    InMux I__10977 (
            .O(N__56594),
            .I(N__56554));
    InMux I__10976 (
            .O(N__56591),
            .I(N__56554));
    LocalMux I__10975 (
            .O(N__56588),
            .I(N__56543));
    Span4Mux_v I__10974 (
            .O(N__56581),
            .I(N__56540));
    InMux I__10973 (
            .O(N__56580),
            .I(N__56536));
    Span4Mux_v I__10972 (
            .O(N__56577),
            .I(N__56532));
    InMux I__10971 (
            .O(N__56576),
            .I(N__56529));
    CascadeMux I__10970 (
            .O(N__56575),
            .I(N__56525));
    LocalMux I__10969 (
            .O(N__56570),
            .I(N__56520));
    LocalMux I__10968 (
            .O(N__56559),
            .I(N__56515));
    LocalMux I__10967 (
            .O(N__56554),
            .I(N__56515));
    CascadeMux I__10966 (
            .O(N__56553),
            .I(N__56511));
    CascadeMux I__10965 (
            .O(N__56552),
            .I(N__56508));
    CascadeMux I__10964 (
            .O(N__56551),
            .I(N__56503));
    CascadeMux I__10963 (
            .O(N__56550),
            .I(N__56500));
    CascadeMux I__10962 (
            .O(N__56549),
            .I(N__56497));
    CascadeMux I__10961 (
            .O(N__56548),
            .I(N__56494));
    CascadeMux I__10960 (
            .O(N__56547),
            .I(N__56491));
    IoInMux I__10959 (
            .O(N__56546),
            .I(N__56488));
    Span4Mux_v I__10958 (
            .O(N__56543),
            .I(N__56485));
    Span4Mux_h I__10957 (
            .O(N__56540),
            .I(N__56480));
    InMux I__10956 (
            .O(N__56539),
            .I(N__56477));
    LocalMux I__10955 (
            .O(N__56536),
            .I(N__56474));
    InMux I__10954 (
            .O(N__56535),
            .I(N__56471));
    Span4Mux_v I__10953 (
            .O(N__56532),
            .I(N__56466));
    LocalMux I__10952 (
            .O(N__56529),
            .I(N__56466));
    InMux I__10951 (
            .O(N__56528),
            .I(N__56463));
    InMux I__10950 (
            .O(N__56525),
            .I(N__56460));
    CascadeMux I__10949 (
            .O(N__56524),
            .I(N__56456));
    CascadeMux I__10948 (
            .O(N__56523),
            .I(N__56453));
    Span4Mux_v I__10947 (
            .O(N__56520),
            .I(N__56448));
    Span4Mux_v I__10946 (
            .O(N__56515),
            .I(N__56448));
    InMux I__10945 (
            .O(N__56514),
            .I(N__56441));
    InMux I__10944 (
            .O(N__56511),
            .I(N__56441));
    InMux I__10943 (
            .O(N__56508),
            .I(N__56441));
    CascadeMux I__10942 (
            .O(N__56507),
            .I(N__56438));
    InMux I__10941 (
            .O(N__56506),
            .I(N__56435));
    InMux I__10940 (
            .O(N__56503),
            .I(N__56432));
    InMux I__10939 (
            .O(N__56500),
            .I(N__56429));
    InMux I__10938 (
            .O(N__56497),
            .I(N__56426));
    InMux I__10937 (
            .O(N__56494),
            .I(N__56421));
    InMux I__10936 (
            .O(N__56491),
            .I(N__56421));
    LocalMux I__10935 (
            .O(N__56488),
            .I(N__56418));
    Span4Mux_h I__10934 (
            .O(N__56485),
            .I(N__56415));
    InMux I__10933 (
            .O(N__56484),
            .I(N__56412));
    CascadeMux I__10932 (
            .O(N__56483),
            .I(N__56409));
    Span4Mux_h I__10931 (
            .O(N__56480),
            .I(N__56406));
    LocalMux I__10930 (
            .O(N__56477),
            .I(N__56403));
    Span4Mux_s1_h I__10929 (
            .O(N__56474),
            .I(N__56400));
    LocalMux I__10928 (
            .O(N__56471),
            .I(N__56397));
    Span4Mux_v I__10927 (
            .O(N__56466),
            .I(N__56392));
    LocalMux I__10926 (
            .O(N__56463),
            .I(N__56392));
    LocalMux I__10925 (
            .O(N__56460),
            .I(N__56389));
    InMux I__10924 (
            .O(N__56459),
            .I(N__56382));
    InMux I__10923 (
            .O(N__56456),
            .I(N__56382));
    InMux I__10922 (
            .O(N__56453),
            .I(N__56382));
    Span4Mux_v I__10921 (
            .O(N__56448),
            .I(N__56377));
    LocalMux I__10920 (
            .O(N__56441),
            .I(N__56377));
    InMux I__10919 (
            .O(N__56438),
            .I(N__56374));
    LocalMux I__10918 (
            .O(N__56435),
            .I(N__56371));
    LocalMux I__10917 (
            .O(N__56432),
            .I(N__56362));
    LocalMux I__10916 (
            .O(N__56429),
            .I(N__56362));
    LocalMux I__10915 (
            .O(N__56426),
            .I(N__56362));
    LocalMux I__10914 (
            .O(N__56421),
            .I(N__56362));
    Span12Mux_s8_v I__10913 (
            .O(N__56418),
            .I(N__56359));
    Sp12to4 I__10912 (
            .O(N__56415),
            .I(N__56354));
    LocalMux I__10911 (
            .O(N__56412),
            .I(N__56354));
    InMux I__10910 (
            .O(N__56409),
            .I(N__56351));
    Span4Mux_h I__10909 (
            .O(N__56406),
            .I(N__56348));
    Span4Mux_v I__10908 (
            .O(N__56403),
            .I(N__56339));
    Span4Mux_v I__10907 (
            .O(N__56400),
            .I(N__56339));
    Span4Mux_v I__10906 (
            .O(N__56397),
            .I(N__56339));
    Span4Mux_v I__10905 (
            .O(N__56392),
            .I(N__56339));
    Span4Mux_h I__10904 (
            .O(N__56389),
            .I(N__56334));
    LocalMux I__10903 (
            .O(N__56382),
            .I(N__56334));
    Span4Mux_h I__10902 (
            .O(N__56377),
            .I(N__56329));
    LocalMux I__10901 (
            .O(N__56374),
            .I(N__56329));
    Span12Mux_s7_h I__10900 (
            .O(N__56371),
            .I(N__56326));
    Span4Mux_v I__10899 (
            .O(N__56362),
            .I(N__56323));
    Span12Mux_v I__10898 (
            .O(N__56359),
            .I(N__56316));
    Span12Mux_v I__10897 (
            .O(N__56354),
            .I(N__56316));
    LocalMux I__10896 (
            .O(N__56351),
            .I(N__56316));
    Span4Mux_h I__10895 (
            .O(N__56348),
            .I(N__56309));
    Span4Mux_h I__10894 (
            .O(N__56339),
            .I(N__56309));
    Span4Mux_v I__10893 (
            .O(N__56334),
            .I(N__56309));
    Span4Mux_h I__10892 (
            .O(N__56329),
            .I(N__56306));
    Odrv12 I__10891 (
            .O(N__56326),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__10890 (
            .O(N__56323),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__10889 (
            .O(N__56316),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__10888 (
            .O(N__56309),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__10887 (
            .O(N__56306),
            .I(CONSTANT_ONE_NET));
    InMux I__10886 (
            .O(N__56295),
            .I(N__56292));
    LocalMux I__10885 (
            .O(N__56292),
            .I(N__56288));
    InMux I__10884 (
            .O(N__56291),
            .I(N__56285));
    Span4Mux_h I__10883 (
            .O(N__56288),
            .I(N__56280));
    LocalMux I__10882 (
            .O(N__56285),
            .I(N__56280));
    Span4Mux_v I__10881 (
            .O(N__56280),
            .I(N__56276));
    InMux I__10880 (
            .O(N__56279),
            .I(N__56273));
    Span4Mux_h I__10879 (
            .O(N__56276),
            .I(N__56270));
    LocalMux I__10878 (
            .O(N__56273),
            .I(\pid_front.error_i_reg_esr_RNI8KHVZ0Z_25 ));
    Odrv4 I__10877 (
            .O(N__56270),
            .I(\pid_front.error_i_reg_esr_RNI8KHVZ0Z_25 ));
    CascadeMux I__10876 (
            .O(N__56265),
            .I(N__56261));
    InMux I__10875 (
            .O(N__56264),
            .I(N__56256));
    InMux I__10874 (
            .O(N__56261),
            .I(N__56256));
    LocalMux I__10873 (
            .O(N__56256),
            .I(\pid_front.error_i_acumm_preregZ0Z_25 ));
    InMux I__10872 (
            .O(N__56253),
            .I(N__56248));
    InMux I__10871 (
            .O(N__56252),
            .I(N__56245));
    InMux I__10870 (
            .O(N__56251),
            .I(N__56242));
    LocalMux I__10869 (
            .O(N__56248),
            .I(N__56239));
    LocalMux I__10868 (
            .O(N__56245),
            .I(N__56236));
    LocalMux I__10867 (
            .O(N__56242),
            .I(N__56233));
    Span12Mux_v I__10866 (
            .O(N__56239),
            .I(N__56230));
    Span4Mux_h I__10865 (
            .O(N__56236),
            .I(N__56227));
    Odrv4 I__10864 (
            .O(N__56233),
            .I(\pid_front.error_i_reg_esr_RNI4EFVZ0Z_23 ));
    Odrv12 I__10863 (
            .O(N__56230),
            .I(\pid_front.error_i_reg_esr_RNI4EFVZ0Z_23 ));
    Odrv4 I__10862 (
            .O(N__56227),
            .I(\pid_front.error_i_reg_esr_RNI4EFVZ0Z_23 ));
    InMux I__10861 (
            .O(N__56220),
            .I(N__56214));
    InMux I__10860 (
            .O(N__56219),
            .I(N__56214));
    LocalMux I__10859 (
            .O(N__56214),
            .I(\pid_front.error_i_acumm_preregZ0Z_23 ));
    InMux I__10858 (
            .O(N__56211),
            .I(N__56205));
    InMux I__10857 (
            .O(N__56210),
            .I(N__56205));
    LocalMux I__10856 (
            .O(N__56205),
            .I(N__56202));
    Span4Mux_h I__10855 (
            .O(N__56202),
            .I(N__56199));
    Span4Mux_v I__10854 (
            .O(N__56199),
            .I(N__56195));
    InMux I__10853 (
            .O(N__56198),
            .I(N__56192));
    Span4Mux_h I__10852 (
            .O(N__56195),
            .I(N__56189));
    LocalMux I__10851 (
            .O(N__56192),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_26_c_RNICQJV ));
    Odrv4 I__10850 (
            .O(N__56189),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_26_c_RNICQJV ));
    InMux I__10849 (
            .O(N__56184),
            .I(N__56178));
    InMux I__10848 (
            .O(N__56183),
            .I(N__56178));
    LocalMux I__10847 (
            .O(N__56178),
            .I(\pid_front.error_i_acumm_preregZ0Z_27 ));
    InMux I__10846 (
            .O(N__56175),
            .I(N__56170));
    InMux I__10845 (
            .O(N__56174),
            .I(N__56165));
    InMux I__10844 (
            .O(N__56173),
            .I(N__56165));
    LocalMux I__10843 (
            .O(N__56170),
            .I(N__56162));
    LocalMux I__10842 (
            .O(N__56165),
            .I(N__56159));
    Odrv4 I__10841 (
            .O(N__56162),
            .I(\pid_front.error_i_reg_esr_RNIALFUZ0Z_17 ));
    Odrv12 I__10840 (
            .O(N__56159),
            .I(\pid_front.error_i_reg_esr_RNIALFUZ0Z_17 ));
    CascadeMux I__10839 (
            .O(N__56154),
            .I(N__56150));
    InMux I__10838 (
            .O(N__56153),
            .I(N__56145));
    InMux I__10837 (
            .O(N__56150),
            .I(N__56145));
    LocalMux I__10836 (
            .O(N__56145),
            .I(N__56142));
    Odrv4 I__10835 (
            .O(N__56142),
            .I(\pid_front.error_i_acumm_preregZ0Z_17 ));
    InMux I__10834 (
            .O(N__56139),
            .I(N__56136));
    LocalMux I__10833 (
            .O(N__56136),
            .I(N__56133));
    Span4Mux_s3_v I__10832 (
            .O(N__56133),
            .I(N__56130));
    Span4Mux_v I__10831 (
            .O(N__56130),
            .I(N__56126));
    InMux I__10830 (
            .O(N__56129),
            .I(N__56123));
    Odrv4 I__10829 (
            .O(N__56126),
            .I(\pid_front.error_i_acummZ0Z_0 ));
    LocalMux I__10828 (
            .O(N__56123),
            .I(\pid_front.error_i_acummZ0Z_0 ));
    InMux I__10827 (
            .O(N__56118),
            .I(N__56114));
    InMux I__10826 (
            .O(N__56117),
            .I(N__56111));
    LocalMux I__10825 (
            .O(N__56114),
            .I(N__56108));
    LocalMux I__10824 (
            .O(N__56111),
            .I(N__56105));
    Span4Mux_v I__10823 (
            .O(N__56108),
            .I(N__56100));
    Span4Mux_h I__10822 (
            .O(N__56105),
            .I(N__56100));
    Span4Mux_v I__10821 (
            .O(N__56100),
            .I(N__56097));
    Odrv4 I__10820 (
            .O(N__56097),
            .I(\pid_front.error_i_acumm_preregZ0Z_0 ));
    InMux I__10819 (
            .O(N__56094),
            .I(N__56088));
    InMux I__10818 (
            .O(N__56093),
            .I(N__56088));
    LocalMux I__10817 (
            .O(N__56088),
            .I(N__56072));
    CEMux I__10816 (
            .O(N__56087),
            .I(N__56043));
    CEMux I__10815 (
            .O(N__56086),
            .I(N__56043));
    CEMux I__10814 (
            .O(N__56085),
            .I(N__56043));
    CEMux I__10813 (
            .O(N__56084),
            .I(N__56043));
    CEMux I__10812 (
            .O(N__56083),
            .I(N__56043));
    CEMux I__10811 (
            .O(N__56082),
            .I(N__56043));
    CEMux I__10810 (
            .O(N__56081),
            .I(N__56043));
    CEMux I__10809 (
            .O(N__56080),
            .I(N__56043));
    CEMux I__10808 (
            .O(N__56079),
            .I(N__56043));
    CEMux I__10807 (
            .O(N__56078),
            .I(N__56043));
    CEMux I__10806 (
            .O(N__56077),
            .I(N__56043));
    CEMux I__10805 (
            .O(N__56076),
            .I(N__56043));
    CEMux I__10804 (
            .O(N__56075),
            .I(N__56043));
    Glb2LocalMux I__10803 (
            .O(N__56072),
            .I(N__56043));
    GlobalMux I__10802 (
            .O(N__56043),
            .I(N__56040));
    gio2CtrlBuf I__10801 (
            .O(N__56040),
            .I(\pid_front.N_764_g ));
    InMux I__10800 (
            .O(N__56037),
            .I(N__56034));
    LocalMux I__10799 (
            .O(N__56034),
            .I(N__56031));
    Span4Mux_v I__10798 (
            .O(N__56031),
            .I(N__56027));
    InMux I__10797 (
            .O(N__56030),
            .I(N__56024));
    Span4Mux_v I__10796 (
            .O(N__56027),
            .I(N__56021));
    LocalMux I__10795 (
            .O(N__56024),
            .I(N__56015));
    Span4Mux_v I__10794 (
            .O(N__56021),
            .I(N__56012));
    CascadeMux I__10793 (
            .O(N__56020),
            .I(N__56009));
    InMux I__10792 (
            .O(N__56019),
            .I(N__56004));
    InMux I__10791 (
            .O(N__56018),
            .I(N__56004));
    Span4Mux_v I__10790 (
            .O(N__56015),
            .I(N__55999));
    Span4Mux_v I__10789 (
            .O(N__56012),
            .I(N__55999));
    InMux I__10788 (
            .O(N__56009),
            .I(N__55996));
    LocalMux I__10787 (
            .O(N__56004),
            .I(\pid_alt.stateZ0Z_0 ));
    Odrv4 I__10786 (
            .O(N__55999),
            .I(\pid_alt.stateZ0Z_0 ));
    LocalMux I__10785 (
            .O(N__55996),
            .I(\pid_alt.stateZ0Z_0 ));
    IoInMux I__10784 (
            .O(N__55989),
            .I(N__55986));
    LocalMux I__10783 (
            .O(N__55986),
            .I(N__55983));
    Odrv4 I__10782 (
            .O(N__55983),
            .I(\pid_alt.state_0_0 ));
    InMux I__10781 (
            .O(N__55980),
            .I(N__55977));
    LocalMux I__10780 (
            .O(N__55977),
            .I(N__55974));
    Sp12to4 I__10779 (
            .O(N__55974),
            .I(N__55971));
    Span12Mux_s10_v I__10778 (
            .O(N__55971),
            .I(N__55968));
    Odrv12 I__10777 (
            .O(N__55968),
            .I(\ppm_encoder_1.un1_init_pulses_11_0 ));
    InMux I__10776 (
            .O(N__55965),
            .I(N__55962));
    LocalMux I__10775 (
            .O(N__55962),
            .I(N__55959));
    Odrv4 I__10774 (
            .O(N__55959),
            .I(\ppm_encoder_1.un1_init_pulses_10_0 ));
    CascadeMux I__10773 (
            .O(N__55956),
            .I(N__55948));
    CascadeMux I__10772 (
            .O(N__55955),
            .I(N__55945));
    CascadeMux I__10771 (
            .O(N__55954),
            .I(N__55933));
    CascadeMux I__10770 (
            .O(N__55953),
            .I(N__55930));
    CascadeMux I__10769 (
            .O(N__55952),
            .I(N__55927));
    CascadeMux I__10768 (
            .O(N__55951),
            .I(N__55924));
    InMux I__10767 (
            .O(N__55948),
            .I(N__55909));
    InMux I__10766 (
            .O(N__55945),
            .I(N__55909));
    InMux I__10765 (
            .O(N__55944),
            .I(N__55909));
    InMux I__10764 (
            .O(N__55943),
            .I(N__55909));
    InMux I__10763 (
            .O(N__55942),
            .I(N__55909));
    InMux I__10762 (
            .O(N__55941),
            .I(N__55909));
    InMux I__10761 (
            .O(N__55940),
            .I(N__55909));
    CascadeMux I__10760 (
            .O(N__55939),
            .I(N__55905));
    CascadeMux I__10759 (
            .O(N__55938),
            .I(N__55902));
    CascadeMux I__10758 (
            .O(N__55937),
            .I(N__55899));
    CascadeMux I__10757 (
            .O(N__55936),
            .I(N__55896));
    InMux I__10756 (
            .O(N__55933),
            .I(N__55891));
    InMux I__10755 (
            .O(N__55930),
            .I(N__55886));
    InMux I__10754 (
            .O(N__55927),
            .I(N__55886));
    InMux I__10753 (
            .O(N__55924),
            .I(N__55883));
    LocalMux I__10752 (
            .O(N__55909),
            .I(N__55880));
    CascadeMux I__10751 (
            .O(N__55908),
            .I(N__55877));
    InMux I__10750 (
            .O(N__55905),
            .I(N__55873));
    InMux I__10749 (
            .O(N__55902),
            .I(N__55862));
    InMux I__10748 (
            .O(N__55899),
            .I(N__55862));
    InMux I__10747 (
            .O(N__55896),
            .I(N__55862));
    InMux I__10746 (
            .O(N__55895),
            .I(N__55862));
    InMux I__10745 (
            .O(N__55894),
            .I(N__55862));
    LocalMux I__10744 (
            .O(N__55891),
            .I(N__55859));
    LocalMux I__10743 (
            .O(N__55886),
            .I(N__55854));
    LocalMux I__10742 (
            .O(N__55883),
            .I(N__55854));
    Span4Mux_v I__10741 (
            .O(N__55880),
            .I(N__55851));
    InMux I__10740 (
            .O(N__55877),
            .I(N__55846));
    InMux I__10739 (
            .O(N__55876),
            .I(N__55846));
    LocalMux I__10738 (
            .O(N__55873),
            .I(N__55841));
    LocalMux I__10737 (
            .O(N__55862),
            .I(N__55841));
    Span4Mux_h I__10736 (
            .O(N__55859),
            .I(N__55834));
    Span4Mux_h I__10735 (
            .O(N__55854),
            .I(N__55834));
    Span4Mux_s0_v I__10734 (
            .O(N__55851),
            .I(N__55834));
    LocalMux I__10733 (
            .O(N__55846),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_RNIB7481Z0Z_3 ));
    Odrv4 I__10732 (
            .O(N__55841),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_RNIB7481Z0Z_3 ));
    Odrv4 I__10731 (
            .O(N__55834),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_RNIB7481Z0Z_3 ));
    InMux I__10730 (
            .O(N__55827),
            .I(N__55824));
    LocalMux I__10729 (
            .O(N__55824),
            .I(N__55819));
    InMux I__10728 (
            .O(N__55823),
            .I(N__55814));
    InMux I__10727 (
            .O(N__55822),
            .I(N__55814));
    Span4Mux_s1_v I__10726 (
            .O(N__55819),
            .I(N__55809));
    LocalMux I__10725 (
            .O(N__55814),
            .I(N__55809));
    Span4Mux_h I__10724 (
            .O(N__55809),
            .I(N__55800));
    InMux I__10723 (
            .O(N__55808),
            .I(N__55797));
    InMux I__10722 (
            .O(N__55807),
            .I(N__55792));
    InMux I__10721 (
            .O(N__55806),
            .I(N__55792));
    CascadeMux I__10720 (
            .O(N__55805),
            .I(N__55788));
    CascadeMux I__10719 (
            .O(N__55804),
            .I(N__55784));
    CascadeMux I__10718 (
            .O(N__55803),
            .I(N__55777));
    Span4Mux_s1_v I__10717 (
            .O(N__55800),
            .I(N__55770));
    LocalMux I__10716 (
            .O(N__55797),
            .I(N__55765));
    LocalMux I__10715 (
            .O(N__55792),
            .I(N__55765));
    InMux I__10714 (
            .O(N__55791),
            .I(N__55752));
    InMux I__10713 (
            .O(N__55788),
            .I(N__55752));
    InMux I__10712 (
            .O(N__55787),
            .I(N__55752));
    InMux I__10711 (
            .O(N__55784),
            .I(N__55752));
    InMux I__10710 (
            .O(N__55783),
            .I(N__55752));
    InMux I__10709 (
            .O(N__55782),
            .I(N__55752));
    InMux I__10708 (
            .O(N__55781),
            .I(N__55737));
    InMux I__10707 (
            .O(N__55780),
            .I(N__55737));
    InMux I__10706 (
            .O(N__55777),
            .I(N__55737));
    InMux I__10705 (
            .O(N__55776),
            .I(N__55737));
    InMux I__10704 (
            .O(N__55775),
            .I(N__55737));
    InMux I__10703 (
            .O(N__55774),
            .I(N__55737));
    InMux I__10702 (
            .O(N__55773),
            .I(N__55737));
    Odrv4 I__10701 (
            .O(N__55770),
            .I(\ppm_encoder_1.counter24_0_I_57_c_RNIV9SJZ0Z1 ));
    Odrv4 I__10700 (
            .O(N__55765),
            .I(\ppm_encoder_1.counter24_0_I_57_c_RNIV9SJZ0Z1 ));
    LocalMux I__10699 (
            .O(N__55752),
            .I(\ppm_encoder_1.counter24_0_I_57_c_RNIV9SJZ0Z1 ));
    LocalMux I__10698 (
            .O(N__55737),
            .I(\ppm_encoder_1.counter24_0_I_57_c_RNIV9SJZ0Z1 ));
    InMux I__10697 (
            .O(N__55728),
            .I(N__55725));
    LocalMux I__10696 (
            .O(N__55725),
            .I(N__55721));
    InMux I__10695 (
            .O(N__55724),
            .I(N__55718));
    Span4Mux_h I__10694 (
            .O(N__55721),
            .I(N__55713));
    LocalMux I__10693 (
            .O(N__55718),
            .I(N__55713));
    Span4Mux_h I__10692 (
            .O(N__55713),
            .I(N__55709));
    InMux I__10691 (
            .O(N__55712),
            .I(N__55706));
    Span4Mux_v I__10690 (
            .O(N__55709),
            .I(N__55703));
    LocalMux I__10689 (
            .O(N__55706),
            .I(\pid_front.error_i_reg_esr_RNI08DVZ0Z_21 ));
    Odrv4 I__10688 (
            .O(N__55703),
            .I(\pid_front.error_i_reg_esr_RNI08DVZ0Z_21 ));
    InMux I__10687 (
            .O(N__55698),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_20 ));
    InMux I__10686 (
            .O(N__55695),
            .I(N__55689));
    InMux I__10685 (
            .O(N__55694),
            .I(N__55689));
    LocalMux I__10684 (
            .O(N__55689),
            .I(N__55686));
    Span4Mux_h I__10683 (
            .O(N__55686),
            .I(N__55682));
    InMux I__10682 (
            .O(N__55685),
            .I(N__55679));
    Span4Mux_v I__10681 (
            .O(N__55682),
            .I(N__55676));
    LocalMux I__10680 (
            .O(N__55679),
            .I(\pid_front.error_i_reg_esr_RNI2BEVZ0Z_22 ));
    Odrv4 I__10679 (
            .O(N__55676),
            .I(\pid_front.error_i_reg_esr_RNI2BEVZ0Z_22 ));
    InMux I__10678 (
            .O(N__55671),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_21 ));
    InMux I__10677 (
            .O(N__55668),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_22 ));
    InMux I__10676 (
            .O(N__55665),
            .I(N__55659));
    InMux I__10675 (
            .O(N__55664),
            .I(N__55659));
    LocalMux I__10674 (
            .O(N__55659),
            .I(N__55656));
    Span4Mux_v I__10673 (
            .O(N__55656),
            .I(N__55652));
    InMux I__10672 (
            .O(N__55655),
            .I(N__55649));
    Span4Mux_h I__10671 (
            .O(N__55652),
            .I(N__55646));
    LocalMux I__10670 (
            .O(N__55649),
            .I(\pid_front.error_i_reg_esr_RNI6HGVZ0Z_24 ));
    Odrv4 I__10669 (
            .O(N__55646),
            .I(\pid_front.error_i_reg_esr_RNI6HGVZ0Z_24 ));
    InMux I__10668 (
            .O(N__55641),
            .I(bfn_13_26_0_));
    InMux I__10667 (
            .O(N__55638),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_24 ));
    InMux I__10666 (
            .O(N__55635),
            .I(N__55629));
    InMux I__10665 (
            .O(N__55634),
            .I(N__55629));
    LocalMux I__10664 (
            .O(N__55629),
            .I(N__55626));
    Span4Mux_v I__10663 (
            .O(N__55626),
            .I(N__55622));
    InMux I__10662 (
            .O(N__55625),
            .I(N__55619));
    Span4Mux_h I__10661 (
            .O(N__55622),
            .I(N__55616));
    LocalMux I__10660 (
            .O(N__55619),
            .I(\pid_front.error_i_reg_esr_RNIANIVZ0Z_26 ));
    Odrv4 I__10659 (
            .O(N__55616),
            .I(\pid_front.error_i_reg_esr_RNIANIVZ0Z_26 ));
    InMux I__10658 (
            .O(N__55611),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_25 ));
    InMux I__10657 (
            .O(N__55608),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_26 ));
    CascadeMux I__10656 (
            .O(N__55605),
            .I(N__55600));
    CascadeMux I__10655 (
            .O(N__55604),
            .I(N__55596));
    InMux I__10654 (
            .O(N__55603),
            .I(N__55579));
    InMux I__10653 (
            .O(N__55600),
            .I(N__55579));
    InMux I__10652 (
            .O(N__55599),
            .I(N__55579));
    InMux I__10651 (
            .O(N__55596),
            .I(N__55579));
    InMux I__10650 (
            .O(N__55595),
            .I(N__55579));
    CascadeMux I__10649 (
            .O(N__55594),
            .I(N__55576));
    CascadeMux I__10648 (
            .O(N__55593),
            .I(N__55572));
    CascadeMux I__10647 (
            .O(N__55592),
            .I(N__55568));
    CascadeMux I__10646 (
            .O(N__55591),
            .I(N__55564));
    CascadeMux I__10645 (
            .O(N__55590),
            .I(N__55559));
    LocalMux I__10644 (
            .O(N__55579),
            .I(N__55555));
    InMux I__10643 (
            .O(N__55576),
            .I(N__55538));
    InMux I__10642 (
            .O(N__55575),
            .I(N__55538));
    InMux I__10641 (
            .O(N__55572),
            .I(N__55538));
    InMux I__10640 (
            .O(N__55571),
            .I(N__55538));
    InMux I__10639 (
            .O(N__55568),
            .I(N__55538));
    InMux I__10638 (
            .O(N__55567),
            .I(N__55538));
    InMux I__10637 (
            .O(N__55564),
            .I(N__55538));
    InMux I__10636 (
            .O(N__55563),
            .I(N__55538));
    InMux I__10635 (
            .O(N__55562),
            .I(N__55531));
    InMux I__10634 (
            .O(N__55559),
            .I(N__55531));
    InMux I__10633 (
            .O(N__55558),
            .I(N__55531));
    Odrv4 I__10632 (
            .O(N__55555),
            .I(\pid_front.error_i_acummZ0Z_13 ));
    LocalMux I__10631 (
            .O(N__55538),
            .I(\pid_front.error_i_acummZ0Z_13 ));
    LocalMux I__10630 (
            .O(N__55531),
            .I(\pid_front.error_i_acummZ0Z_13 ));
    InMux I__10629 (
            .O(N__55524),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_27 ));
    InMux I__10628 (
            .O(N__55521),
            .I(N__55515));
    InMux I__10627 (
            .O(N__55520),
            .I(N__55515));
    LocalMux I__10626 (
            .O(N__55515),
            .I(N__55512));
    Span4Mux_v I__10625 (
            .O(N__55512),
            .I(N__55508));
    InMux I__10624 (
            .O(N__55511),
            .I(N__55505));
    Span4Mux_h I__10623 (
            .O(N__55508),
            .I(N__55502));
    LocalMux I__10622 (
            .O(N__55505),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_27_c_RNIDSKV ));
    Odrv4 I__10621 (
            .O(N__55502),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_27_c_RNIDSKV ));
    InMux I__10620 (
            .O(N__55497),
            .I(N__55493));
    CascadeMux I__10619 (
            .O(N__55496),
            .I(N__55489));
    LocalMux I__10618 (
            .O(N__55493),
            .I(N__55486));
    InMux I__10617 (
            .O(N__55492),
            .I(N__55481));
    InMux I__10616 (
            .O(N__55489),
            .I(N__55481));
    Span4Mux_h I__10615 (
            .O(N__55486),
            .I(N__55478));
    LocalMux I__10614 (
            .O(N__55481),
            .I(N__55475));
    Span4Mux_v I__10613 (
            .O(N__55478),
            .I(N__55472));
    Span4Mux_h I__10612 (
            .O(N__55475),
            .I(N__55469));
    Odrv4 I__10611 (
            .O(N__55472),
            .I(\pid_front.error_i_acumm_preregZ0Z_28 ));
    Odrv4 I__10610 (
            .O(N__55469),
            .I(\pid_front.error_i_acumm_preregZ0Z_28 ));
    InMux I__10609 (
            .O(N__55464),
            .I(N__55461));
    LocalMux I__10608 (
            .O(N__55461),
            .I(N__55455));
    InMux I__10607 (
            .O(N__55460),
            .I(N__55452));
    InMux I__10606 (
            .O(N__55459),
            .I(N__55449));
    InMux I__10605 (
            .O(N__55458),
            .I(N__55446));
    Span4Mux_h I__10604 (
            .O(N__55455),
            .I(N__55441));
    LocalMux I__10603 (
            .O(N__55452),
            .I(N__55441));
    LocalMux I__10602 (
            .O(N__55449),
            .I(N__55438));
    LocalMux I__10601 (
            .O(N__55446),
            .I(N__55435));
    Span4Mux_v I__10600 (
            .O(N__55441),
            .I(N__55432));
    Sp12to4 I__10599 (
            .O(N__55438),
            .I(N__55429));
    Odrv4 I__10598 (
            .O(N__55435),
            .I(\pid_front.error_i_reg_esr_RNI29BUZ0Z_13 ));
    Odrv4 I__10597 (
            .O(N__55432),
            .I(\pid_front.error_i_reg_esr_RNI29BUZ0Z_13 ));
    Odrv12 I__10596 (
            .O(N__55429),
            .I(\pid_front.error_i_reg_esr_RNI29BUZ0Z_13 ));
    InMux I__10595 (
            .O(N__55422),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_12 ));
    InMux I__10594 (
            .O(N__55419),
            .I(N__55415));
    InMux I__10593 (
            .O(N__55418),
            .I(N__55411));
    LocalMux I__10592 (
            .O(N__55415),
            .I(N__55408));
    InMux I__10591 (
            .O(N__55414),
            .I(N__55405));
    LocalMux I__10590 (
            .O(N__55411),
            .I(N__55402));
    Span4Mux_h I__10589 (
            .O(N__55408),
            .I(N__55399));
    LocalMux I__10588 (
            .O(N__55405),
            .I(N__55396));
    Span4Mux_v I__10587 (
            .O(N__55402),
            .I(N__55391));
    Span4Mux_v I__10586 (
            .O(N__55399),
            .I(N__55391));
    Span4Mux_h I__10585 (
            .O(N__55396),
            .I(N__55388));
    Odrv4 I__10584 (
            .O(N__55391),
            .I(\pid_front.error_i_reg_esr_RNI4CCUZ0Z_14 ));
    Odrv4 I__10583 (
            .O(N__55388),
            .I(\pid_front.error_i_reg_esr_RNI4CCUZ0Z_14 ));
    InMux I__10582 (
            .O(N__55383),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_13 ));
    InMux I__10581 (
            .O(N__55380),
            .I(N__55375));
    InMux I__10580 (
            .O(N__55379),
            .I(N__55370));
    InMux I__10579 (
            .O(N__55378),
            .I(N__55370));
    LocalMux I__10578 (
            .O(N__55375),
            .I(N__55367));
    LocalMux I__10577 (
            .O(N__55370),
            .I(N__55364));
    Span4Mux_h I__10576 (
            .O(N__55367),
            .I(N__55361));
    Span4Mux_h I__10575 (
            .O(N__55364),
            .I(N__55358));
    Odrv4 I__10574 (
            .O(N__55361),
            .I(\pid_front.error_i_reg_esr_RNI6FDUZ0Z_15 ));
    Odrv4 I__10573 (
            .O(N__55358),
            .I(\pid_front.error_i_reg_esr_RNI6FDUZ0Z_15 ));
    InMux I__10572 (
            .O(N__55353),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_14 ));
    InMux I__10571 (
            .O(N__55350),
            .I(N__55347));
    LocalMux I__10570 (
            .O(N__55347),
            .I(N__55342));
    InMux I__10569 (
            .O(N__55346),
            .I(N__55339));
    InMux I__10568 (
            .O(N__55345),
            .I(N__55336));
    Span12Mux_v I__10567 (
            .O(N__55342),
            .I(N__55331));
    LocalMux I__10566 (
            .O(N__55339),
            .I(N__55331));
    LocalMux I__10565 (
            .O(N__55336),
            .I(\pid_front.error_i_reg_esr_RNI8IEUZ0Z_16 ));
    Odrv12 I__10564 (
            .O(N__55331),
            .I(\pid_front.error_i_reg_esr_RNI8IEUZ0Z_16 ));
    InMux I__10563 (
            .O(N__55326),
            .I(bfn_13_25_0_));
    InMux I__10562 (
            .O(N__55323),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_16 ));
    InMux I__10561 (
            .O(N__55320),
            .I(N__55316));
    InMux I__10560 (
            .O(N__55319),
            .I(N__55313));
    LocalMux I__10559 (
            .O(N__55316),
            .I(N__55309));
    LocalMux I__10558 (
            .O(N__55313),
            .I(N__55306));
    InMux I__10557 (
            .O(N__55312),
            .I(N__55303));
    Span4Mux_h I__10556 (
            .O(N__55309),
            .I(N__55298));
    Span4Mux_v I__10555 (
            .O(N__55306),
            .I(N__55298));
    LocalMux I__10554 (
            .O(N__55303),
            .I(N__55295));
    Odrv4 I__10553 (
            .O(N__55298),
            .I(\pid_front.error_i_reg_esr_RNICOGUZ0Z_18 ));
    Odrv12 I__10552 (
            .O(N__55295),
            .I(\pid_front.error_i_reg_esr_RNICOGUZ0Z_18 ));
    InMux I__10551 (
            .O(N__55290),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_17 ));
    InMux I__10550 (
            .O(N__55287),
            .I(N__55283));
    InMux I__10549 (
            .O(N__55286),
            .I(N__55279));
    LocalMux I__10548 (
            .O(N__55283),
            .I(N__55276));
    InMux I__10547 (
            .O(N__55282),
            .I(N__55273));
    LocalMux I__10546 (
            .O(N__55279),
            .I(N__55270));
    Span4Mux_v I__10545 (
            .O(N__55276),
            .I(N__55267));
    LocalMux I__10544 (
            .O(N__55273),
            .I(N__55264));
    Span4Mux_h I__10543 (
            .O(N__55270),
            .I(N__55257));
    Span4Mux_h I__10542 (
            .O(N__55267),
            .I(N__55257));
    Span4Mux_v I__10541 (
            .O(N__55264),
            .I(N__55257));
    Odrv4 I__10540 (
            .O(N__55257),
            .I(\pid_front.error_i_reg_esr_RNIERHUZ0Z_19 ));
    InMux I__10539 (
            .O(N__55254),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_18 ));
    InMux I__10538 (
            .O(N__55251),
            .I(N__55245));
    InMux I__10537 (
            .O(N__55250),
            .I(N__55245));
    LocalMux I__10536 (
            .O(N__55245),
            .I(N__55242));
    Span4Mux_v I__10535 (
            .O(N__55242),
            .I(N__55238));
    InMux I__10534 (
            .O(N__55241),
            .I(N__55235));
    Span4Mux_h I__10533 (
            .O(N__55238),
            .I(N__55232));
    LocalMux I__10532 (
            .O(N__55235),
            .I(\pid_front.error_i_reg_esr_RNI7MJUZ0Z_20 ));
    Odrv4 I__10531 (
            .O(N__55232),
            .I(\pid_front.error_i_reg_esr_RNI7MJUZ0Z_20 ));
    InMux I__10530 (
            .O(N__55227),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_19 ));
    InMux I__10529 (
            .O(N__55224),
            .I(N__55221));
    LocalMux I__10528 (
            .O(N__55221),
            .I(\pid_front.error_i_acummZ0Z_5 ));
    CascadeMux I__10527 (
            .O(N__55218),
            .I(N__55215));
    InMux I__10526 (
            .O(N__55215),
            .I(N__55212));
    LocalMux I__10525 (
            .O(N__55212),
            .I(N__55208));
    InMux I__10524 (
            .O(N__55211),
            .I(N__55205));
    Span4Mux_h I__10523 (
            .O(N__55208),
            .I(N__55202));
    LocalMux I__10522 (
            .O(N__55205),
            .I(\pid_front.error_i_regZ0Z_5 ));
    Odrv4 I__10521 (
            .O(N__55202),
            .I(\pid_front.error_i_regZ0Z_5 ));
    InMux I__10520 (
            .O(N__55197),
            .I(N__55191));
    InMux I__10519 (
            .O(N__55196),
            .I(N__55186));
    InMux I__10518 (
            .O(N__55195),
            .I(N__55186));
    InMux I__10517 (
            .O(N__55194),
            .I(N__55183));
    LocalMux I__10516 (
            .O(N__55191),
            .I(N__55178));
    LocalMux I__10515 (
            .O(N__55186),
            .I(N__55178));
    LocalMux I__10514 (
            .O(N__55183),
            .I(N__55175));
    Span4Mux_v I__10513 (
            .O(N__55178),
            .I(N__55172));
    Span4Mux_h I__10512 (
            .O(N__55175),
            .I(N__55169));
    Span4Mux_h I__10511 (
            .O(N__55172),
            .I(N__55166));
    Odrv4 I__10510 (
            .O(N__55169),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_4_c_RNICGQM ));
    Odrv4 I__10509 (
            .O(N__55166),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_4_c_RNICGQM ));
    InMux I__10508 (
            .O(N__55161),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_4 ));
    InMux I__10507 (
            .O(N__55158),
            .I(N__55155));
    LocalMux I__10506 (
            .O(N__55155),
            .I(\pid_front.error_i_acummZ0Z_6 ));
    InMux I__10505 (
            .O(N__55152),
            .I(N__55145));
    InMux I__10504 (
            .O(N__55151),
            .I(N__55145));
    InMux I__10503 (
            .O(N__55150),
            .I(N__55142));
    LocalMux I__10502 (
            .O(N__55145),
            .I(N__55139));
    LocalMux I__10501 (
            .O(N__55142),
            .I(N__55136));
    Span4Mux_h I__10500 (
            .O(N__55139),
            .I(N__55133));
    Span4Mux_h I__10499 (
            .O(N__55136),
            .I(N__55128));
    Span4Mux_v I__10498 (
            .O(N__55133),
            .I(N__55128));
    Odrv4 I__10497 (
            .O(N__55128),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_5_c_RNIOULE ));
    InMux I__10496 (
            .O(N__55125),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_5 ));
    InMux I__10495 (
            .O(N__55122),
            .I(N__55119));
    LocalMux I__10494 (
            .O(N__55119),
            .I(\pid_front.error_i_acummZ0Z_7 ));
    InMux I__10493 (
            .O(N__55116),
            .I(N__55111));
    InMux I__10492 (
            .O(N__55115),
            .I(N__55106));
    InMux I__10491 (
            .O(N__55114),
            .I(N__55106));
    LocalMux I__10490 (
            .O(N__55111),
            .I(N__55103));
    LocalMux I__10489 (
            .O(N__55106),
            .I(N__55100));
    Span4Mux_h I__10488 (
            .O(N__55103),
            .I(N__55095));
    Span4Mux_h I__10487 (
            .O(N__55100),
            .I(N__55095));
    Odrv4 I__10486 (
            .O(N__55095),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_6_c_RNIR2NE ));
    InMux I__10485 (
            .O(N__55092),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_6 ));
    InMux I__10484 (
            .O(N__55089),
            .I(N__55086));
    LocalMux I__10483 (
            .O(N__55086),
            .I(\pid_front.error_i_acummZ0Z_8 ));
    InMux I__10482 (
            .O(N__55083),
            .I(N__55077));
    InMux I__10481 (
            .O(N__55082),
            .I(N__55077));
    LocalMux I__10480 (
            .O(N__55077),
            .I(N__55073));
    InMux I__10479 (
            .O(N__55076),
            .I(N__55070));
    Span4Mux_h I__10478 (
            .O(N__55073),
            .I(N__55067));
    LocalMux I__10477 (
            .O(N__55070),
            .I(N__55064));
    Span4Mux_v I__10476 (
            .O(N__55067),
            .I(N__55061));
    Odrv4 I__10475 (
            .O(N__55064),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_7_c_RNIU6OE ));
    Odrv4 I__10474 (
            .O(N__55061),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_7_c_RNIU6OE ));
    InMux I__10473 (
            .O(N__55056),
            .I(bfn_13_24_0_));
    InMux I__10472 (
            .O(N__55053),
            .I(N__55050));
    LocalMux I__10471 (
            .O(N__55050),
            .I(\pid_front.error_i_acummZ0Z_9 ));
    InMux I__10470 (
            .O(N__55047),
            .I(N__55044));
    LocalMux I__10469 (
            .O(N__55044),
            .I(N__55039));
    InMux I__10468 (
            .O(N__55043),
            .I(N__55034));
    InMux I__10467 (
            .O(N__55042),
            .I(N__55034));
    Span4Mux_h I__10466 (
            .O(N__55039),
            .I(N__55031));
    LocalMux I__10465 (
            .O(N__55034),
            .I(N__55028));
    Span4Mux_v I__10464 (
            .O(N__55031),
            .I(N__55025));
    Span12Mux_v I__10463 (
            .O(N__55028),
            .I(N__55022));
    Odrv4 I__10462 (
            .O(N__55025),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_8_c_RNI1BPE ));
    Odrv12 I__10461 (
            .O(N__55022),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_8_c_RNI1BPE ));
    InMux I__10460 (
            .O(N__55017),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_8 ));
    InMux I__10459 (
            .O(N__55014),
            .I(N__55011));
    LocalMux I__10458 (
            .O(N__55011),
            .I(\pid_front.error_i_acummZ0Z_10 ));
    InMux I__10457 (
            .O(N__55008),
            .I(N__55001));
    InMux I__10456 (
            .O(N__55007),
            .I(N__55001));
    InMux I__10455 (
            .O(N__55006),
            .I(N__54998));
    LocalMux I__10454 (
            .O(N__55001),
            .I(N__54995));
    LocalMux I__10453 (
            .O(N__54998),
            .I(N__54992));
    Span4Mux_v I__10452 (
            .O(N__54995),
            .I(N__54989));
    Span4Mux_h I__10451 (
            .O(N__54992),
            .I(N__54984));
    Span4Mux_h I__10450 (
            .O(N__54989),
            .I(N__54984));
    Odrv4 I__10449 (
            .O(N__54984),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_9_c_RNIIPQK ));
    InMux I__10448 (
            .O(N__54981),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_9 ));
    InMux I__10447 (
            .O(N__54978),
            .I(N__54975));
    LocalMux I__10446 (
            .O(N__54975),
            .I(\pid_front.error_i_acummZ0Z_11 ));
    InMux I__10445 (
            .O(N__54972),
            .I(N__54968));
    InMux I__10444 (
            .O(N__54971),
            .I(N__54965));
    LocalMux I__10443 (
            .O(N__54968),
            .I(N__54960));
    LocalMux I__10442 (
            .O(N__54965),
            .I(N__54957));
    InMux I__10441 (
            .O(N__54964),
            .I(N__54952));
    InMux I__10440 (
            .O(N__54963),
            .I(N__54952));
    Span4Mux_v I__10439 (
            .O(N__54960),
            .I(N__54945));
    Span4Mux_v I__10438 (
            .O(N__54957),
            .I(N__54945));
    LocalMux I__10437 (
            .O(N__54952),
            .I(N__54945));
    Odrv4 I__10436 (
            .O(N__54945),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_10_c_RNIJD4S ));
    InMux I__10435 (
            .O(N__54942),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_10 ));
    InMux I__10434 (
            .O(N__54939),
            .I(N__54936));
    LocalMux I__10433 (
            .O(N__54936),
            .I(\pid_front.error_i_acummZ0Z_12 ));
    InMux I__10432 (
            .O(N__54933),
            .I(N__54926));
    InMux I__10431 (
            .O(N__54932),
            .I(N__54926));
    InMux I__10430 (
            .O(N__54931),
            .I(N__54923));
    LocalMux I__10429 (
            .O(N__54926),
            .I(N__54920));
    LocalMux I__10428 (
            .O(N__54923),
            .I(N__54915));
    Span4Mux_h I__10427 (
            .O(N__54920),
            .I(N__54915));
    Odrv4 I__10426 (
            .O(N__54915),
            .I(\pid_front.error_i_reg_esr_RNIV4AUZ0Z_12 ));
    InMux I__10425 (
            .O(N__54912),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_11 ));
    InMux I__10424 (
            .O(N__54909),
            .I(N__54906));
    LocalMux I__10423 (
            .O(N__54906),
            .I(N__54903));
    Span4Mux_v I__10422 (
            .O(N__54903),
            .I(N__54900));
    Odrv4 I__10421 (
            .O(N__54900),
            .I(drone_H_disp_front_i_12));
    CascadeMux I__10420 (
            .O(N__54897),
            .I(N__54894));
    InMux I__10419 (
            .O(N__54894),
            .I(N__54890));
    InMux I__10418 (
            .O(N__54893),
            .I(N__54887));
    LocalMux I__10417 (
            .O(N__54890),
            .I(drone_H_disp_front_13));
    LocalMux I__10416 (
            .O(N__54887),
            .I(drone_H_disp_front_13));
    InMux I__10415 (
            .O(N__54882),
            .I(\pid_front.error_cry_8 ));
    InMux I__10414 (
            .O(N__54879),
            .I(N__54876));
    LocalMux I__10413 (
            .O(N__54876),
            .I(drone_H_disp_front_i_13));
    InMux I__10412 (
            .O(N__54873),
            .I(\pid_front.error_cry_9 ));
    InMux I__10411 (
            .O(N__54870),
            .I(N__54867));
    LocalMux I__10410 (
            .O(N__54867),
            .I(drone_H_disp_front_15));
    CascadeMux I__10409 (
            .O(N__54864),
            .I(N__54860));
    InMux I__10408 (
            .O(N__54863),
            .I(N__54855));
    InMux I__10407 (
            .O(N__54860),
            .I(N__54855));
    LocalMux I__10406 (
            .O(N__54855),
            .I(drone_H_disp_front_14));
    InMux I__10405 (
            .O(N__54852),
            .I(\pid_front.error_cry_10 ));
    CascadeMux I__10404 (
            .O(N__54849),
            .I(N__54846));
    InMux I__10403 (
            .O(N__54846),
            .I(N__54842));
    InMux I__10402 (
            .O(N__54845),
            .I(N__54839));
    LocalMux I__10401 (
            .O(N__54842),
            .I(N__54836));
    LocalMux I__10400 (
            .O(N__54839),
            .I(N__54833));
    Span4Mux_h I__10399 (
            .O(N__54836),
            .I(N__54830));
    Span4Mux_v I__10398 (
            .O(N__54833),
            .I(N__54827));
    Sp12to4 I__10397 (
            .O(N__54830),
            .I(N__54824));
    Odrv4 I__10396 (
            .O(N__54827),
            .I(\pid_front.un1_pid_prereg_0 ));
    Odrv12 I__10395 (
            .O(N__54824),
            .I(\pid_front.un1_pid_prereg_0 ));
    InMux I__10394 (
            .O(N__54819),
            .I(N__54816));
    LocalMux I__10393 (
            .O(N__54816),
            .I(\pid_front.error_i_acummZ0Z_1 ));
    CascadeMux I__10392 (
            .O(N__54813),
            .I(N__54810));
    InMux I__10391 (
            .O(N__54810),
            .I(N__54805));
    InMux I__10390 (
            .O(N__54809),
            .I(N__54802));
    InMux I__10389 (
            .O(N__54808),
            .I(N__54799));
    LocalMux I__10388 (
            .O(N__54805),
            .I(N__54796));
    LocalMux I__10387 (
            .O(N__54802),
            .I(N__54793));
    LocalMux I__10386 (
            .O(N__54799),
            .I(N__54790));
    Span4Mux_v I__10385 (
            .O(N__54796),
            .I(N__54787));
    Span4Mux_v I__10384 (
            .O(N__54793),
            .I(N__54784));
    Span4Mux_h I__10383 (
            .O(N__54790),
            .I(N__54779));
    Span4Mux_h I__10382 (
            .O(N__54787),
            .I(N__54779));
    Odrv4 I__10381 (
            .O(N__54784),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_0_c_RNI9AGE ));
    Odrv4 I__10380 (
            .O(N__54779),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_0_c_RNI9AGE ));
    InMux I__10379 (
            .O(N__54774),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_0 ));
    InMux I__10378 (
            .O(N__54771),
            .I(N__54768));
    LocalMux I__10377 (
            .O(N__54768),
            .I(\pid_front.error_i_acummZ0Z_2 ));
    CascadeMux I__10376 (
            .O(N__54765),
            .I(N__54762));
    InMux I__10375 (
            .O(N__54762),
            .I(N__54758));
    InMux I__10374 (
            .O(N__54761),
            .I(N__54754));
    LocalMux I__10373 (
            .O(N__54758),
            .I(N__54751));
    InMux I__10372 (
            .O(N__54757),
            .I(N__54748));
    LocalMux I__10371 (
            .O(N__54754),
            .I(N__54745));
    Span4Mux_v I__10370 (
            .O(N__54751),
            .I(N__54742));
    LocalMux I__10369 (
            .O(N__54748),
            .I(N__54739));
    Span4Mux_v I__10368 (
            .O(N__54745),
            .I(N__54736));
    Span4Mux_h I__10367 (
            .O(N__54742),
            .I(N__54733));
    Odrv4 I__10366 (
            .O(N__54739),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_1_c_RNICEHE ));
    Odrv4 I__10365 (
            .O(N__54736),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_1_c_RNICEHE ));
    Odrv4 I__10364 (
            .O(N__54733),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_1_c_RNICEHE ));
    InMux I__10363 (
            .O(N__54726),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_1 ));
    InMux I__10362 (
            .O(N__54723),
            .I(N__54720));
    LocalMux I__10361 (
            .O(N__54720),
            .I(\pid_front.error_i_acummZ0Z_3 ));
    InMux I__10360 (
            .O(N__54717),
            .I(N__54712));
    InMux I__10359 (
            .O(N__54716),
            .I(N__54707));
    InMux I__10358 (
            .O(N__54715),
            .I(N__54707));
    LocalMux I__10357 (
            .O(N__54712),
            .I(N__54704));
    LocalMux I__10356 (
            .O(N__54707),
            .I(N__54701));
    Span4Mux_h I__10355 (
            .O(N__54704),
            .I(N__54696));
    Span4Mux_v I__10354 (
            .O(N__54701),
            .I(N__54696));
    Odrv4 I__10353 (
            .O(N__54696),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_2_c_RNIFIIE ));
    InMux I__10352 (
            .O(N__54693),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_2 ));
    InMux I__10351 (
            .O(N__54690),
            .I(N__54687));
    LocalMux I__10350 (
            .O(N__54687),
            .I(\pid_front.error_i_acummZ0Z_4 ));
    InMux I__10349 (
            .O(N__54684),
            .I(N__54677));
    InMux I__10348 (
            .O(N__54683),
            .I(N__54677));
    InMux I__10347 (
            .O(N__54682),
            .I(N__54674));
    LocalMux I__10346 (
            .O(N__54677),
            .I(N__54671));
    LocalMux I__10345 (
            .O(N__54674),
            .I(N__54668));
    Span4Mux_v I__10344 (
            .O(N__54671),
            .I(N__54665));
    Span4Mux_h I__10343 (
            .O(N__54668),
            .I(N__54662));
    Span4Mux_h I__10342 (
            .O(N__54665),
            .I(N__54659));
    Odrv4 I__10341 (
            .O(N__54662),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_3_c_RNIIMJE ));
    Odrv4 I__10340 (
            .O(N__54659),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_3_c_RNIIMJE ));
    InMux I__10339 (
            .O(N__54654),
            .I(\pid_front.un1_error_i_acumm_prereg_cry_3 ));
    InMux I__10338 (
            .O(N__54651),
            .I(N__54648));
    LocalMux I__10337 (
            .O(N__54648),
            .I(drone_H_disp_front_i_5));
    CascadeMux I__10336 (
            .O(N__54645),
            .I(N__54642));
    InMux I__10335 (
            .O(N__54642),
            .I(N__54639));
    LocalMux I__10334 (
            .O(N__54639),
            .I(front_command_1));
    InMux I__10333 (
            .O(N__54636),
            .I(\pid_front.error_cry_0_0 ));
    InMux I__10332 (
            .O(N__54633),
            .I(N__54630));
    LocalMux I__10331 (
            .O(N__54630),
            .I(drone_H_disp_front_i_6));
    CascadeMux I__10330 (
            .O(N__54627),
            .I(N__54624));
    InMux I__10329 (
            .O(N__54624),
            .I(N__54621));
    LocalMux I__10328 (
            .O(N__54621),
            .I(front_command_2));
    InMux I__10327 (
            .O(N__54618),
            .I(\pid_front.error_cry_1_0 ));
    InMux I__10326 (
            .O(N__54615),
            .I(N__54612));
    LocalMux I__10325 (
            .O(N__54612),
            .I(drone_H_disp_front_i_7));
    CascadeMux I__10324 (
            .O(N__54609),
            .I(N__54606));
    InMux I__10323 (
            .O(N__54606),
            .I(N__54603));
    LocalMux I__10322 (
            .O(N__54603),
            .I(front_command_3));
    InMux I__10321 (
            .O(N__54600),
            .I(\pid_front.error_cry_2_0 ));
    InMux I__10320 (
            .O(N__54597),
            .I(N__54594));
    LocalMux I__10319 (
            .O(N__54594),
            .I(drone_H_disp_front_i_8));
    CascadeMux I__10318 (
            .O(N__54591),
            .I(N__54588));
    InMux I__10317 (
            .O(N__54588),
            .I(N__54585));
    LocalMux I__10316 (
            .O(N__54585),
            .I(N__54582));
    Odrv4 I__10315 (
            .O(N__54582),
            .I(front_command_4));
    InMux I__10314 (
            .O(N__54579),
            .I(bfn_13_22_0_));
    InMux I__10313 (
            .O(N__54576),
            .I(N__54573));
    LocalMux I__10312 (
            .O(N__54573),
            .I(drone_H_disp_front_i_9));
    CascadeMux I__10311 (
            .O(N__54570),
            .I(N__54567));
    InMux I__10310 (
            .O(N__54567),
            .I(N__54564));
    LocalMux I__10309 (
            .O(N__54564),
            .I(N__54561));
    Span4Mux_h I__10308 (
            .O(N__54561),
            .I(N__54558));
    Odrv4 I__10307 (
            .O(N__54558),
            .I(front_command_5));
    InMux I__10306 (
            .O(N__54555),
            .I(\pid_front.error_cry_4 ));
    InMux I__10305 (
            .O(N__54552),
            .I(N__54549));
    LocalMux I__10304 (
            .O(N__54549),
            .I(N__54546));
    Odrv4 I__10303 (
            .O(N__54546),
            .I(front_command_6));
    CascadeMux I__10302 (
            .O(N__54543),
            .I(N__54540));
    InMux I__10301 (
            .O(N__54540),
            .I(N__54537));
    LocalMux I__10300 (
            .O(N__54537),
            .I(drone_H_disp_front_i_10));
    InMux I__10299 (
            .O(N__54534),
            .I(\pid_front.error_cry_5 ));
    InMux I__10298 (
            .O(N__54531),
            .I(N__54528));
    LocalMux I__10297 (
            .O(N__54528),
            .I(N__54525));
    Span4Mux_v I__10296 (
            .O(N__54525),
            .I(N__54522));
    Odrv4 I__10295 (
            .O(N__54522),
            .I(\pid_front.error_axbZ0Z_7 ));
    InMux I__10294 (
            .O(N__54519),
            .I(\pid_front.error_cry_6 ));
    InMux I__10293 (
            .O(N__54516),
            .I(N__54513));
    LocalMux I__10292 (
            .O(N__54513),
            .I(N__54510));
    Odrv4 I__10291 (
            .O(N__54510),
            .I(\pid_front.error_axb_8_l_ofx_0 ));
    CascadeMux I__10290 (
            .O(N__54507),
            .I(N__54502));
    InMux I__10289 (
            .O(N__54506),
            .I(N__54499));
    InMux I__10288 (
            .O(N__54505),
            .I(N__54496));
    InMux I__10287 (
            .O(N__54502),
            .I(N__54493));
    LocalMux I__10286 (
            .O(N__54499),
            .I(N__54490));
    LocalMux I__10285 (
            .O(N__54496),
            .I(drone_H_disp_front_12));
    LocalMux I__10284 (
            .O(N__54493),
            .I(drone_H_disp_front_12));
    Odrv4 I__10283 (
            .O(N__54490),
            .I(drone_H_disp_front_12));
    InMux I__10282 (
            .O(N__54483),
            .I(\pid_front.error_cry_7 ));
    InMux I__10281 (
            .O(N__54480),
            .I(N__54477));
    LocalMux I__10280 (
            .O(N__54477),
            .I(N__54473));
    InMux I__10279 (
            .O(N__54476),
            .I(N__54470));
    Span4Mux_h I__10278 (
            .O(N__54473),
            .I(N__54467));
    LocalMux I__10277 (
            .O(N__54470),
            .I(front_command_7));
    Odrv4 I__10276 (
            .O(N__54467),
            .I(front_command_7));
    InMux I__10275 (
            .O(N__54462),
            .I(N__54458));
    InMux I__10274 (
            .O(N__54461),
            .I(N__54455));
    LocalMux I__10273 (
            .O(N__54458),
            .I(N__54452));
    LocalMux I__10272 (
            .O(N__54455),
            .I(drone_H_disp_front_11));
    Odrv4 I__10271 (
            .O(N__54452),
            .I(drone_H_disp_front_11));
    CascadeMux I__10270 (
            .O(N__54447),
            .I(N__54444));
    InMux I__10269 (
            .O(N__54444),
            .I(N__54441));
    LocalMux I__10268 (
            .O(N__54441),
            .I(\pid_front.error_axb_0 ));
    InMux I__10267 (
            .O(N__54438),
            .I(N__54435));
    LocalMux I__10266 (
            .O(N__54435),
            .I(N__54432));
    Odrv4 I__10265 (
            .O(N__54432),
            .I(\pid_front.error_axbZ0Z_1 ));
    InMux I__10264 (
            .O(N__54429),
            .I(\pid_front.error_cry_0 ));
    InMux I__10263 (
            .O(N__54426),
            .I(N__54423));
    LocalMux I__10262 (
            .O(N__54423),
            .I(N__54420));
    Odrv4 I__10261 (
            .O(N__54420),
            .I(\pid_front.error_axbZ0Z_2 ));
    InMux I__10260 (
            .O(N__54417),
            .I(\pid_front.error_cry_1 ));
    InMux I__10259 (
            .O(N__54414),
            .I(N__54411));
    LocalMux I__10258 (
            .O(N__54411),
            .I(N__54408));
    Odrv4 I__10257 (
            .O(N__54408),
            .I(\pid_front.error_axbZ0Z_3 ));
    InMux I__10256 (
            .O(N__54405),
            .I(\pid_front.error_cry_2 ));
    InMux I__10255 (
            .O(N__54402),
            .I(N__54399));
    LocalMux I__10254 (
            .O(N__54399),
            .I(drone_H_disp_front_i_4));
    CascadeMux I__10253 (
            .O(N__54396),
            .I(N__54393));
    InMux I__10252 (
            .O(N__54393),
            .I(N__54390));
    LocalMux I__10251 (
            .O(N__54390),
            .I(front_command_0));
    InMux I__10250 (
            .O(N__54387),
            .I(\pid_front.error_cry_3 ));
    InMux I__10249 (
            .O(N__54384),
            .I(N__54381));
    LocalMux I__10248 (
            .O(N__54381),
            .I(drone_H_disp_side_1));
    InMux I__10247 (
            .O(N__54378),
            .I(N__54374));
    InMux I__10246 (
            .O(N__54377),
            .I(N__54371));
    LocalMux I__10245 (
            .O(N__54374),
            .I(N__54368));
    LocalMux I__10244 (
            .O(N__54371),
            .I(N__54365));
    Span12Mux_v I__10243 (
            .O(N__54368),
            .I(N__54362));
    Span12Mux_v I__10242 (
            .O(N__54365),
            .I(N__54359));
    Span12Mux_h I__10241 (
            .O(N__54362),
            .I(N__54356));
    Span12Mux_h I__10240 (
            .O(N__54359),
            .I(N__54353));
    Odrv12 I__10239 (
            .O(N__54356),
            .I(xy_kd_2));
    Odrv12 I__10238 (
            .O(N__54353),
            .I(xy_kd_2));
    InMux I__10237 (
            .O(N__54348),
            .I(N__54344));
    InMux I__10236 (
            .O(N__54347),
            .I(N__54341));
    LocalMux I__10235 (
            .O(N__54344),
            .I(N__54338));
    LocalMux I__10234 (
            .O(N__54341),
            .I(N__54335));
    Sp12to4 I__10233 (
            .O(N__54338),
            .I(N__54330));
    Span12Mux_v I__10232 (
            .O(N__54335),
            .I(N__54330));
    Span12Mux_h I__10231 (
            .O(N__54330),
            .I(N__54327));
    Odrv12 I__10230 (
            .O(N__54327),
            .I(xy_kd_6));
    InMux I__10229 (
            .O(N__54324),
            .I(N__54321));
    LocalMux I__10228 (
            .O(N__54321),
            .I(N__54318));
    Odrv12 I__10227 (
            .O(N__54318),
            .I(\dron_frame_decoder_1.drone_altitude_11 ));
    InMux I__10226 (
            .O(N__54315),
            .I(N__54312));
    LocalMux I__10225 (
            .O(N__54312),
            .I(N__54309));
    Span12Mux_s10_h I__10224 (
            .O(N__54309),
            .I(N__54306));
    Odrv12 I__10223 (
            .O(N__54306),
            .I(drone_altitude_i_11));
    InMux I__10222 (
            .O(N__54303),
            .I(N__54298));
    InMux I__10221 (
            .O(N__54302),
            .I(N__54295));
    InMux I__10220 (
            .O(N__54301),
            .I(N__54292));
    LocalMux I__10219 (
            .O(N__54298),
            .I(N__54286));
    LocalMux I__10218 (
            .O(N__54295),
            .I(N__54286));
    LocalMux I__10217 (
            .O(N__54292),
            .I(N__54283));
    InMux I__10216 (
            .O(N__54291),
            .I(N__54280));
    Span4Mux_v I__10215 (
            .O(N__54286),
            .I(N__54277));
    Odrv4 I__10214 (
            .O(N__54283),
            .I(\pid_front.error_d_reg_prevZ0Z_14 ));
    LocalMux I__10213 (
            .O(N__54280),
            .I(\pid_front.error_d_reg_prevZ0Z_14 ));
    Odrv4 I__10212 (
            .O(N__54277),
            .I(\pid_front.error_d_reg_prevZ0Z_14 ));
    InMux I__10211 (
            .O(N__54270),
            .I(N__54265));
    CascadeMux I__10210 (
            .O(N__54269),
            .I(N__54262));
    InMux I__10209 (
            .O(N__54268),
            .I(N__54259));
    LocalMux I__10208 (
            .O(N__54265),
            .I(N__54256));
    InMux I__10207 (
            .O(N__54262),
            .I(N__54252));
    LocalMux I__10206 (
            .O(N__54259),
            .I(N__54249));
    Span4Mux_v I__10205 (
            .O(N__54256),
            .I(N__54246));
    InMux I__10204 (
            .O(N__54255),
            .I(N__54243));
    LocalMux I__10203 (
            .O(N__54252),
            .I(N__54240));
    Span4Mux_h I__10202 (
            .O(N__54249),
            .I(N__54237));
    Span4Mux_h I__10201 (
            .O(N__54246),
            .I(N__54232));
    LocalMux I__10200 (
            .O(N__54243),
            .I(N__54232));
    Span4Mux_h I__10199 (
            .O(N__54240),
            .I(N__54227));
    Span4Mux_h I__10198 (
            .O(N__54237),
            .I(N__54227));
    Span4Mux_h I__10197 (
            .O(N__54232),
            .I(N__54224));
    Sp12to4 I__10196 (
            .O(N__54227),
            .I(N__54219));
    Sp12to4 I__10195 (
            .O(N__54224),
            .I(N__54219));
    Span12Mux_v I__10194 (
            .O(N__54219),
            .I(N__54216));
    Odrv12 I__10193 (
            .O(N__54216),
            .I(\pid_front.error_p_regZ0Z_14 ));
    InMux I__10192 (
            .O(N__54213),
            .I(N__54210));
    LocalMux I__10191 (
            .O(N__54210),
            .I(N__54207));
    Span12Mux_h I__10190 (
            .O(N__54207),
            .I(N__54204));
    Odrv12 I__10189 (
            .O(N__54204),
            .I(\pid_front.error_p_reg_esr_RNIH0C61_0Z0Z_14 ));
    InMux I__10188 (
            .O(N__54201),
            .I(N__54198));
    LocalMux I__10187 (
            .O(N__54198),
            .I(drone_H_disp_side_3));
    CEMux I__10186 (
            .O(N__54195),
            .I(N__54191));
    CEMux I__10185 (
            .O(N__54194),
            .I(N__54188));
    LocalMux I__10184 (
            .O(N__54191),
            .I(N__54185));
    LocalMux I__10183 (
            .O(N__54188),
            .I(N__54182));
    Span4Mux_h I__10182 (
            .O(N__54185),
            .I(N__54179));
    Sp12to4 I__10181 (
            .O(N__54182),
            .I(N__54176));
    Span4Mux_h I__10180 (
            .O(N__54179),
            .I(N__54173));
    Span12Mux_h I__10179 (
            .O(N__54176),
            .I(N__54170));
    Odrv4 I__10178 (
            .O(N__54173),
            .I(\dron_frame_decoder_1.N_724_0 ));
    Odrv12 I__10177 (
            .O(N__54170),
            .I(\dron_frame_decoder_1.N_724_0 ));
    InMux I__10176 (
            .O(N__54165),
            .I(N__54162));
    LocalMux I__10175 (
            .O(N__54162),
            .I(N__54159));
    Span12Mux_s9_h I__10174 (
            .O(N__54159),
            .I(N__54156));
    Odrv12 I__10173 (
            .O(N__54156),
            .I(\pid_alt.error_axbZ0Z_2 ));
    InMux I__10172 (
            .O(N__54153),
            .I(N__54150));
    LocalMux I__10171 (
            .O(N__54150),
            .I(drone_altitude_2));
    InMux I__10170 (
            .O(N__54147),
            .I(N__54144));
    LocalMux I__10169 (
            .O(N__54144),
            .I(N__54141));
    Span12Mux_s7_h I__10168 (
            .O(N__54141),
            .I(N__54138));
    Odrv12 I__10167 (
            .O(N__54138),
            .I(\pid_alt.error_axbZ0Z_3 ));
    InMux I__10166 (
            .O(N__54135),
            .I(N__54132));
    LocalMux I__10165 (
            .O(N__54132),
            .I(drone_altitude_3));
    CEMux I__10164 (
            .O(N__54129),
            .I(N__54126));
    LocalMux I__10163 (
            .O(N__54126),
            .I(N__54122));
    CEMux I__10162 (
            .O(N__54125),
            .I(N__54119));
    Span4Mux_v I__10161 (
            .O(N__54122),
            .I(N__54116));
    LocalMux I__10160 (
            .O(N__54119),
            .I(N__54113));
    Span4Mux_h I__10159 (
            .O(N__54116),
            .I(N__54110));
    Span4Mux_h I__10158 (
            .O(N__54113),
            .I(N__54107));
    Span4Mux_h I__10157 (
            .O(N__54110),
            .I(N__54102));
    Span4Mux_v I__10156 (
            .O(N__54107),
            .I(N__54102));
    Odrv4 I__10155 (
            .O(N__54102),
            .I(\dron_frame_decoder_1.N_740_0 ));
    CascadeMux I__10154 (
            .O(N__54099),
            .I(\pid_side.error_i_reg_9_rn_0_26_cascade_ ));
    CascadeMux I__10153 (
            .O(N__54096),
            .I(\pid_side.m6_2_03_cascade_ ));
    InMux I__10152 (
            .O(N__54093),
            .I(N__54087));
    InMux I__10151 (
            .O(N__54092),
            .I(N__54087));
    LocalMux I__10150 (
            .O(N__54087),
            .I(\pid_side.N_39_1 ));
    CascadeMux I__10149 (
            .O(N__54084),
            .I(\pid_side.error_i_reg_9_rn_0_18_cascade_ ));
    InMux I__10148 (
            .O(N__54081),
            .I(N__54078));
    LocalMux I__10147 (
            .O(N__54078),
            .I(drone_H_disp_side_2));
    InMux I__10146 (
            .O(N__54075),
            .I(N__54072));
    LocalMux I__10145 (
            .O(N__54072),
            .I(\pid_side.m36_1_ns_1 ));
    CascadeMux I__10144 (
            .O(N__54069),
            .I(\pid_side.N_37_1_cascade_ ));
    CascadeMux I__10143 (
            .O(N__54066),
            .I(\pid_side.N_39_1_cascade_ ));
    CascadeMux I__10142 (
            .O(N__54063),
            .I(\pid_side.N_126_0_cascade_ ));
    CascadeMux I__10141 (
            .O(N__54060),
            .I(\pid_side.m2_0_03_3_i_0_cascade_ ));
    InMux I__10140 (
            .O(N__54057),
            .I(N__54054));
    LocalMux I__10139 (
            .O(N__54054),
            .I(\pid_side.N_41_0 ));
    CascadeMux I__10138 (
            .O(N__54051),
            .I(\pid_side.N_41_0_cascade_ ));
    InMux I__10137 (
            .O(N__54048),
            .I(N__54045));
    LocalMux I__10136 (
            .O(N__54045),
            .I(\pid_side.error_p_reg_esr_RNISPTC1Z0Z_8 ));
    InMux I__10135 (
            .O(N__54042),
            .I(N__54036));
    InMux I__10134 (
            .O(N__54041),
            .I(N__54036));
    LocalMux I__10133 (
            .O(N__54036),
            .I(\pid_side.error_p_reg_esr_RNI1VTC1_0Z0Z_9 ));
    InMux I__10132 (
            .O(N__54033),
            .I(N__54030));
    LocalMux I__10131 (
            .O(N__54030),
            .I(\pid_side.N_2374_i ));
    InMux I__10130 (
            .O(N__54027),
            .I(N__54023));
    CascadeMux I__10129 (
            .O(N__54026),
            .I(N__54020));
    LocalMux I__10128 (
            .O(N__54023),
            .I(N__54016));
    InMux I__10127 (
            .O(N__54020),
            .I(N__54011));
    InMux I__10126 (
            .O(N__54019),
            .I(N__54011));
    Span4Mux_v I__10125 (
            .O(N__54016),
            .I(N__54008));
    LocalMux I__10124 (
            .O(N__54011),
            .I(\pid_side.error_d_reg_prevZ0Z_7 ));
    Odrv4 I__10123 (
            .O(N__54008),
            .I(\pid_side.error_d_reg_prevZ0Z_7 ));
    CascadeMux I__10122 (
            .O(N__54003),
            .I(\pid_side.N_2374_i_cascade_ ));
    InMux I__10121 (
            .O(N__54000),
            .I(N__53993));
    InMux I__10120 (
            .O(N__53999),
            .I(N__53993));
    InMux I__10119 (
            .O(N__53998),
            .I(N__53990));
    LocalMux I__10118 (
            .O(N__53993),
            .I(\pid_side.error_d_reg_prevZ0Z_8 ));
    LocalMux I__10117 (
            .O(N__53990),
            .I(\pid_side.error_d_reg_prevZ0Z_8 ));
    CascadeMux I__10116 (
            .O(N__53985),
            .I(\pid_side.error_i_reg_esr_RNO_0Z0Z_22_cascade_ ));
    InMux I__10115 (
            .O(N__53982),
            .I(N__53979));
    LocalMux I__10114 (
            .O(N__53979),
            .I(N__53975));
    CascadeMux I__10113 (
            .O(N__53978),
            .I(N__53972));
    Span4Mux_v I__10112 (
            .O(N__53975),
            .I(N__53969));
    InMux I__10111 (
            .O(N__53972),
            .I(N__53966));
    Span4Mux_v I__10110 (
            .O(N__53969),
            .I(N__53958));
    LocalMux I__10109 (
            .O(N__53966),
            .I(N__53958));
    CascadeMux I__10108 (
            .O(N__53965),
            .I(N__53955));
    InMux I__10107 (
            .O(N__53964),
            .I(N__53950));
    InMux I__10106 (
            .O(N__53963),
            .I(N__53950));
    Span4Mux_h I__10105 (
            .O(N__53958),
            .I(N__53947));
    InMux I__10104 (
            .O(N__53955),
            .I(N__53944));
    LocalMux I__10103 (
            .O(N__53950),
            .I(N__53939));
    Span4Mux_h I__10102 (
            .O(N__53947),
            .I(N__53939));
    LocalMux I__10101 (
            .O(N__53944),
            .I(\ppm_encoder_1.N_257_i_i ));
    Odrv4 I__10100 (
            .O(N__53939),
            .I(\ppm_encoder_1.N_257_i_i ));
    InMux I__10099 (
            .O(N__53934),
            .I(N__53931));
    LocalMux I__10098 (
            .O(N__53931),
            .I(N__53927));
    InMux I__10097 (
            .O(N__53930),
            .I(N__53924));
    Span4Mux_v I__10096 (
            .O(N__53927),
            .I(N__53921));
    LocalMux I__10095 (
            .O(N__53924),
            .I(N__53918));
    Sp12to4 I__10094 (
            .O(N__53921),
            .I(N__53913));
    Span12Mux_v I__10093 (
            .O(N__53918),
            .I(N__53913));
    Odrv12 I__10092 (
            .O(N__53913),
            .I(frame_decoder_OFF4data_7));
    InMux I__10091 (
            .O(N__53910),
            .I(N__53907));
    LocalMux I__10090 (
            .O(N__53907),
            .I(N__53904));
    Span4Mux_v I__10089 (
            .O(N__53904),
            .I(N__53901));
    Span4Mux_h I__10088 (
            .O(N__53901),
            .I(N__53898));
    Span4Mux_h I__10087 (
            .O(N__53898),
            .I(N__53894));
    InMux I__10086 (
            .O(N__53897),
            .I(N__53891));
    Odrv4 I__10085 (
            .O(N__53894),
            .I(frame_decoder_CH4data_7));
    LocalMux I__10084 (
            .O(N__53891),
            .I(frame_decoder_CH4data_7));
    InMux I__10083 (
            .O(N__53886),
            .I(N__53883));
    LocalMux I__10082 (
            .O(N__53883),
            .I(N__53880));
    Span4Mux_v I__10081 (
            .O(N__53880),
            .I(N__53877));
    Odrv4 I__10080 (
            .O(N__53877),
            .I(\scaler_4.N_2725_i_l_ofxZ0 ));
    CascadeMux I__10079 (
            .O(N__53874),
            .I(\pid_side.error_p_reg_esr_RNISPTC1Z0Z_8_cascade_ ));
    InMux I__10078 (
            .O(N__53871),
            .I(N__53867));
    InMux I__10077 (
            .O(N__53870),
            .I(N__53864));
    LocalMux I__10076 (
            .O(N__53867),
            .I(N__53861));
    LocalMux I__10075 (
            .O(N__53864),
            .I(side_order_3));
    Odrv4 I__10074 (
            .O(N__53861),
            .I(side_order_3));
    InMux I__10073 (
            .O(N__53856),
            .I(N__53852));
    InMux I__10072 (
            .O(N__53855),
            .I(N__53849));
    LocalMux I__10071 (
            .O(N__53852),
            .I(N__53846));
    LocalMux I__10070 (
            .O(N__53849),
            .I(N__53843));
    Span4Mux_v I__10069 (
            .O(N__53846),
            .I(N__53840));
    Span4Mux_h I__10068 (
            .O(N__53843),
            .I(N__53837));
    Odrv4 I__10067 (
            .O(N__53840),
            .I(side_order_11));
    Odrv4 I__10066 (
            .O(N__53837),
            .I(side_order_11));
    InMux I__10065 (
            .O(N__53832),
            .I(N__53829));
    LocalMux I__10064 (
            .O(N__53829),
            .I(N__53825));
    InMux I__10063 (
            .O(N__53828),
            .I(N__53822));
    Sp12to4 I__10062 (
            .O(N__53825),
            .I(N__53819));
    LocalMux I__10061 (
            .O(N__53822),
            .I(N__53816));
    Odrv12 I__10060 (
            .O(N__53819),
            .I(side_order_1));
    Odrv4 I__10059 (
            .O(N__53816),
            .I(side_order_1));
    InMux I__10058 (
            .O(N__53811),
            .I(N__53807));
    InMux I__10057 (
            .O(N__53810),
            .I(N__53804));
    LocalMux I__10056 (
            .O(N__53807),
            .I(N__53801));
    LocalMux I__10055 (
            .O(N__53804),
            .I(N__53798));
    Odrv12 I__10054 (
            .O(N__53801),
            .I(side_order_0));
    Odrv4 I__10053 (
            .O(N__53798),
            .I(side_order_0));
    InMux I__10052 (
            .O(N__53793),
            .I(N__53790));
    LocalMux I__10051 (
            .O(N__53790),
            .I(N__53787));
    Span4Mux_h I__10050 (
            .O(N__53787),
            .I(N__53783));
    InMux I__10049 (
            .O(N__53786),
            .I(N__53780));
    Span4Mux_v I__10048 (
            .O(N__53783),
            .I(N__53775));
    LocalMux I__10047 (
            .O(N__53780),
            .I(N__53775));
    Span4Mux_h I__10046 (
            .O(N__53775),
            .I(N__53772));
    Odrv4 I__10045 (
            .O(N__53772),
            .I(side_order_10));
    CascadeMux I__10044 (
            .O(N__53769),
            .I(N__53765));
    InMux I__10043 (
            .O(N__53768),
            .I(N__53762));
    InMux I__10042 (
            .O(N__53765),
            .I(N__53759));
    LocalMux I__10041 (
            .O(N__53762),
            .I(N__53756));
    LocalMux I__10040 (
            .O(N__53759),
            .I(N__53753));
    Odrv4 I__10039 (
            .O(N__53756),
            .I(side_order_4));
    Odrv4 I__10038 (
            .O(N__53753),
            .I(side_order_4));
    InMux I__10037 (
            .O(N__53748),
            .I(N__53745));
    LocalMux I__10036 (
            .O(N__53745),
            .I(N__53741));
    InMux I__10035 (
            .O(N__53744),
            .I(N__53738));
    Span4Mux_v I__10034 (
            .O(N__53741),
            .I(N__53733));
    LocalMux I__10033 (
            .O(N__53738),
            .I(N__53733));
    Odrv4 I__10032 (
            .O(N__53733),
            .I(side_order_8));
    InMux I__10031 (
            .O(N__53730),
            .I(N__53727));
    LocalMux I__10030 (
            .O(N__53727),
            .I(N__53723));
    InMux I__10029 (
            .O(N__53726),
            .I(N__53720));
    Span4Mux_v I__10028 (
            .O(N__53723),
            .I(N__53715));
    LocalMux I__10027 (
            .O(N__53720),
            .I(N__53715));
    Odrv4 I__10026 (
            .O(N__53715),
            .I(side_order_9));
    InMux I__10025 (
            .O(N__53712),
            .I(N__53709));
    LocalMux I__10024 (
            .O(N__53709),
            .I(N__53705));
    InMux I__10023 (
            .O(N__53708),
            .I(N__53702));
    Span4Mux_v I__10022 (
            .O(N__53705),
            .I(N__53699));
    LocalMux I__10021 (
            .O(N__53702),
            .I(N__53696));
    Odrv4 I__10020 (
            .O(N__53699),
            .I(scaler_4_data_13));
    Odrv4 I__10019 (
            .O(N__53696),
            .I(scaler_4_data_13));
    InMux I__10018 (
            .O(N__53691),
            .I(N__53688));
    LocalMux I__10017 (
            .O(N__53688),
            .I(N__53685));
    Span4Mux_h I__10016 (
            .O(N__53685),
            .I(N__53682));
    Odrv4 I__10015 (
            .O(N__53682),
            .I(\ppm_encoder_1.un1_rudder_cry_12_THRU_CO ));
    CascadeMux I__10014 (
            .O(N__53679),
            .I(N__53675));
    InMux I__10013 (
            .O(N__53678),
            .I(N__53672));
    InMux I__10012 (
            .O(N__53675),
            .I(N__53668));
    LocalMux I__10011 (
            .O(N__53672),
            .I(N__53665));
    InMux I__10010 (
            .O(N__53671),
            .I(N__53662));
    LocalMux I__10009 (
            .O(N__53668),
            .I(N__53657));
    Span4Mux_h I__10008 (
            .O(N__53665),
            .I(N__53657));
    LocalMux I__10007 (
            .O(N__53662),
            .I(\ppm_encoder_1.aileronZ0Z_7 ));
    Odrv4 I__10006 (
            .O(N__53657),
            .I(\ppm_encoder_1.aileronZ0Z_7 ));
    CascadeMux I__10005 (
            .O(N__53652),
            .I(N__53648));
    CascadeMux I__10004 (
            .O(N__53651),
            .I(N__53644));
    InMux I__10003 (
            .O(N__53648),
            .I(N__53641));
    InMux I__10002 (
            .O(N__53647),
            .I(N__53638));
    InMux I__10001 (
            .O(N__53644),
            .I(N__53635));
    LocalMux I__10000 (
            .O(N__53641),
            .I(N__53632));
    LocalMux I__9999 (
            .O(N__53638),
            .I(N__53625));
    LocalMux I__9998 (
            .O(N__53635),
            .I(N__53625));
    Span4Mux_v I__9997 (
            .O(N__53632),
            .I(N__53625));
    Odrv4 I__9996 (
            .O(N__53625),
            .I(\ppm_encoder_1.throttleZ0Z_7 ));
    InMux I__9995 (
            .O(N__53622),
            .I(N__53619));
    LocalMux I__9994 (
            .O(N__53619),
            .I(N__53615));
    InMux I__9993 (
            .O(N__53618),
            .I(N__53612));
    Span4Mux_v I__9992 (
            .O(N__53615),
            .I(N__53608));
    LocalMux I__9991 (
            .O(N__53612),
            .I(N__53605));
    InMux I__9990 (
            .O(N__53611),
            .I(N__53602));
    Span4Mux_v I__9989 (
            .O(N__53608),
            .I(N__53597));
    Span4Mux_s1_v I__9988 (
            .O(N__53605),
            .I(N__53597));
    LocalMux I__9987 (
            .O(N__53602),
            .I(\ppm_encoder_1.rudderZ0Z_11 ));
    Odrv4 I__9986 (
            .O(N__53597),
            .I(\ppm_encoder_1.rudderZ0Z_11 ));
    InMux I__9985 (
            .O(N__53592),
            .I(N__53589));
    LocalMux I__9984 (
            .O(N__53589),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_11 ));
    InMux I__9983 (
            .O(N__53586),
            .I(N__53583));
    LocalMux I__9982 (
            .O(N__53583),
            .I(N__53580));
    Sp12to4 I__9981 (
            .O(N__53580),
            .I(N__53575));
    InMux I__9980 (
            .O(N__53579),
            .I(N__53572));
    InMux I__9979 (
            .O(N__53578),
            .I(N__53569));
    Span12Mux_s1_v I__9978 (
            .O(N__53575),
            .I(N__53564));
    LocalMux I__9977 (
            .O(N__53572),
            .I(N__53564));
    LocalMux I__9976 (
            .O(N__53569),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_3 ));
    Odrv12 I__9975 (
            .O(N__53564),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_3 ));
    CascadeMux I__9974 (
            .O(N__53559),
            .I(N__53556));
    InMux I__9973 (
            .O(N__53556),
            .I(N__53552));
    InMux I__9972 (
            .O(N__53555),
            .I(N__53549));
    LocalMux I__9971 (
            .O(N__53552),
            .I(\ppm_encoder_1.rudderZ0Z_13 ));
    LocalMux I__9970 (
            .O(N__53549),
            .I(\ppm_encoder_1.rudderZ0Z_13 ));
    InMux I__9969 (
            .O(N__53544),
            .I(N__53538));
    InMux I__9968 (
            .O(N__53543),
            .I(N__53538));
    LocalMux I__9967 (
            .O(N__53538),
            .I(\ppm_encoder_1.rudder_RNIN2KQZ0Z_13 ));
    InMux I__9966 (
            .O(N__53535),
            .I(N__53531));
    CascadeMux I__9965 (
            .O(N__53534),
            .I(N__53528));
    LocalMux I__9964 (
            .O(N__53531),
            .I(N__53525));
    InMux I__9963 (
            .O(N__53528),
            .I(N__53522));
    Span4Mux_h I__9962 (
            .O(N__53525),
            .I(N__53519));
    LocalMux I__9961 (
            .O(N__53522),
            .I(N__53516));
    Odrv4 I__9960 (
            .O(N__53519),
            .I(side_order_5));
    Odrv12 I__9959 (
            .O(N__53516),
            .I(side_order_5));
    InMux I__9958 (
            .O(N__53511),
            .I(N__53507));
    InMux I__9957 (
            .O(N__53510),
            .I(N__53504));
    LocalMux I__9956 (
            .O(N__53507),
            .I(N__53501));
    LocalMux I__9955 (
            .O(N__53504),
            .I(side_order_7));
    Odrv4 I__9954 (
            .O(N__53501),
            .I(side_order_7));
    CascadeMux I__9953 (
            .O(N__53496),
            .I(\ppm_encoder_1.un2_throttle_iv_0_0_1_7_cascade_ ));
    InMux I__9952 (
            .O(N__53493),
            .I(N__53490));
    LocalMux I__9951 (
            .O(N__53490),
            .I(\ppm_encoder_1.un2_throttle_iv_0_0_0_7 ));
    CascadeMux I__9950 (
            .O(N__53487),
            .I(N__53484));
    InMux I__9949 (
            .O(N__53484),
            .I(N__53481));
    LocalMux I__9948 (
            .O(N__53481),
            .I(N__53478));
    Span4Mux_v I__9947 (
            .O(N__53478),
            .I(N__53475));
    Odrv4 I__9946 (
            .O(N__53475),
            .I(\ppm_encoder_1.N_263_i_i ));
    CascadeMux I__9945 (
            .O(N__53472),
            .I(\ppm_encoder_1.N_263_i_i_cascade_ ));
    InMux I__9944 (
            .O(N__53469),
            .I(N__53466));
    LocalMux I__9943 (
            .O(N__53466),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_7 ));
    InMux I__9942 (
            .O(N__53463),
            .I(N__53460));
    LocalMux I__9941 (
            .O(N__53460),
            .I(N__53457));
    Span4Mux_h I__9940 (
            .O(N__53457),
            .I(N__53454));
    Odrv4 I__9939 (
            .O(N__53454),
            .I(\ppm_encoder_1.init_pulses_RNI2VJU5Z0Z_7 ));
    CascadeMux I__9938 (
            .O(N__53451),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_13_cascade_ ));
    CascadeMux I__9937 (
            .O(N__53448),
            .I(N__53445));
    InMux I__9936 (
            .O(N__53445),
            .I(N__53441));
    InMux I__9935 (
            .O(N__53444),
            .I(N__53438));
    LocalMux I__9934 (
            .O(N__53441),
            .I(N__53434));
    LocalMux I__9933 (
            .O(N__53438),
            .I(N__53431));
    InMux I__9932 (
            .O(N__53437),
            .I(N__53428));
    Span4Mux_v I__9931 (
            .O(N__53434),
            .I(N__53425));
    Span4Mux_v I__9930 (
            .O(N__53431),
            .I(N__53422));
    LocalMux I__9929 (
            .O(N__53428),
            .I(\ppm_encoder_1.N_268_i_i ));
    Odrv4 I__9928 (
            .O(N__53425),
            .I(\ppm_encoder_1.N_268_i_i ));
    Odrv4 I__9927 (
            .O(N__53422),
            .I(\ppm_encoder_1.N_268_i_i ));
    InMux I__9926 (
            .O(N__53415),
            .I(N__53412));
    LocalMux I__9925 (
            .O(N__53412),
            .I(N__53409));
    Span4Mux_h I__9924 (
            .O(N__53409),
            .I(N__53406));
    Odrv4 I__9923 (
            .O(N__53406),
            .I(\ppm_encoder_1.init_pulses_RNIFVPF5Z0Z_13 ));
    InMux I__9922 (
            .O(N__53403),
            .I(N__53400));
    LocalMux I__9921 (
            .O(N__53400),
            .I(\ppm_encoder_1.un2_throttle_iv_0_1_13 ));
    InMux I__9920 (
            .O(N__53397),
            .I(N__53394));
    LocalMux I__9919 (
            .O(N__53394),
            .I(\ppm_encoder_1.un2_throttle_iv_0_0_13 ));
    InMux I__9918 (
            .O(N__53391),
            .I(N__53385));
    InMux I__9917 (
            .O(N__53390),
            .I(N__53385));
    LocalMux I__9916 (
            .O(N__53385),
            .I(\ppm_encoder_1.elevator_RNIRHGEZ0Z_13 ));
    CascadeMux I__9915 (
            .O(N__53382),
            .I(N__53378));
    InMux I__9914 (
            .O(N__53381),
            .I(N__53373));
    InMux I__9913 (
            .O(N__53378),
            .I(N__53373));
    LocalMux I__9912 (
            .O(N__53373),
            .I(N__53369));
    InMux I__9911 (
            .O(N__53372),
            .I(N__53365));
    Span4Mux_v I__9910 (
            .O(N__53369),
            .I(N__53362));
    InMux I__9909 (
            .O(N__53368),
            .I(N__53359));
    LocalMux I__9908 (
            .O(N__53365),
            .I(\ppm_encoder_1.init_pulsesZ0Z_13 ));
    Odrv4 I__9907 (
            .O(N__53362),
            .I(\ppm_encoder_1.init_pulsesZ0Z_13 ));
    LocalMux I__9906 (
            .O(N__53359),
            .I(\ppm_encoder_1.init_pulsesZ0Z_13 ));
    CascadeMux I__9905 (
            .O(N__53352),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIHO7DZ0Z_0_cascade_ ));
    InMux I__9904 (
            .O(N__53349),
            .I(N__53346));
    LocalMux I__9903 (
            .O(N__53346),
            .I(\ppm_encoder_1.un2_throttle_iv_0_1_10 ));
    InMux I__9902 (
            .O(N__53343),
            .I(N__53340));
    LocalMux I__9901 (
            .O(N__53340),
            .I(N__53336));
    InMux I__9900 (
            .O(N__53339),
            .I(N__53333));
    Span4Mux_h I__9899 (
            .O(N__53336),
            .I(N__53329));
    LocalMux I__9898 (
            .O(N__53333),
            .I(N__53326));
    InMux I__9897 (
            .O(N__53332),
            .I(N__53323));
    Span4Mux_v I__9896 (
            .O(N__53329),
            .I(N__53318));
    Span4Mux_h I__9895 (
            .O(N__53326),
            .I(N__53318));
    LocalMux I__9894 (
            .O(N__53323),
            .I(\ppm_encoder_1.throttleZ0Z_2 ));
    Odrv4 I__9893 (
            .O(N__53318),
            .I(\ppm_encoder_1.throttleZ0Z_2 ));
    CascadeMux I__9892 (
            .O(N__53313),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIJQ7DZ0Z_1_cascade_ ));
    CascadeMux I__9891 (
            .O(N__53310),
            .I(\ppm_encoder_1.un2_throttle_iv_i_i_0_14_cascade_ ));
    CascadeMux I__9890 (
            .O(N__53307),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_14_cascade_ ));
    InMux I__9889 (
            .O(N__53304),
            .I(N__53301));
    LocalMux I__9888 (
            .O(N__53301),
            .I(N__53298));
    Odrv4 I__9887 (
            .O(N__53298),
            .I(\ppm_encoder_1.init_pulses_RNIE8336Z0Z_14 ));
    CascadeMux I__9886 (
            .O(N__53295),
            .I(\ppm_encoder_1.PPM_STATE_RNIV4V5Z0Z_1_cascade_ ));
    CascadeMux I__9885 (
            .O(N__53292),
            .I(N__53289));
    InMux I__9884 (
            .O(N__53289),
            .I(N__53286));
    LocalMux I__9883 (
            .O(N__53286),
            .I(N__53282));
    InMux I__9882 (
            .O(N__53285),
            .I(N__53279));
    Odrv12 I__9881 (
            .O(N__53282),
            .I(\ppm_encoder_1.N_269_i_i ));
    LocalMux I__9880 (
            .O(N__53279),
            .I(\ppm_encoder_1.N_269_i_i ));
    InMux I__9879 (
            .O(N__53274),
            .I(N__53271));
    LocalMux I__9878 (
            .O(N__53271),
            .I(\ppm_encoder_1.N_269_i ));
    InMux I__9877 (
            .O(N__53268),
            .I(N__53265));
    LocalMux I__9876 (
            .O(N__53265),
            .I(N__53262));
    Span4Mux_h I__9875 (
            .O(N__53262),
            .I(N__53259));
    Odrv4 I__9874 (
            .O(N__53259),
            .I(\ppm_encoder_1.counter24_0_I_57_c_RNIJMMDZ0 ));
    CascadeMux I__9873 (
            .O(N__53256),
            .I(N__53252));
    InMux I__9872 (
            .O(N__53255),
            .I(N__53248));
    InMux I__9871 (
            .O(N__53252),
            .I(N__53245));
    InMux I__9870 (
            .O(N__53251),
            .I(N__53242));
    LocalMux I__9869 (
            .O(N__53248),
            .I(\ppm_encoder_1.aileronZ0Z_1 ));
    LocalMux I__9868 (
            .O(N__53245),
            .I(\ppm_encoder_1.aileronZ0Z_1 ));
    LocalMux I__9867 (
            .O(N__53242),
            .I(\ppm_encoder_1.aileronZ0Z_1 ));
    CascadeMux I__9866 (
            .O(N__53235),
            .I(\ppm_encoder_1.pulses2count_9_0_0_0_3_cascade_ ));
    CascadeMux I__9865 (
            .O(N__53232),
            .I(N__53227));
    InMux I__9864 (
            .O(N__53231),
            .I(N__53223));
    InMux I__9863 (
            .O(N__53230),
            .I(N__53218));
    InMux I__9862 (
            .O(N__53227),
            .I(N__53218));
    InMux I__9861 (
            .O(N__53226),
            .I(N__53215));
    LocalMux I__9860 (
            .O(N__53223),
            .I(N__53212));
    LocalMux I__9859 (
            .O(N__53218),
            .I(N__53209));
    LocalMux I__9858 (
            .O(N__53215),
            .I(N__53206));
    Span4Mux_s1_v I__9857 (
            .O(N__53212),
            .I(N__53203));
    Span4Mux_h I__9856 (
            .O(N__53209),
            .I(N__53200));
    Odrv4 I__9855 (
            .O(N__53206),
            .I(\ppm_encoder_1.init_pulsesZ0Z_3 ));
    Odrv4 I__9854 (
            .O(N__53203),
            .I(\ppm_encoder_1.init_pulsesZ0Z_3 ));
    Odrv4 I__9853 (
            .O(N__53200),
            .I(\ppm_encoder_1.init_pulsesZ0Z_3 ));
    CascadeMux I__9852 (
            .O(N__53193),
            .I(\ppm_encoder_1.un2_throttle_iv_0_0_0_cascade_ ));
    InMux I__9851 (
            .O(N__53190),
            .I(N__53187));
    LocalMux I__9850 (
            .O(N__53187),
            .I(N__53184));
    Odrv12 I__9849 (
            .O(N__53184),
            .I(\ppm_encoder_1.throttle_RNI25564Z0Z_0 ));
    InMux I__9848 (
            .O(N__53181),
            .I(N__53178));
    LocalMux I__9847 (
            .O(N__53178),
            .I(\ppm_encoder_1.un2_throttle_iv_0_1_0 ));
    InMux I__9846 (
            .O(N__53175),
            .I(N__53172));
    LocalMux I__9845 (
            .O(N__53172),
            .I(\ppm_encoder_1.un2_throttle_iv_0_0_0 ));
    CascadeMux I__9844 (
            .O(N__53169),
            .I(\ppm_encoder_1.un2_throttle_iv_0_1_0_cascade_ ));
    InMux I__9843 (
            .O(N__53166),
            .I(N__53163));
    LocalMux I__9842 (
            .O(N__53163),
            .I(N__53160));
    Span4Mux_s3_v I__9841 (
            .O(N__53160),
            .I(N__53157));
    Span4Mux_v I__9840 (
            .O(N__53157),
            .I(N__53153));
    InMux I__9839 (
            .O(N__53156),
            .I(N__53150));
    Span4Mux_h I__9838 (
            .O(N__53153),
            .I(N__53145));
    LocalMux I__9837 (
            .O(N__53150),
            .I(N__53145));
    Span4Mux_h I__9836 (
            .O(N__53145),
            .I(N__53142));
    Odrv4 I__9835 (
            .O(N__53142),
            .I(throttle_order_0));
    InMux I__9834 (
            .O(N__53139),
            .I(N__53130));
    InMux I__9833 (
            .O(N__53138),
            .I(N__53130));
    InMux I__9832 (
            .O(N__53137),
            .I(N__53130));
    LocalMux I__9831 (
            .O(N__53130),
            .I(\ppm_encoder_1.aileronZ0Z_0 ));
    CascadeMux I__9830 (
            .O(N__53127),
            .I(N__53122));
    CascadeMux I__9829 (
            .O(N__53126),
            .I(N__53119));
    InMux I__9828 (
            .O(N__53125),
            .I(N__53112));
    InMux I__9827 (
            .O(N__53122),
            .I(N__53112));
    InMux I__9826 (
            .O(N__53119),
            .I(N__53112));
    LocalMux I__9825 (
            .O(N__53112),
            .I(\ppm_encoder_1.throttleZ0Z_0 ));
    InMux I__9824 (
            .O(N__53109),
            .I(N__53106));
    LocalMux I__9823 (
            .O(N__53106),
            .I(N__53102));
    InMux I__9822 (
            .O(N__53105),
            .I(N__53099));
    Span12Mux_h I__9821 (
            .O(N__53102),
            .I(N__53096));
    LocalMux I__9820 (
            .O(N__53099),
            .I(N__53093));
    Span12Mux_v I__9819 (
            .O(N__53096),
            .I(N__53090));
    Span4Mux_v I__9818 (
            .O(N__53093),
            .I(N__53087));
    Odrv12 I__9817 (
            .O(N__53090),
            .I(front_order_0));
    Odrv4 I__9816 (
            .O(N__53087),
            .I(front_order_0));
    CascadeMux I__9815 (
            .O(N__53082),
            .I(\ppm_encoder_1.un2_throttle_iv_0_2_11_cascade_ ));
    CascadeMux I__9814 (
            .O(N__53079),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_11_cascade_ ));
    InMux I__9813 (
            .O(N__53076),
            .I(N__53073));
    LocalMux I__9812 (
            .O(N__53073),
            .I(N__53070));
    Span4Mux_h I__9811 (
            .O(N__53070),
            .I(N__53067));
    Odrv4 I__9810 (
            .O(N__53067),
            .I(\ppm_encoder_1.init_pulses_RNI4JPF5Z0Z_11 ));
    CascadeMux I__9809 (
            .O(N__53064),
            .I(N__53059));
    InMux I__9808 (
            .O(N__53063),
            .I(N__53056));
    InMux I__9807 (
            .O(N__53062),
            .I(N__53050));
    InMux I__9806 (
            .O(N__53059),
            .I(N__53050));
    LocalMux I__9805 (
            .O(N__53056),
            .I(N__53047));
    CascadeMux I__9804 (
            .O(N__53055),
            .I(N__53044));
    LocalMux I__9803 (
            .O(N__53050),
            .I(N__53041));
    Span12Mux_h I__9802 (
            .O(N__53047),
            .I(N__53038));
    InMux I__9801 (
            .O(N__53044),
            .I(N__53035));
    Span4Mux_s1_v I__9800 (
            .O(N__53041),
            .I(N__53032));
    Odrv12 I__9799 (
            .O(N__53038),
            .I(\ppm_encoder_1.init_pulsesZ0Z_11 ));
    LocalMux I__9798 (
            .O(N__53035),
            .I(\ppm_encoder_1.init_pulsesZ0Z_11 ));
    Odrv4 I__9797 (
            .O(N__53032),
            .I(\ppm_encoder_1.init_pulsesZ0Z_11 ));
    CascadeMux I__9796 (
            .O(N__53025),
            .I(N__53022));
    InMux I__9795 (
            .O(N__53022),
            .I(N__53019));
    LocalMux I__9794 (
            .O(N__53019),
            .I(N__53016));
    Span4Mux_h I__9793 (
            .O(N__53016),
            .I(N__53012));
    InMux I__9792 (
            .O(N__53015),
            .I(N__53009));
    Odrv4 I__9791 (
            .O(N__53012),
            .I(\ppm_encoder_1.N_266_i_i ));
    LocalMux I__9790 (
            .O(N__53009),
            .I(\ppm_encoder_1.N_266_i_i ));
    InMux I__9789 (
            .O(N__53004),
            .I(N__53001));
    LocalMux I__9788 (
            .O(N__53001),
            .I(N__52998));
    Odrv12 I__9787 (
            .O(N__52998),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_4 ));
    InMux I__9786 (
            .O(N__52995),
            .I(N__52992));
    LocalMux I__9785 (
            .O(N__52992),
            .I(N__52989));
    Odrv4 I__9784 (
            .O(N__52989),
            .I(\ppm_encoder_1.un1_init_pulses_11_13 ));
    InMux I__9783 (
            .O(N__52986),
            .I(N__52983));
    LocalMux I__9782 (
            .O(N__52983),
            .I(N__52980));
    Span4Mux_h I__9781 (
            .O(N__52980),
            .I(N__52977));
    Odrv4 I__9780 (
            .O(N__52977),
            .I(\ppm_encoder_1.un1_init_pulses_10_13 ));
    InMux I__9779 (
            .O(N__52974),
            .I(N__52971));
    LocalMux I__9778 (
            .O(N__52971),
            .I(N__52968));
    Span4Mux_h I__9777 (
            .O(N__52968),
            .I(N__52965));
    Odrv4 I__9776 (
            .O(N__52965),
            .I(\ppm_encoder_1.un1_init_pulses_11_2 ));
    CascadeMux I__9775 (
            .O(N__52962),
            .I(N__52959));
    InMux I__9774 (
            .O(N__52959),
            .I(N__52956));
    LocalMux I__9773 (
            .O(N__52956),
            .I(N__52953));
    Span4Mux_s2_v I__9772 (
            .O(N__52953),
            .I(N__52950));
    Odrv4 I__9771 (
            .O(N__52950),
            .I(\ppm_encoder_1.un1_init_pulses_10_2 ));
    InMux I__9770 (
            .O(N__52947),
            .I(N__52938));
    InMux I__9769 (
            .O(N__52946),
            .I(N__52938));
    InMux I__9768 (
            .O(N__52945),
            .I(N__52935));
    InMux I__9767 (
            .O(N__52944),
            .I(N__52931));
    InMux I__9766 (
            .O(N__52943),
            .I(N__52928));
    LocalMux I__9765 (
            .O(N__52938),
            .I(N__52923));
    LocalMux I__9764 (
            .O(N__52935),
            .I(N__52923));
    InMux I__9763 (
            .O(N__52934),
            .I(N__52920));
    LocalMux I__9762 (
            .O(N__52931),
            .I(N__52917));
    LocalMux I__9761 (
            .O(N__52928),
            .I(N__52914));
    Span12Mux_s4_v I__9760 (
            .O(N__52923),
            .I(N__52905));
    LocalMux I__9759 (
            .O(N__52920),
            .I(N__52902));
    Span4Mux_h I__9758 (
            .O(N__52917),
            .I(N__52899));
    Span4Mux_h I__9757 (
            .O(N__52914),
            .I(N__52896));
    InMux I__9756 (
            .O(N__52913),
            .I(N__52893));
    InMux I__9755 (
            .O(N__52912),
            .I(N__52890));
    InMux I__9754 (
            .O(N__52911),
            .I(N__52881));
    InMux I__9753 (
            .O(N__52910),
            .I(N__52881));
    InMux I__9752 (
            .O(N__52909),
            .I(N__52881));
    InMux I__9751 (
            .O(N__52908),
            .I(N__52881));
    Odrv12 I__9750 (
            .O(N__52905),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1 ));
    Odrv4 I__9749 (
            .O(N__52902),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1 ));
    Odrv4 I__9748 (
            .O(N__52899),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1 ));
    Odrv4 I__9747 (
            .O(N__52896),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1 ));
    LocalMux I__9746 (
            .O(N__52893),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1 ));
    LocalMux I__9745 (
            .O(N__52890),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1 ));
    LocalMux I__9744 (
            .O(N__52881),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1 ));
    InMux I__9743 (
            .O(N__52866),
            .I(N__52862));
    CascadeMux I__9742 (
            .O(N__52865),
            .I(N__52859));
    LocalMux I__9741 (
            .O(N__52862),
            .I(N__52856));
    InMux I__9740 (
            .O(N__52859),
            .I(N__52853));
    Span4Mux_s3_v I__9739 (
            .O(N__52856),
            .I(N__52849));
    LocalMux I__9738 (
            .O(N__52853),
            .I(N__52846));
    InMux I__9737 (
            .O(N__52852),
            .I(N__52843));
    Span4Mux_h I__9736 (
            .O(N__52849),
            .I(N__52838));
    Span4Mux_h I__9735 (
            .O(N__52846),
            .I(N__52838));
    LocalMux I__9734 (
            .O(N__52843),
            .I(\ppm_encoder_1.elevatorZ0Z_3 ));
    Odrv4 I__9733 (
            .O(N__52838),
            .I(\ppm_encoder_1.elevatorZ0Z_3 ));
    CascadeMux I__9732 (
            .O(N__52833),
            .I(N__52830));
    InMux I__9731 (
            .O(N__52830),
            .I(N__52821));
    InMux I__9730 (
            .O(N__52829),
            .I(N__52821));
    InMux I__9729 (
            .O(N__52828),
            .I(N__52818));
    InMux I__9728 (
            .O(N__52827),
            .I(N__52814));
    InMux I__9727 (
            .O(N__52826),
            .I(N__52811));
    LocalMux I__9726 (
            .O(N__52821),
            .I(N__52806));
    LocalMux I__9725 (
            .O(N__52818),
            .I(N__52806));
    InMux I__9724 (
            .O(N__52817),
            .I(N__52803));
    LocalMux I__9723 (
            .O(N__52814),
            .I(N__52800));
    LocalMux I__9722 (
            .O(N__52811),
            .I(N__52797));
    Span4Mux_s1_v I__9721 (
            .O(N__52806),
            .I(N__52788));
    LocalMux I__9720 (
            .O(N__52803),
            .I(N__52783));
    Span4Mux_h I__9719 (
            .O(N__52800),
            .I(N__52783));
    Span4Mux_h I__9718 (
            .O(N__52797),
            .I(N__52780));
    InMux I__9717 (
            .O(N__52796),
            .I(N__52777));
    InMux I__9716 (
            .O(N__52795),
            .I(N__52772));
    InMux I__9715 (
            .O(N__52794),
            .I(N__52772));
    InMux I__9714 (
            .O(N__52793),
            .I(N__52765));
    InMux I__9713 (
            .O(N__52792),
            .I(N__52765));
    InMux I__9712 (
            .O(N__52791),
            .I(N__52765));
    Odrv4 I__9711 (
            .O(N__52788),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1 ));
    Odrv4 I__9710 (
            .O(N__52783),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1 ));
    Odrv4 I__9709 (
            .O(N__52780),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1 ));
    LocalMux I__9708 (
            .O(N__52777),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1 ));
    LocalMux I__9707 (
            .O(N__52772),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1 ));
    LocalMux I__9706 (
            .O(N__52765),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1 ));
    InMux I__9705 (
            .O(N__52752),
            .I(N__52748));
    InMux I__9704 (
            .O(N__52751),
            .I(N__52744));
    LocalMux I__9703 (
            .O(N__52748),
            .I(N__52741));
    InMux I__9702 (
            .O(N__52747),
            .I(N__52738));
    LocalMux I__9701 (
            .O(N__52744),
            .I(N__52735));
    Odrv12 I__9700 (
            .O(N__52741),
            .I(\pid_front.un10lto12 ));
    LocalMux I__9699 (
            .O(N__52738),
            .I(\pid_front.un10lto12 ));
    Odrv4 I__9698 (
            .O(N__52735),
            .I(\pid_front.un10lto12 ));
    InMux I__9697 (
            .O(N__52728),
            .I(N__52725));
    LocalMux I__9696 (
            .O(N__52725),
            .I(\pid_front.error_i_acumm16lto27_10 ));
    InMux I__9695 (
            .O(N__52722),
            .I(N__52719));
    LocalMux I__9694 (
            .O(N__52719),
            .I(N__52716));
    Odrv4 I__9693 (
            .O(N__52716),
            .I(\pid_front.error_i_acumm16lto27_9 ));
    CascadeMux I__9692 (
            .O(N__52713),
            .I(\pid_front.error_i_acumm16lto27_7_cascade_ ));
    InMux I__9691 (
            .O(N__52710),
            .I(N__52707));
    LocalMux I__9690 (
            .O(N__52707),
            .I(\pid_front.error_i_acumm16lto27_8 ));
    InMux I__9689 (
            .O(N__52704),
            .I(N__52701));
    LocalMux I__9688 (
            .O(N__52701),
            .I(N__52698));
    Odrv12 I__9687 (
            .O(N__52698),
            .I(\pid_front.error_i_acumm16lto27_13 ));
    InMux I__9686 (
            .O(N__52695),
            .I(N__52689));
    InMux I__9685 (
            .O(N__52694),
            .I(N__52689));
    LocalMux I__9684 (
            .O(N__52689),
            .I(\pid_front.error_i_acumm_preregZ0Z_22 ));
    CascadeMux I__9683 (
            .O(N__52686),
            .I(N__52683));
    InMux I__9682 (
            .O(N__52683),
            .I(N__52677));
    InMux I__9681 (
            .O(N__52682),
            .I(N__52677));
    LocalMux I__9680 (
            .O(N__52677),
            .I(\pid_front.error_i_acumm_preregZ0Z_24 ));
    InMux I__9679 (
            .O(N__52674),
            .I(N__52671));
    LocalMux I__9678 (
            .O(N__52671),
            .I(N__52666));
    InMux I__9677 (
            .O(N__52670),
            .I(N__52661));
    InMux I__9676 (
            .O(N__52669),
            .I(N__52661));
    Odrv12 I__9675 (
            .O(N__52666),
            .I(\pid_front.error_i_acumm_preregZ0Z_13 ));
    LocalMux I__9674 (
            .O(N__52661),
            .I(\pid_front.error_i_acumm_preregZ0Z_13 ));
    CascadeMux I__9673 (
            .O(N__52656),
            .I(\pid_front.un10lto27_8_cascade_ ));
    InMux I__9672 (
            .O(N__52653),
            .I(N__52650));
    LocalMux I__9671 (
            .O(N__52650),
            .I(\pid_front.un10lto27_11 ));
    CascadeMux I__9670 (
            .O(N__52647),
            .I(N__52644));
    InMux I__9669 (
            .O(N__52644),
            .I(N__52638));
    InMux I__9668 (
            .O(N__52643),
            .I(N__52638));
    LocalMux I__9667 (
            .O(N__52638),
            .I(\pid_front.error_i_acumm_preregZ0Z_26 ));
    InMux I__9666 (
            .O(N__52635),
            .I(N__52631));
    InMux I__9665 (
            .O(N__52634),
            .I(N__52627));
    LocalMux I__9664 (
            .O(N__52631),
            .I(N__52624));
    CascadeMux I__9663 (
            .O(N__52630),
            .I(N__52621));
    LocalMux I__9662 (
            .O(N__52627),
            .I(N__52618));
    Span4Mux_s3_v I__9661 (
            .O(N__52624),
            .I(N__52615));
    InMux I__9660 (
            .O(N__52621),
            .I(N__52612));
    Span4Mux_v I__9659 (
            .O(N__52618),
            .I(N__52609));
    Span4Mux_h I__9658 (
            .O(N__52615),
            .I(N__52606));
    LocalMux I__9657 (
            .O(N__52612),
            .I(\ppm_encoder_1.elevatorZ0Z_11 ));
    Odrv4 I__9656 (
            .O(N__52609),
            .I(\ppm_encoder_1.elevatorZ0Z_11 ));
    Odrv4 I__9655 (
            .O(N__52606),
            .I(\ppm_encoder_1.elevatorZ0Z_11 ));
    CascadeMux I__9654 (
            .O(N__52599),
            .I(\ppm_encoder_1.elevator_RNIPFGEZ0Z_11_cascade_ ));
    InMux I__9653 (
            .O(N__52596),
            .I(N__52593));
    LocalMux I__9652 (
            .O(N__52593),
            .I(\pid_front.error_d_reg_prev_esr_RNIQHN6Z0Z_1 ));
    InMux I__9651 (
            .O(N__52590),
            .I(N__52582));
    InMux I__9650 (
            .O(N__52589),
            .I(N__52571));
    InMux I__9649 (
            .O(N__52588),
            .I(N__52571));
    InMux I__9648 (
            .O(N__52587),
            .I(N__52571));
    InMux I__9647 (
            .O(N__52586),
            .I(N__52571));
    InMux I__9646 (
            .O(N__52585),
            .I(N__52571));
    LocalMux I__9645 (
            .O(N__52582),
            .I(\pid_front.error_d_regZ0Z_1 ));
    LocalMux I__9644 (
            .O(N__52571),
            .I(\pid_front.error_d_regZ0Z_1 ));
    InMux I__9643 (
            .O(N__52566),
            .I(N__52562));
    CascadeMux I__9642 (
            .O(N__52565),
            .I(N__52559));
    LocalMux I__9641 (
            .O(N__52562),
            .I(N__52554));
    InMux I__9640 (
            .O(N__52559),
            .I(N__52547));
    InMux I__9639 (
            .O(N__52558),
            .I(N__52547));
    InMux I__9638 (
            .O(N__52557),
            .I(N__52547));
    Odrv4 I__9637 (
            .O(N__52554),
            .I(\pid_front.error_d_reg_prevZ0Z_1 ));
    LocalMux I__9636 (
            .O(N__52547),
            .I(\pid_front.error_d_reg_prevZ0Z_1 ));
    CascadeMux I__9635 (
            .O(N__52542),
            .I(N__52538));
    CascadeMux I__9634 (
            .O(N__52541),
            .I(N__52535));
    InMux I__9633 (
            .O(N__52538),
            .I(N__52532));
    InMux I__9632 (
            .O(N__52535),
            .I(N__52529));
    LocalMux I__9631 (
            .O(N__52532),
            .I(\pid_front.error_i_acumm_preregZ0Z_21 ));
    LocalMux I__9630 (
            .O(N__52529),
            .I(\pid_front.error_i_acumm_preregZ0Z_21 ));
    InMux I__9629 (
            .O(N__52524),
            .I(N__52519));
    InMux I__9628 (
            .O(N__52523),
            .I(N__52516));
    InMux I__9627 (
            .O(N__52522),
            .I(N__52513));
    LocalMux I__9626 (
            .O(N__52519),
            .I(N__52506));
    LocalMux I__9625 (
            .O(N__52516),
            .I(N__52506));
    LocalMux I__9624 (
            .O(N__52513),
            .I(N__52506));
    Odrv4 I__9623 (
            .O(N__52506),
            .I(\pid_front.error_i_acumm_preregZ0Z_8 ));
    InMux I__9622 (
            .O(N__52503),
            .I(N__52497));
    InMux I__9621 (
            .O(N__52502),
            .I(N__52497));
    LocalMux I__9620 (
            .O(N__52497),
            .I(\pid_front.error_i_acumm_preregZ0Z_16 ));
    InMux I__9619 (
            .O(N__52494),
            .I(N__52491));
    LocalMux I__9618 (
            .O(N__52491),
            .I(N__52487));
    InMux I__9617 (
            .O(N__52490),
            .I(N__52484));
    Odrv4 I__9616 (
            .O(N__52487),
            .I(\pid_front.error_i_acumm_preregZ0Z_20 ));
    LocalMux I__9615 (
            .O(N__52484),
            .I(\pid_front.error_i_acumm_preregZ0Z_20 ));
    CascadeMux I__9614 (
            .O(N__52479),
            .I(N__52476));
    InMux I__9613 (
            .O(N__52476),
            .I(N__52473));
    LocalMux I__9612 (
            .O(N__52473),
            .I(N__52470));
    Span4Mux_h I__9611 (
            .O(N__52470),
            .I(N__52465));
    InMux I__9610 (
            .O(N__52469),
            .I(N__52460));
    InMux I__9609 (
            .O(N__52468),
            .I(N__52460));
    Odrv4 I__9608 (
            .O(N__52465),
            .I(\pid_front.error_i_acumm_preregZ0Z_6 ));
    LocalMux I__9607 (
            .O(N__52460),
            .I(\pid_front.error_i_acumm_preregZ0Z_6 ));
    InMux I__9606 (
            .O(N__52455),
            .I(N__52452));
    LocalMux I__9605 (
            .O(N__52452),
            .I(N__52448));
    InMux I__9604 (
            .O(N__52451),
            .I(N__52444));
    Span4Mux_v I__9603 (
            .O(N__52448),
            .I(N__52441));
    InMux I__9602 (
            .O(N__52447),
            .I(N__52438));
    LocalMux I__9601 (
            .O(N__52444),
            .I(N__52433));
    Span4Mux_v I__9600 (
            .O(N__52441),
            .I(N__52433));
    LocalMux I__9599 (
            .O(N__52438),
            .I(N__52428));
    Span4Mux_v I__9598 (
            .O(N__52433),
            .I(N__52428));
    Odrv4 I__9597 (
            .O(N__52428),
            .I(\pid_front.error_i_acumm_preregZ0Z_11 ));
    CascadeMux I__9596 (
            .O(N__52425),
            .I(N__52421));
    CascadeMux I__9595 (
            .O(N__52424),
            .I(N__52418));
    InMux I__9594 (
            .O(N__52421),
            .I(N__52401));
    InMux I__9593 (
            .O(N__52418),
            .I(N__52401));
    InMux I__9592 (
            .O(N__52417),
            .I(N__52401));
    InMux I__9591 (
            .O(N__52416),
            .I(N__52401));
    InMux I__9590 (
            .O(N__52415),
            .I(N__52401));
    InMux I__9589 (
            .O(N__52414),
            .I(N__52401));
    LocalMux I__9588 (
            .O(N__52401),
            .I(\pid_front.error_i_acumm_2_sqmuxa_1 ));
    InMux I__9587 (
            .O(N__52398),
            .I(N__52369));
    InMux I__9586 (
            .O(N__52397),
            .I(N__52369));
    InMux I__9585 (
            .O(N__52396),
            .I(N__52369));
    InMux I__9584 (
            .O(N__52395),
            .I(N__52369));
    InMux I__9583 (
            .O(N__52394),
            .I(N__52369));
    InMux I__9582 (
            .O(N__52393),
            .I(N__52369));
    InMux I__9581 (
            .O(N__52392),
            .I(N__52369));
    InMux I__9580 (
            .O(N__52391),
            .I(N__52369));
    InMux I__9579 (
            .O(N__52390),
            .I(N__52358));
    InMux I__9578 (
            .O(N__52389),
            .I(N__52358));
    InMux I__9577 (
            .O(N__52388),
            .I(N__52358));
    InMux I__9576 (
            .O(N__52387),
            .I(N__52358));
    InMux I__9575 (
            .O(N__52386),
            .I(N__52358));
    LocalMux I__9574 (
            .O(N__52369),
            .I(\pid_front.error_i_acumm_2_sqmuxa ));
    LocalMux I__9573 (
            .O(N__52358),
            .I(\pid_front.error_i_acumm_2_sqmuxa ));
    CascadeMux I__9572 (
            .O(N__52353),
            .I(\pid_front.error_p_reg_esr_RNI2BC9_0Z0Z_1_cascade_ ));
    CascadeMux I__9571 (
            .O(N__52350),
            .I(\pid_front.error_d_reg_prev_esr_RNIFSHOZ0Z_1_cascade_ ));
    InMux I__9570 (
            .O(N__52347),
            .I(N__52344));
    LocalMux I__9569 (
            .O(N__52344),
            .I(N__52341));
    Span4Mux_h I__9568 (
            .O(N__52341),
            .I(N__52338));
    Span4Mux_v I__9567 (
            .O(N__52338),
            .I(N__52335));
    Odrv4 I__9566 (
            .O(N__52335),
            .I(\pid_front.error_d_reg_prev_esr_RNID19M1Z0Z_1 ));
    InMux I__9565 (
            .O(N__52332),
            .I(N__52328));
    InMux I__9564 (
            .O(N__52331),
            .I(N__52325));
    LocalMux I__9563 (
            .O(N__52328),
            .I(N__52320));
    LocalMux I__9562 (
            .O(N__52325),
            .I(N__52320));
    Span12Mux_s8_v I__9561 (
            .O(N__52320),
            .I(N__52317));
    Odrv12 I__9560 (
            .O(N__52317),
            .I(\pid_front.error_p_reg_esr_RNIO4E8_0Z0Z_2 ));
    InMux I__9559 (
            .O(N__52314),
            .I(N__52311));
    LocalMux I__9558 (
            .O(N__52311),
            .I(\pid_front.error_d_reg_prev_esr_RNIFSHOZ0Z_1 ));
    CascadeMux I__9557 (
            .O(N__52308),
            .I(N__52305));
    InMux I__9556 (
            .O(N__52305),
            .I(N__52301));
    InMux I__9555 (
            .O(N__52304),
            .I(N__52298));
    LocalMux I__9554 (
            .O(N__52301),
            .I(N__52295));
    LocalMux I__9553 (
            .O(N__52298),
            .I(N__52292));
    Span4Mux_h I__9552 (
            .O(N__52295),
            .I(N__52287));
    Span4Mux_h I__9551 (
            .O(N__52292),
            .I(N__52287));
    Span4Mux_v I__9550 (
            .O(N__52287),
            .I(N__52284));
    Odrv4 I__9549 (
            .O(N__52284),
            .I(\pid_front.error_d_reg_prev_esr_RNI1JN71Z0Z_1 ));
    CascadeMux I__9548 (
            .O(N__52281),
            .I(N__52276));
    CascadeMux I__9547 (
            .O(N__52280),
            .I(N__52273));
    InMux I__9546 (
            .O(N__52279),
            .I(N__52270));
    InMux I__9545 (
            .O(N__52276),
            .I(N__52265));
    InMux I__9544 (
            .O(N__52273),
            .I(N__52265));
    LocalMux I__9543 (
            .O(N__52270),
            .I(\pid_front.error_p_regZ0Z_1 ));
    LocalMux I__9542 (
            .O(N__52265),
            .I(\pid_front.error_p_regZ0Z_1 ));
    InMux I__9541 (
            .O(N__52260),
            .I(N__52257));
    LocalMux I__9540 (
            .O(N__52257),
            .I(\pid_front.error_p_reg_esr_RNI2BC9Z0Z_1 ));
    InMux I__9539 (
            .O(N__52254),
            .I(N__52245));
    InMux I__9538 (
            .O(N__52253),
            .I(N__52245));
    InMux I__9537 (
            .O(N__52252),
            .I(N__52238));
    InMux I__9536 (
            .O(N__52251),
            .I(N__52238));
    InMux I__9535 (
            .O(N__52250),
            .I(N__52238));
    LocalMux I__9534 (
            .O(N__52245),
            .I(\pid_front.error_d_regZ0Z_0 ));
    LocalMux I__9533 (
            .O(N__52238),
            .I(\pid_front.error_d_regZ0Z_0 ));
    InMux I__9532 (
            .O(N__52233),
            .I(N__52225));
    InMux I__9531 (
            .O(N__52232),
            .I(N__52225));
    InMux I__9530 (
            .O(N__52231),
            .I(N__52220));
    InMux I__9529 (
            .O(N__52230),
            .I(N__52220));
    LocalMux I__9528 (
            .O(N__52225),
            .I(\pid_front.error_d_reg_prevZ0Z_0 ));
    LocalMux I__9527 (
            .O(N__52220),
            .I(\pid_front.error_d_reg_prevZ0Z_0 ));
    InMux I__9526 (
            .O(N__52215),
            .I(N__52211));
    InMux I__9525 (
            .O(N__52214),
            .I(N__52208));
    LocalMux I__9524 (
            .O(N__52211),
            .I(\pid_front.error_i_acumm_preregZ0Z_1 ));
    LocalMux I__9523 (
            .O(N__52208),
            .I(\pid_front.error_i_acumm_preregZ0Z_1 ));
    InMux I__9522 (
            .O(N__52203),
            .I(N__52200));
    LocalMux I__9521 (
            .O(N__52200),
            .I(N__52196));
    CascadeMux I__9520 (
            .O(N__52199),
            .I(N__52193));
    Span4Mux_h I__9519 (
            .O(N__52196),
            .I(N__52190));
    InMux I__9518 (
            .O(N__52193),
            .I(N__52187));
    Odrv4 I__9517 (
            .O(N__52190),
            .I(\pid_front.error_i_acumm_preregZ0Z_2 ));
    LocalMux I__9516 (
            .O(N__52187),
            .I(\pid_front.error_i_acumm_preregZ0Z_2 ));
    InMux I__9515 (
            .O(N__52182),
            .I(N__52178));
    InMux I__9514 (
            .O(N__52181),
            .I(N__52175));
    LocalMux I__9513 (
            .O(N__52178),
            .I(\pid_front.error_i_acumm16lto3 ));
    LocalMux I__9512 (
            .O(N__52175),
            .I(\pid_front.error_i_acumm16lto3 ));
    InMux I__9511 (
            .O(N__52170),
            .I(N__52167));
    LocalMux I__9510 (
            .O(N__52167),
            .I(\pid_front.error_i_acumm_prereg_esr_RNIV9S71Z0Z_12 ));
    CascadeMux I__9509 (
            .O(N__52164),
            .I(\pid_front.error_i_acumm_2_sqmuxa_1_cascade_ ));
    InMux I__9508 (
            .O(N__52161),
            .I(N__52158));
    LocalMux I__9507 (
            .O(N__52158),
            .I(\pid_front.error_i_acumm_prereg_esr_RNI0I2H5Z0Z_12 ));
    CascadeMux I__9506 (
            .O(N__52155),
            .I(\pid_front.error_i_acumm_2_sqmuxa_cascade_ ));
    InMux I__9505 (
            .O(N__52152),
            .I(N__52149));
    LocalMux I__9504 (
            .O(N__52149),
            .I(N__52145));
    InMux I__9503 (
            .O(N__52148),
            .I(N__52142));
    Span4Mux_h I__9502 (
            .O(N__52145),
            .I(N__52139));
    LocalMux I__9501 (
            .O(N__52142),
            .I(N__52135));
    Span4Mux_v I__9500 (
            .O(N__52139),
            .I(N__52132));
    InMux I__9499 (
            .O(N__52138),
            .I(N__52129));
    Span4Mux_h I__9498 (
            .O(N__52135),
            .I(N__52124));
    Span4Mux_v I__9497 (
            .O(N__52132),
            .I(N__52124));
    LocalMux I__9496 (
            .O(N__52129),
            .I(\pid_front.error_i_acumm_preregZ0Z_10 ));
    Odrv4 I__9495 (
            .O(N__52124),
            .I(\pid_front.error_i_acumm_preregZ0Z_10 ));
    CascadeMux I__9494 (
            .O(N__52119),
            .I(N__52116));
    InMux I__9493 (
            .O(N__52116),
            .I(N__52113));
    LocalMux I__9492 (
            .O(N__52113),
            .I(N__52110));
    Span4Mux_h I__9491 (
            .O(N__52110),
            .I(N__52105));
    InMux I__9490 (
            .O(N__52109),
            .I(N__52100));
    InMux I__9489 (
            .O(N__52108),
            .I(N__52100));
    Odrv4 I__9488 (
            .O(N__52105),
            .I(\pid_front.error_i_acumm_preregZ0Z_4 ));
    LocalMux I__9487 (
            .O(N__52100),
            .I(\pid_front.error_i_acumm_preregZ0Z_4 ));
    InMux I__9486 (
            .O(N__52095),
            .I(N__52092));
    LocalMux I__9485 (
            .O(N__52092),
            .I(N__52087));
    InMux I__9484 (
            .O(N__52091),
            .I(N__52082));
    InMux I__9483 (
            .O(N__52090),
            .I(N__52082));
    Span4Mux_h I__9482 (
            .O(N__52087),
            .I(N__52079));
    LocalMux I__9481 (
            .O(N__52082),
            .I(N__52076));
    Odrv4 I__9480 (
            .O(N__52079),
            .I(\pid_front.error_i_acumm_preregZ0Z_5 ));
    Odrv4 I__9479 (
            .O(N__52076),
            .I(\pid_front.error_i_acumm_preregZ0Z_5 ));
    InMux I__9478 (
            .O(N__52071),
            .I(N__52068));
    LocalMux I__9477 (
            .O(N__52068),
            .I(\dron_frame_decoder_1.drone_H_disp_front_10 ));
    CascadeMux I__9476 (
            .O(N__52065),
            .I(\pid_front.N_3_cascade_ ));
    CascadeMux I__9475 (
            .O(N__52062),
            .I(\pid_front.m2_0_03_3_i_0_cascade_ ));
    InMux I__9474 (
            .O(N__52059),
            .I(N__52056));
    LocalMux I__9473 (
            .O(N__52056),
            .I(\dron_frame_decoder_1.drone_H_disp_front_9 ));
    InMux I__9472 (
            .O(N__52053),
            .I(N__52050));
    LocalMux I__9471 (
            .O(N__52050),
            .I(N__52047));
    Span4Mux_h I__9470 (
            .O(N__52047),
            .I(N__52042));
    InMux I__9469 (
            .O(N__52046),
            .I(N__52037));
    InMux I__9468 (
            .O(N__52045),
            .I(N__52037));
    Odrv4 I__9467 (
            .O(N__52042),
            .I(\pid_front.error_i_acumm_preregZ0Z_7 ));
    LocalMux I__9466 (
            .O(N__52037),
            .I(\pid_front.error_i_acumm_preregZ0Z_7 ));
    InMux I__9465 (
            .O(N__52032),
            .I(N__52020));
    InMux I__9464 (
            .O(N__52031),
            .I(N__52020));
    InMux I__9463 (
            .O(N__52030),
            .I(N__52020));
    InMux I__9462 (
            .O(N__52029),
            .I(N__52020));
    LocalMux I__9461 (
            .O(N__52020),
            .I(\pid_front.error_i_acumm_3_sqmuxa ));
    InMux I__9460 (
            .O(N__52017),
            .I(N__52014));
    LocalMux I__9459 (
            .O(N__52014),
            .I(N__52009));
    InMux I__9458 (
            .O(N__52013),
            .I(N__52004));
    InMux I__9457 (
            .O(N__52012),
            .I(N__52004));
    Span4Mux_v I__9456 (
            .O(N__52009),
            .I(N__51999));
    LocalMux I__9455 (
            .O(N__52004),
            .I(N__51999));
    Span4Mux_h I__9454 (
            .O(N__51999),
            .I(N__51996));
    Span4Mux_v I__9453 (
            .O(N__51996),
            .I(N__51993));
    Odrv4 I__9452 (
            .O(N__51993),
            .I(\pid_front.error_i_acumm_preregZ0Z_9 ));
    CEMux I__9451 (
            .O(N__51990),
            .I(N__51987));
    LocalMux I__9450 (
            .O(N__51987),
            .I(N__51984));
    Span4Mux_v I__9449 (
            .O(N__51984),
            .I(N__51981));
    Span4Mux_v I__9448 (
            .O(N__51981),
            .I(N__51978));
    Odrv4 I__9447 (
            .O(N__51978),
            .I(\dron_frame_decoder_1.N_700_0 ));
    InMux I__9446 (
            .O(N__51975),
            .I(N__51972));
    LocalMux I__9445 (
            .O(N__51972),
            .I(\dron_frame_decoder_1.drone_H_disp_front_8 ));
    CascadeMux I__9444 (
            .O(N__51969),
            .I(\pid_front.un1_pid_prereg_0_7_cascade_ ));
    InMux I__9443 (
            .O(N__51966),
            .I(N__51963));
    LocalMux I__9442 (
            .O(N__51963),
            .I(N__51959));
    InMux I__9441 (
            .O(N__51962),
            .I(N__51956));
    Odrv12 I__9440 (
            .O(N__51959),
            .I(\pid_front.un1_pid_prereg_0_6 ));
    LocalMux I__9439 (
            .O(N__51956),
            .I(\pid_front.un1_pid_prereg_0_6 ));
    CascadeMux I__9438 (
            .O(N__51951),
            .I(N__51948));
    InMux I__9437 (
            .O(N__51948),
            .I(N__51945));
    LocalMux I__9436 (
            .O(N__51945),
            .I(N__51942));
    Odrv12 I__9435 (
            .O(N__51942),
            .I(\pid_front.error_p_reg_esr_RNIE7KM6Z0Z_17 ));
    CEMux I__9434 (
            .O(N__51939),
            .I(N__51936));
    LocalMux I__9433 (
            .O(N__51936),
            .I(N__51933));
    Span4Mux_v I__9432 (
            .O(N__51933),
            .I(N__51930));
    Odrv4 I__9431 (
            .O(N__51930),
            .I(\Commands_frame_decoder.source_CH3data_1_sqmuxa_0 ));
    InMux I__9430 (
            .O(N__51927),
            .I(N__51923));
    CascadeMux I__9429 (
            .O(N__51926),
            .I(N__51920));
    LocalMux I__9428 (
            .O(N__51923),
            .I(N__51916));
    InMux I__9427 (
            .O(N__51920),
            .I(N__51910));
    InMux I__9426 (
            .O(N__51919),
            .I(N__51910));
    Span4Mux_v I__9425 (
            .O(N__51916),
            .I(N__51907));
    InMux I__9424 (
            .O(N__51915),
            .I(N__51904));
    LocalMux I__9423 (
            .O(N__51910),
            .I(N__51901));
    Span4Mux_h I__9422 (
            .O(N__51907),
            .I(N__51896));
    LocalMux I__9421 (
            .O(N__51904),
            .I(N__51896));
    Odrv4 I__9420 (
            .O(N__51901),
            .I(\pid_front.error_p_reg_esr_RNIETB61_4Z0Z_13 ));
    Odrv4 I__9419 (
            .O(N__51896),
            .I(\pid_front.error_p_reg_esr_RNIETB61_4Z0Z_13 ));
    InMux I__9418 (
            .O(N__51891),
            .I(N__51888));
    LocalMux I__9417 (
            .O(N__51888),
            .I(\pid_front.error_d_reg_prev_esr_RNIOLN44Z0Z_12 ));
    CascadeMux I__9416 (
            .O(N__51885),
            .I(N__51882));
    InMux I__9415 (
            .O(N__51882),
            .I(N__51879));
    LocalMux I__9414 (
            .O(N__51879),
            .I(N__51875));
    InMux I__9413 (
            .O(N__51878),
            .I(N__51872));
    Span4Mux_v I__9412 (
            .O(N__51875),
            .I(N__51867));
    LocalMux I__9411 (
            .O(N__51872),
            .I(N__51867));
    Odrv4 I__9410 (
            .O(N__51867),
            .I(\pid_front.error_d_reg_prev_esr_RNI8SE96Z0Z_12 ));
    InMux I__9409 (
            .O(N__51864),
            .I(N__51861));
    LocalMux I__9408 (
            .O(N__51861),
            .I(N__51858));
    Span4Mux_v I__9407 (
            .O(N__51858),
            .I(N__51855));
    Span4Mux_v I__9406 (
            .O(N__51855),
            .I(N__51852));
    Span4Mux_h I__9405 (
            .O(N__51852),
            .I(N__51849));
    Odrv4 I__9404 (
            .O(N__51849),
            .I(\pid_front.error_p_reg_esr_RNIQ9C61Z0Z_17 ));
    CascadeMux I__9403 (
            .O(N__51846),
            .I(\pid_front.error_p_reg_esr_RNIQ9C61Z0Z_17_cascade_ ));
    InMux I__9402 (
            .O(N__51843),
            .I(N__51840));
    LocalMux I__9401 (
            .O(N__51840),
            .I(N__51837));
    Span4Mux_h I__9400 (
            .O(N__51837),
            .I(N__51833));
    InMux I__9399 (
            .O(N__51836),
            .I(N__51830));
    Span4Mux_v I__9398 (
            .O(N__51833),
            .I(N__51827));
    LocalMux I__9397 (
            .O(N__51830),
            .I(\pid_front.error_p_reg_esr_RNITCC61_0Z0Z_18 ));
    Odrv4 I__9396 (
            .O(N__51827),
            .I(\pid_front.error_p_reg_esr_RNITCC61_0Z0Z_18 ));
    InMux I__9395 (
            .O(N__51822),
            .I(N__51819));
    LocalMux I__9394 (
            .O(N__51819),
            .I(N__51816));
    Span4Mux_v I__9393 (
            .O(N__51816),
            .I(N__51813));
    Span4Mux_v I__9392 (
            .O(N__51813),
            .I(N__51809));
    InMux I__9391 (
            .O(N__51812),
            .I(N__51806));
    Odrv4 I__9390 (
            .O(N__51809),
            .I(\pid_front.un1_pid_prereg_0_4 ));
    LocalMux I__9389 (
            .O(N__51806),
            .I(\pid_front.un1_pid_prereg_0_4 ));
    InMux I__9388 (
            .O(N__51801),
            .I(N__51798));
    LocalMux I__9387 (
            .O(N__51798),
            .I(N__51795));
    Span4Mux_h I__9386 (
            .O(N__51795),
            .I(N__51792));
    Span4Mux_v I__9385 (
            .O(N__51792),
            .I(N__51788));
    InMux I__9384 (
            .O(N__51791),
            .I(N__51785));
    Odrv4 I__9383 (
            .O(N__51788),
            .I(\pid_front.un1_pid_prereg_0_5 ));
    LocalMux I__9382 (
            .O(N__51785),
            .I(\pid_front.un1_pid_prereg_0_5 ));
    CascadeMux I__9381 (
            .O(N__51780),
            .I(\pid_front.un1_pid_prereg_0_6_cascade_ ));
    InMux I__9380 (
            .O(N__51777),
            .I(N__51774));
    LocalMux I__9379 (
            .O(N__51774),
            .I(N__51771));
    Odrv12 I__9378 (
            .O(N__51771),
            .I(\pid_front.error_p_reg_esr_RNICS5DDZ0Z_16 ));
    InMux I__9377 (
            .O(N__51768),
            .I(N__51762));
    InMux I__9376 (
            .O(N__51767),
            .I(N__51762));
    LocalMux I__9375 (
            .O(N__51762),
            .I(N__51759));
    Span4Mux_v I__9374 (
            .O(N__51759),
            .I(N__51756));
    Span4Mux_h I__9373 (
            .O(N__51756),
            .I(N__51753));
    Odrv4 I__9372 (
            .O(N__51753),
            .I(\pid_front.error_p_regZ0Z_17 ));
    CascadeMux I__9371 (
            .O(N__51750),
            .I(N__51747));
    InMux I__9370 (
            .O(N__51747),
            .I(N__51741));
    InMux I__9369 (
            .O(N__51746),
            .I(N__51741));
    LocalMux I__9368 (
            .O(N__51741),
            .I(\pid_front.error_d_reg_prevZ0Z_17 ));
    InMux I__9367 (
            .O(N__51738),
            .I(N__51732));
    InMux I__9366 (
            .O(N__51737),
            .I(N__51732));
    LocalMux I__9365 (
            .O(N__51732),
            .I(N__51729));
    Span4Mux_h I__9364 (
            .O(N__51729),
            .I(N__51726));
    Span4Mux_v I__9363 (
            .O(N__51726),
            .I(N__51723));
    Odrv4 I__9362 (
            .O(N__51723),
            .I(\pid_front.error_p_reg_esr_RNIQ9C61_0Z0Z_17 ));
    InMux I__9361 (
            .O(N__51720),
            .I(N__51716));
    CascadeMux I__9360 (
            .O(N__51719),
            .I(N__51713));
    LocalMux I__9359 (
            .O(N__51716),
            .I(N__51710));
    InMux I__9358 (
            .O(N__51713),
            .I(N__51707));
    Span4Mux_v I__9357 (
            .O(N__51710),
            .I(N__51704));
    LocalMux I__9356 (
            .O(N__51707),
            .I(N__51701));
    Odrv4 I__9355 (
            .O(N__51704),
            .I(\pid_front.error_p_reg_esr_RNI0GC61_0Z0Z_19 ));
    Odrv4 I__9354 (
            .O(N__51701),
            .I(\pid_front.error_p_reg_esr_RNI0GC61_0Z0Z_19 ));
    InMux I__9353 (
            .O(N__51696),
            .I(N__51693));
    LocalMux I__9352 (
            .O(N__51693),
            .I(N__51689));
    InMux I__9351 (
            .O(N__51692),
            .I(N__51686));
    Odrv12 I__9350 (
            .O(N__51689),
            .I(\pid_front.un1_pid_prereg_0_7 ));
    LocalMux I__9349 (
            .O(N__51686),
            .I(\pid_front.un1_pid_prereg_0_7 ));
    InMux I__9348 (
            .O(N__51681),
            .I(N__51675));
    InMux I__9347 (
            .O(N__51680),
            .I(N__51675));
    LocalMux I__9346 (
            .O(N__51675),
            .I(N__51672));
    Span4Mux_h I__9345 (
            .O(N__51672),
            .I(N__51669));
    Span4Mux_h I__9344 (
            .O(N__51669),
            .I(N__51666));
    Span4Mux_h I__9343 (
            .O(N__51666),
            .I(N__51663));
    Odrv4 I__9342 (
            .O(N__51663),
            .I(\pid_front.error_p_regZ0Z_2 ));
    InMux I__9341 (
            .O(N__51660),
            .I(N__51654));
    InMux I__9340 (
            .O(N__51659),
            .I(N__51654));
    LocalMux I__9339 (
            .O(N__51654),
            .I(\pid_front.error_d_reg_prevZ0Z_2 ));
    InMux I__9338 (
            .O(N__51651),
            .I(N__51645));
    InMux I__9337 (
            .O(N__51650),
            .I(N__51645));
    LocalMux I__9336 (
            .O(N__51645),
            .I(N__51642));
    Span4Mux_h I__9335 (
            .O(N__51642),
            .I(N__51639));
    Span4Mux_h I__9334 (
            .O(N__51639),
            .I(N__51636));
    Odrv4 I__9333 (
            .O(N__51636),
            .I(\pid_front.error_p_regZ0Z_3 ));
    InMux I__9332 (
            .O(N__51633),
            .I(N__51627));
    InMux I__9331 (
            .O(N__51632),
            .I(N__51627));
    LocalMux I__9330 (
            .O(N__51627),
            .I(\pid_front.error_d_reg_prevZ0Z_3 ));
    InMux I__9329 (
            .O(N__51624),
            .I(N__51618));
    InMux I__9328 (
            .O(N__51623),
            .I(N__51618));
    LocalMux I__9327 (
            .O(N__51618),
            .I(N__51615));
    Span4Mux_h I__9326 (
            .O(N__51615),
            .I(N__51612));
    Odrv4 I__9325 (
            .O(N__51612),
            .I(\pid_front.error_p_reg_esr_RNIR7E8Z0Z_3 ));
    InMux I__9324 (
            .O(N__51609),
            .I(N__51606));
    LocalMux I__9323 (
            .O(N__51606),
            .I(N__51602));
    InMux I__9322 (
            .O(N__51605),
            .I(N__51599));
    Span4Mux_h I__9321 (
            .O(N__51602),
            .I(N__51596));
    LocalMux I__9320 (
            .O(N__51599),
            .I(N__51593));
    Span4Mux_v I__9319 (
            .O(N__51596),
            .I(N__51590));
    Span4Mux_h I__9318 (
            .O(N__51593),
            .I(N__51587));
    Sp12to4 I__9317 (
            .O(N__51590),
            .I(N__51584));
    Span4Mux_v I__9316 (
            .O(N__51587),
            .I(N__51581));
    Odrv12 I__9315 (
            .O(N__51584),
            .I(\pid_alt.error_p_regZ0Z_15 ));
    Odrv4 I__9314 (
            .O(N__51581),
            .I(\pid_alt.error_p_regZ0Z_15 ));
    InMux I__9313 (
            .O(N__51576),
            .I(N__51570));
    InMux I__9312 (
            .O(N__51575),
            .I(N__51570));
    LocalMux I__9311 (
            .O(N__51570),
            .I(N__51567));
    Span4Mux_v I__9310 (
            .O(N__51567),
            .I(N__51564));
    Span4Mux_h I__9309 (
            .O(N__51564),
            .I(N__51561));
    Span4Mux_h I__9308 (
            .O(N__51561),
            .I(N__51558));
    Odrv4 I__9307 (
            .O(N__51558),
            .I(\pid_alt.error_d_reg_prev_esr_RNISPHMZ0Z_15 ));
    InMux I__9306 (
            .O(N__51555),
            .I(N__51548));
    InMux I__9305 (
            .O(N__51554),
            .I(N__51548));
    InMux I__9304 (
            .O(N__51553),
            .I(N__51545));
    LocalMux I__9303 (
            .O(N__51548),
            .I(N__51542));
    LocalMux I__9302 (
            .O(N__51545),
            .I(N__51539));
    Span4Mux_v I__9301 (
            .O(N__51542),
            .I(N__51536));
    Span4Mux_v I__9300 (
            .O(N__51539),
            .I(N__51533));
    Span4Mux_h I__9299 (
            .O(N__51536),
            .I(N__51530));
    Span4Mux_h I__9298 (
            .O(N__51533),
            .I(N__51525));
    Span4Mux_h I__9297 (
            .O(N__51530),
            .I(N__51525));
    Span4Mux_v I__9296 (
            .O(N__51525),
            .I(N__51522));
    Span4Mux_v I__9295 (
            .O(N__51522),
            .I(N__51519));
    Odrv4 I__9294 (
            .O(N__51519),
            .I(\pid_alt.error_d_regZ0Z_15 ));
    InMux I__9293 (
            .O(N__51516),
            .I(N__51513));
    LocalMux I__9292 (
            .O(N__51513),
            .I(N__51510));
    Span4Mux_h I__9291 (
            .O(N__51510),
            .I(N__51506));
    InMux I__9290 (
            .O(N__51509),
            .I(N__51503));
    Span4Mux_h I__9289 (
            .O(N__51506),
            .I(N__51500));
    LocalMux I__9288 (
            .O(N__51503),
            .I(\pid_alt.error_d_reg_prevZ0Z_15 ));
    Odrv4 I__9287 (
            .O(N__51500),
            .I(\pid_alt.error_d_reg_prevZ0Z_15 ));
    CEMux I__9286 (
            .O(N__51495),
            .I(N__51423));
    CEMux I__9285 (
            .O(N__51494),
            .I(N__51423));
    CEMux I__9284 (
            .O(N__51493),
            .I(N__51423));
    CEMux I__9283 (
            .O(N__51492),
            .I(N__51423));
    CEMux I__9282 (
            .O(N__51491),
            .I(N__51423));
    CEMux I__9281 (
            .O(N__51490),
            .I(N__51423));
    CEMux I__9280 (
            .O(N__51489),
            .I(N__51423));
    CEMux I__9279 (
            .O(N__51488),
            .I(N__51423));
    CEMux I__9278 (
            .O(N__51487),
            .I(N__51423));
    CEMux I__9277 (
            .O(N__51486),
            .I(N__51423));
    CEMux I__9276 (
            .O(N__51485),
            .I(N__51423));
    CEMux I__9275 (
            .O(N__51484),
            .I(N__51423));
    CEMux I__9274 (
            .O(N__51483),
            .I(N__51423));
    CEMux I__9273 (
            .O(N__51482),
            .I(N__51423));
    CEMux I__9272 (
            .O(N__51481),
            .I(N__51423));
    CEMux I__9271 (
            .O(N__51480),
            .I(N__51423));
    CEMux I__9270 (
            .O(N__51479),
            .I(N__51423));
    CEMux I__9269 (
            .O(N__51478),
            .I(N__51423));
    CEMux I__9268 (
            .O(N__51477),
            .I(N__51423));
    CEMux I__9267 (
            .O(N__51476),
            .I(N__51423));
    CEMux I__9266 (
            .O(N__51475),
            .I(N__51423));
    CEMux I__9265 (
            .O(N__51474),
            .I(N__51423));
    CEMux I__9264 (
            .O(N__51473),
            .I(N__51423));
    CEMux I__9263 (
            .O(N__51472),
            .I(N__51423));
    GlobalMux I__9262 (
            .O(N__51423),
            .I(N__51420));
    gio2CtrlBuf I__9261 (
            .O(N__51420),
            .I(\pid_alt.state_0_g_0 ));
    IoInMux I__9260 (
            .O(N__51417),
            .I(N__51414));
    LocalMux I__9259 (
            .O(N__51414),
            .I(N__51411));
    Span12Mux_s3_v I__9258 (
            .O(N__51411),
            .I(N__51408));
    Odrv12 I__9257 (
            .O(N__51408),
            .I(\pid_front.state_RNIM14NZ0Z_0 ));
    InMux I__9256 (
            .O(N__51405),
            .I(N__51402));
    LocalMux I__9255 (
            .O(N__51402),
            .I(N__51399));
    Odrv4 I__9254 (
            .O(N__51399),
            .I(\pid_front.state_RNIVIRQZ0Z_0 ));
    CascadeMux I__9253 (
            .O(N__51396),
            .I(N__51393));
    InMux I__9252 (
            .O(N__51393),
            .I(N__51390));
    LocalMux I__9251 (
            .O(N__51390),
            .I(N__51387));
    Span4Mux_h I__9250 (
            .O(N__51387),
            .I(N__51384));
    Odrv4 I__9249 (
            .O(N__51384),
            .I(\pid_front.error_p_reg_esr_RNI3I672Z0Z_2 ));
    InMux I__9248 (
            .O(N__51381),
            .I(N__51378));
    LocalMux I__9247 (
            .O(N__51378),
            .I(\pid_front.error_p_reg_esr_RNIO4E8Z0Z_2 ));
    CascadeMux I__9246 (
            .O(N__51375),
            .I(\pid_front.error_p_reg_esr_RNIO4E8Z0Z_2_cascade_ ));
    InMux I__9245 (
            .O(N__51372),
            .I(N__51368));
    CascadeMux I__9244 (
            .O(N__51371),
            .I(N__51365));
    LocalMux I__9243 (
            .O(N__51368),
            .I(N__51362));
    InMux I__9242 (
            .O(N__51365),
            .I(N__51359));
    Span4Mux_v I__9241 (
            .O(N__51362),
            .I(N__51356));
    LocalMux I__9240 (
            .O(N__51359),
            .I(N__51353));
    Odrv4 I__9239 (
            .O(N__51356),
            .I(\pid_front.error_p_reg_esr_RNI2VEVZ0Z_2 ));
    Odrv4 I__9238 (
            .O(N__51353),
            .I(\pid_front.error_p_reg_esr_RNI2VEVZ0Z_2 ));
    InMux I__9237 (
            .O(N__51348),
            .I(N__51342));
    InMux I__9236 (
            .O(N__51347),
            .I(N__51342));
    LocalMux I__9235 (
            .O(N__51342),
            .I(\pid_front.error_p_reg_esr_RNIR7E8_0Z0Z_3 ));
    InMux I__9234 (
            .O(N__51339),
            .I(N__51336));
    LocalMux I__9233 (
            .O(N__51336),
            .I(N__51333));
    Span4Mux_v I__9232 (
            .O(N__51333),
            .I(N__51330));
    Span4Mux_h I__9231 (
            .O(N__51330),
            .I(N__51327));
    Span4Mux_v I__9230 (
            .O(N__51327),
            .I(N__51324));
    Sp12to4 I__9229 (
            .O(N__51324),
            .I(N__51321));
    Odrv12 I__9228 (
            .O(N__51321),
            .I(\Commands_frame_decoder.source_CH3data_1_sqmuxa ));
    InMux I__9227 (
            .O(N__51318),
            .I(N__51315));
    LocalMux I__9226 (
            .O(N__51315),
            .I(N__51311));
    InMux I__9225 (
            .O(N__51314),
            .I(N__51308));
    Span12Mux_s1_h I__9224 (
            .O(N__51311),
            .I(N__51305));
    LocalMux I__9223 (
            .O(N__51308),
            .I(N__51302));
    Span12Mux_v I__9222 (
            .O(N__51305),
            .I(N__51299));
    Span12Mux_v I__9221 (
            .O(N__51302),
            .I(N__51296));
    Span12Mux_h I__9220 (
            .O(N__51299),
            .I(N__51291));
    Span12Mux_h I__9219 (
            .O(N__51296),
            .I(N__51291));
    Odrv12 I__9218 (
            .O(N__51291),
            .I(xy_kp_0));
    InMux I__9217 (
            .O(N__51288),
            .I(N__51285));
    LocalMux I__9216 (
            .O(N__51285),
            .I(N__51281));
    InMux I__9215 (
            .O(N__51284),
            .I(N__51278));
    Span4Mux_s0_h I__9214 (
            .O(N__51281),
            .I(N__51275));
    LocalMux I__9213 (
            .O(N__51278),
            .I(N__51272));
    Span4Mux_h I__9212 (
            .O(N__51275),
            .I(N__51269));
    Span4Mux_h I__9211 (
            .O(N__51272),
            .I(N__51266));
    Span4Mux_h I__9210 (
            .O(N__51269),
            .I(N__51263));
    Span4Mux_h I__9209 (
            .O(N__51266),
            .I(N__51260));
    Span4Mux_h I__9208 (
            .O(N__51263),
            .I(N__51257));
    Span4Mux_h I__9207 (
            .O(N__51260),
            .I(N__51254));
    Odrv4 I__9206 (
            .O(N__51257),
            .I(xy_kp_2));
    Odrv4 I__9205 (
            .O(N__51254),
            .I(xy_kp_2));
    InMux I__9204 (
            .O(N__51249),
            .I(N__51246));
    LocalMux I__9203 (
            .O(N__51246),
            .I(N__51243));
    Span4Mux_s2_h I__9202 (
            .O(N__51243),
            .I(N__51239));
    InMux I__9201 (
            .O(N__51242),
            .I(N__51236));
    Span4Mux_v I__9200 (
            .O(N__51239),
            .I(N__51233));
    LocalMux I__9199 (
            .O(N__51236),
            .I(N__51230));
    Span4Mux_h I__9198 (
            .O(N__51233),
            .I(N__51227));
    Span12Mux_v I__9197 (
            .O(N__51230),
            .I(N__51224));
    Span4Mux_h I__9196 (
            .O(N__51227),
            .I(N__51221));
    Span12Mux_h I__9195 (
            .O(N__51224),
            .I(N__51218));
    Odrv4 I__9194 (
            .O(N__51221),
            .I(xy_kp_3));
    Odrv12 I__9193 (
            .O(N__51218),
            .I(xy_kp_3));
    InMux I__9192 (
            .O(N__51213),
            .I(N__51210));
    LocalMux I__9191 (
            .O(N__51210),
            .I(N__51206));
    InMux I__9190 (
            .O(N__51209),
            .I(N__51203));
    Span4Mux_v I__9189 (
            .O(N__51206),
            .I(N__51200));
    LocalMux I__9188 (
            .O(N__51203),
            .I(N__51197));
    Sp12to4 I__9187 (
            .O(N__51200),
            .I(N__51194));
    Span12Mux_v I__9186 (
            .O(N__51197),
            .I(N__51191));
    Span12Mux_h I__9185 (
            .O(N__51194),
            .I(N__51186));
    Span12Mux_h I__9184 (
            .O(N__51191),
            .I(N__51186));
    Odrv12 I__9183 (
            .O(N__51186),
            .I(xy_kp_7));
    InMux I__9182 (
            .O(N__51183),
            .I(N__51180));
    LocalMux I__9181 (
            .O(N__51180),
            .I(N__51176));
    InMux I__9180 (
            .O(N__51179),
            .I(N__51173));
    Odrv4 I__9179 (
            .O(N__51176),
            .I(\dron_frame_decoder_1.state_RNI4N6KZ0Z_2 ));
    LocalMux I__9178 (
            .O(N__51173),
            .I(\dron_frame_decoder_1.state_RNI4N6KZ0Z_2 ));
    InMux I__9177 (
            .O(N__51168),
            .I(N__51161));
    InMux I__9176 (
            .O(N__51167),
            .I(N__51161));
    InMux I__9175 (
            .O(N__51166),
            .I(N__51158));
    LocalMux I__9174 (
            .O(N__51161),
            .I(N__51151));
    LocalMux I__9173 (
            .O(N__51158),
            .I(N__51148));
    InMux I__9172 (
            .O(N__51157),
            .I(N__51143));
    InMux I__9171 (
            .O(N__51156),
            .I(N__51143));
    InMux I__9170 (
            .O(N__51155),
            .I(N__51138));
    InMux I__9169 (
            .O(N__51154),
            .I(N__51138));
    Span4Mux_v I__9168 (
            .O(N__51151),
            .I(N__51135));
    Span4Mux_v I__9167 (
            .O(N__51148),
            .I(N__51128));
    LocalMux I__9166 (
            .O(N__51143),
            .I(N__51128));
    LocalMux I__9165 (
            .O(N__51138),
            .I(N__51128));
    Odrv4 I__9164 (
            .O(N__51135),
            .I(\dron_frame_decoder_1.N_218 ));
    Odrv4 I__9163 (
            .O(N__51128),
            .I(\dron_frame_decoder_1.N_218 ));
    InMux I__9162 (
            .O(N__51123),
            .I(N__51120));
    LocalMux I__9161 (
            .O(N__51120),
            .I(\dron_frame_decoder_1.state_RNI6P6KZ0Z_4 ));
    CascadeMux I__9160 (
            .O(N__51117),
            .I(N__51114));
    InMux I__9159 (
            .O(N__51114),
            .I(N__51109));
    InMux I__9158 (
            .O(N__51113),
            .I(N__51106));
    InMux I__9157 (
            .O(N__51112),
            .I(N__51103));
    LocalMux I__9156 (
            .O(N__51109),
            .I(N__51098));
    LocalMux I__9155 (
            .O(N__51106),
            .I(N__51098));
    LocalMux I__9154 (
            .O(N__51103),
            .I(\dron_frame_decoder_1.stateZ0Z_7 ));
    Odrv4 I__9153 (
            .O(N__51098),
            .I(\dron_frame_decoder_1.stateZ0Z_7 ));
    InMux I__9152 (
            .O(N__51093),
            .I(N__51090));
    LocalMux I__9151 (
            .O(N__51090),
            .I(N__51087));
    Sp12to4 I__9150 (
            .O(N__51087),
            .I(N__51084));
    Odrv12 I__9149 (
            .O(N__51084),
            .I(\pid_front.error_i_acumm_prereg_esr_RNIRU7I_0Z0Z_10 ));
    CascadeMux I__9148 (
            .O(N__51081),
            .I(\dron_frame_decoder_1.state_ns_0_i_a2_0_2_3_cascade_ ));
    CascadeMux I__9147 (
            .O(N__51078),
            .I(N__51074));
    InMux I__9146 (
            .O(N__51077),
            .I(N__51068));
    InMux I__9145 (
            .O(N__51074),
            .I(N__51068));
    InMux I__9144 (
            .O(N__51073),
            .I(N__51065));
    LocalMux I__9143 (
            .O(N__51068),
            .I(N__51062));
    LocalMux I__9142 (
            .O(N__51065),
            .I(N__51057));
    Span4Mux_h I__9141 (
            .O(N__51062),
            .I(N__51057));
    Odrv4 I__9140 (
            .O(N__51057),
            .I(\dron_frame_decoder_1.stateZ0Z_3 ));
    InMux I__9139 (
            .O(N__51054),
            .I(N__51051));
    LocalMux I__9138 (
            .O(N__51051),
            .I(\dron_frame_decoder_1.N_230_5 ));
    InMux I__9137 (
            .O(N__51048),
            .I(N__51045));
    LocalMux I__9136 (
            .O(N__51045),
            .I(\dron_frame_decoder_1.state_ns_0_i_a2_0_3_3 ));
    InMux I__9135 (
            .O(N__51042),
            .I(N__51037));
    InMux I__9134 (
            .O(N__51041),
            .I(N__51032));
    InMux I__9133 (
            .O(N__51040),
            .I(N__51032));
    LocalMux I__9132 (
            .O(N__51037),
            .I(\dron_frame_decoder_1.stateZ0Z_1 ));
    LocalMux I__9131 (
            .O(N__51032),
            .I(\dron_frame_decoder_1.stateZ0Z_1 ));
    CascadeMux I__9130 (
            .O(N__51027),
            .I(N__51024));
    InMux I__9129 (
            .O(N__51024),
            .I(N__51021));
    LocalMux I__9128 (
            .O(N__51021),
            .I(\dron_frame_decoder_1.N_200 ));
    InMux I__9127 (
            .O(N__51018),
            .I(N__51010));
    InMux I__9126 (
            .O(N__51017),
            .I(N__51010));
    InMux I__9125 (
            .O(N__51016),
            .I(N__51005));
    InMux I__9124 (
            .O(N__51015),
            .I(N__51005));
    LocalMux I__9123 (
            .O(N__51010),
            .I(\dron_frame_decoder_1.stateZ0Z_0 ));
    LocalMux I__9122 (
            .O(N__51005),
            .I(\dron_frame_decoder_1.stateZ0Z_0 ));
    InMux I__9121 (
            .O(N__51000),
            .I(N__50997));
    LocalMux I__9120 (
            .O(N__50997),
            .I(\dron_frame_decoder_1.state_ns_i_a2_0_1_0 ));
    CascadeMux I__9119 (
            .O(N__50994),
            .I(N__50987));
    InMux I__9118 (
            .O(N__50993),
            .I(N__50983));
    InMux I__9117 (
            .O(N__50992),
            .I(N__50978));
    InMux I__9116 (
            .O(N__50991),
            .I(N__50978));
    InMux I__9115 (
            .O(N__50990),
            .I(N__50971));
    InMux I__9114 (
            .O(N__50987),
            .I(N__50971));
    InMux I__9113 (
            .O(N__50986),
            .I(N__50971));
    LocalMux I__9112 (
            .O(N__50983),
            .I(\dron_frame_decoder_1.stateZ0Z_6 ));
    LocalMux I__9111 (
            .O(N__50978),
            .I(\dron_frame_decoder_1.stateZ0Z_6 ));
    LocalMux I__9110 (
            .O(N__50971),
            .I(\dron_frame_decoder_1.stateZ0Z_6 ));
    InMux I__9109 (
            .O(N__50964),
            .I(N__50961));
    LocalMux I__9108 (
            .O(N__50961),
            .I(N__50955));
    InMux I__9107 (
            .O(N__50960),
            .I(N__50948));
    InMux I__9106 (
            .O(N__50959),
            .I(N__50948));
    InMux I__9105 (
            .O(N__50958),
            .I(N__50948));
    Span4Mux_v I__9104 (
            .O(N__50955),
            .I(N__50937));
    LocalMux I__9103 (
            .O(N__50948),
            .I(N__50937));
    InMux I__9102 (
            .O(N__50947),
            .I(N__50930));
    InMux I__9101 (
            .O(N__50946),
            .I(N__50930));
    InMux I__9100 (
            .O(N__50945),
            .I(N__50923));
    InMux I__9099 (
            .O(N__50944),
            .I(N__50923));
    InMux I__9098 (
            .O(N__50943),
            .I(N__50918));
    InMux I__9097 (
            .O(N__50942),
            .I(N__50918));
    Span4Mux_h I__9096 (
            .O(N__50937),
            .I(N__50915));
    InMux I__9095 (
            .O(N__50936),
            .I(N__50910));
    InMux I__9094 (
            .O(N__50935),
            .I(N__50910));
    LocalMux I__9093 (
            .O(N__50930),
            .I(N__50907));
    InMux I__9092 (
            .O(N__50929),
            .I(N__50904));
    InMux I__9091 (
            .O(N__50928),
            .I(N__50901));
    LocalMux I__9090 (
            .O(N__50923),
            .I(uart_drone_data_rdy));
    LocalMux I__9089 (
            .O(N__50918),
            .I(uart_drone_data_rdy));
    Odrv4 I__9088 (
            .O(N__50915),
            .I(uart_drone_data_rdy));
    LocalMux I__9087 (
            .O(N__50910),
            .I(uart_drone_data_rdy));
    Odrv4 I__9086 (
            .O(N__50907),
            .I(uart_drone_data_rdy));
    LocalMux I__9085 (
            .O(N__50904),
            .I(uart_drone_data_rdy));
    LocalMux I__9084 (
            .O(N__50901),
            .I(uart_drone_data_rdy));
    CascadeMux I__9083 (
            .O(N__50886),
            .I(N__50883));
    InMux I__9082 (
            .O(N__50883),
            .I(N__50880));
    LocalMux I__9081 (
            .O(N__50880),
            .I(N__50877));
    Odrv4 I__9080 (
            .O(N__50877),
            .I(\uart_drone.CO0 ));
    InMux I__9079 (
            .O(N__50874),
            .I(N__50868));
    InMux I__9078 (
            .O(N__50873),
            .I(N__50868));
    LocalMux I__9077 (
            .O(N__50868),
            .I(N__50865));
    Odrv4 I__9076 (
            .O(N__50865),
            .I(\uart_drone.un1_state_7_0 ));
    CascadeMux I__9075 (
            .O(N__50862),
            .I(N__50859));
    InMux I__9074 (
            .O(N__50859),
            .I(N__50854));
    InMux I__9073 (
            .O(N__50858),
            .I(N__50851));
    InMux I__9072 (
            .O(N__50857),
            .I(N__50848));
    LocalMux I__9071 (
            .O(N__50854),
            .I(N__50843));
    LocalMux I__9070 (
            .O(N__50851),
            .I(N__50843));
    LocalMux I__9069 (
            .O(N__50848),
            .I(\uart_drone.N_152 ));
    Odrv4 I__9068 (
            .O(N__50843),
            .I(\uart_drone.N_152 ));
    InMux I__9067 (
            .O(N__50838),
            .I(N__50835));
    LocalMux I__9066 (
            .O(N__50835),
            .I(N__50829));
    InMux I__9065 (
            .O(N__50834),
            .I(N__50824));
    InMux I__9064 (
            .O(N__50833),
            .I(N__50824));
    InMux I__9063 (
            .O(N__50832),
            .I(N__50820));
    Span4Mux_h I__9062 (
            .O(N__50829),
            .I(N__50815));
    LocalMux I__9061 (
            .O(N__50824),
            .I(N__50815));
    InMux I__9060 (
            .O(N__50823),
            .I(N__50809));
    LocalMux I__9059 (
            .O(N__50820),
            .I(N__50806));
    Span4Mux_h I__9058 (
            .O(N__50815),
            .I(N__50803));
    InMux I__9057 (
            .O(N__50814),
            .I(N__50796));
    InMux I__9056 (
            .O(N__50813),
            .I(N__50796));
    InMux I__9055 (
            .O(N__50812),
            .I(N__50796));
    LocalMux I__9054 (
            .O(N__50809),
            .I(\uart_drone.timer_CountZ1Z_3 ));
    Odrv4 I__9053 (
            .O(N__50806),
            .I(\uart_drone.timer_CountZ1Z_3 ));
    Odrv4 I__9052 (
            .O(N__50803),
            .I(\uart_drone.timer_CountZ1Z_3 ));
    LocalMux I__9051 (
            .O(N__50796),
            .I(\uart_drone.timer_CountZ1Z_3 ));
    InMux I__9050 (
            .O(N__50787),
            .I(N__50779));
    InMux I__9049 (
            .O(N__50786),
            .I(N__50774));
    InMux I__9048 (
            .O(N__50785),
            .I(N__50774));
    InMux I__9047 (
            .O(N__50784),
            .I(N__50771));
    InMux I__9046 (
            .O(N__50783),
            .I(N__50764));
    InMux I__9045 (
            .O(N__50782),
            .I(N__50764));
    LocalMux I__9044 (
            .O(N__50779),
            .I(N__50759));
    LocalMux I__9043 (
            .O(N__50774),
            .I(N__50759));
    LocalMux I__9042 (
            .O(N__50771),
            .I(N__50755));
    InMux I__9041 (
            .O(N__50770),
            .I(N__50750));
    InMux I__9040 (
            .O(N__50769),
            .I(N__50750));
    LocalMux I__9039 (
            .O(N__50764),
            .I(N__50747));
    Span4Mux_h I__9038 (
            .O(N__50759),
            .I(N__50744));
    InMux I__9037 (
            .O(N__50758),
            .I(N__50741));
    Span4Mux_v I__9036 (
            .O(N__50755),
            .I(N__50736));
    LocalMux I__9035 (
            .O(N__50750),
            .I(N__50736));
    Span4Mux_h I__9034 (
            .O(N__50747),
            .I(N__50731));
    Span4Mux_h I__9033 (
            .O(N__50744),
            .I(N__50731));
    LocalMux I__9032 (
            .O(N__50741),
            .I(\uart_drone.timer_CountZ0Z_4 ));
    Odrv4 I__9031 (
            .O(N__50736),
            .I(\uart_drone.timer_CountZ0Z_4 ));
    Odrv4 I__9030 (
            .O(N__50731),
            .I(\uart_drone.timer_CountZ0Z_4 ));
    CascadeMux I__9029 (
            .O(N__50724),
            .I(N__50721));
    InMux I__9028 (
            .O(N__50721),
            .I(N__50718));
    LocalMux I__9027 (
            .O(N__50718),
            .I(N__50714));
    InMux I__9026 (
            .O(N__50717),
            .I(N__50711));
    Span4Mux_h I__9025 (
            .O(N__50714),
            .I(N__50706));
    LocalMux I__9024 (
            .O(N__50711),
            .I(N__50706));
    Odrv4 I__9023 (
            .O(N__50706),
            .I(\uart_drone.N_144_1 ));
    InMux I__9022 (
            .O(N__50703),
            .I(N__50699));
    InMux I__9021 (
            .O(N__50702),
            .I(N__50696));
    LocalMux I__9020 (
            .O(N__50699),
            .I(N__50693));
    LocalMux I__9019 (
            .O(N__50696),
            .I(N__50690));
    Span12Mux_h I__9018 (
            .O(N__50693),
            .I(N__50687));
    Span12Mux_s2_h I__9017 (
            .O(N__50690),
            .I(N__50684));
    Odrv12 I__9016 (
            .O(N__50687),
            .I(xy_kp_5));
    Odrv12 I__9015 (
            .O(N__50684),
            .I(xy_kp_5));
    InMux I__9014 (
            .O(N__50679),
            .I(N__50676));
    LocalMux I__9013 (
            .O(N__50676),
            .I(N__50672));
    InMux I__9012 (
            .O(N__50675),
            .I(N__50669));
    Span12Mux_v I__9011 (
            .O(N__50672),
            .I(N__50666));
    LocalMux I__9010 (
            .O(N__50669),
            .I(N__50663));
    Span12Mux_h I__9009 (
            .O(N__50666),
            .I(N__50660));
    Span12Mux_s3_h I__9008 (
            .O(N__50663),
            .I(N__50657));
    Odrv12 I__9007 (
            .O(N__50660),
            .I(xy_kp_6));
    Odrv12 I__9006 (
            .O(N__50657),
            .I(xy_kp_6));
    IoInMux I__9005 (
            .O(N__50652),
            .I(N__50649));
    LocalMux I__9004 (
            .O(N__50649),
            .I(N__50646));
    Span12Mux_s1_v I__9003 (
            .O(N__50646),
            .I(N__50643));
    Odrv12 I__9002 (
            .O(N__50643),
            .I(\pid_side.state_RNIL5IFZ0Z_0 ));
    InMux I__9001 (
            .O(N__50640),
            .I(N__50637));
    LocalMux I__9000 (
            .O(N__50637),
            .I(N__50634));
    Span4Mux_h I__8999 (
            .O(N__50634),
            .I(N__50631));
    Odrv4 I__8998 (
            .O(N__50631),
            .I(\uart_drone.data_Auxce_0_0_4 ));
    InMux I__8997 (
            .O(N__50628),
            .I(N__50625));
    LocalMux I__8996 (
            .O(N__50625),
            .I(N__50622));
    Span4Mux_h I__8995 (
            .O(N__50622),
            .I(N__50619));
    Odrv4 I__8994 (
            .O(N__50619),
            .I(\uart_drone.data_Auxce_0_5 ));
    InMux I__8993 (
            .O(N__50616),
            .I(N__50613));
    LocalMux I__8992 (
            .O(N__50613),
            .I(N__50610));
    Span4Mux_h I__8991 (
            .O(N__50610),
            .I(N__50607));
    Odrv4 I__8990 (
            .O(N__50607),
            .I(\uart_drone.data_Auxce_0_6 ));
    InMux I__8989 (
            .O(N__50604),
            .I(N__50601));
    LocalMux I__8988 (
            .O(N__50601),
            .I(\ppm_encoder_1.un1_aileron_cry_2_THRU_CO ));
    InMux I__8987 (
            .O(N__50598),
            .I(N__50595));
    LocalMux I__8986 (
            .O(N__50595),
            .I(\ppm_encoder_1.un1_aileron_cry_11_THRU_CO ));
    InMux I__8985 (
            .O(N__50592),
            .I(N__50589));
    LocalMux I__8984 (
            .O(N__50589),
            .I(N__50586));
    Span4Mux_h I__8983 (
            .O(N__50586),
            .I(N__50583));
    Odrv4 I__8982 (
            .O(N__50583),
            .I(\ppm_encoder_1.un1_elevator_cry_5_THRU_CO ));
    InMux I__8981 (
            .O(N__50580),
            .I(N__50577));
    LocalMux I__8980 (
            .O(N__50577),
            .I(N__50574));
    Span4Mux_h I__8979 (
            .O(N__50574),
            .I(N__50570));
    InMux I__8978 (
            .O(N__50573),
            .I(N__50567));
    Span4Mux_v I__8977 (
            .O(N__50570),
            .I(N__50564));
    LocalMux I__8976 (
            .O(N__50567),
            .I(N__50561));
    Odrv4 I__8975 (
            .O(N__50564),
            .I(front_order_6));
    Odrv4 I__8974 (
            .O(N__50561),
            .I(front_order_6));
    CascadeMux I__8973 (
            .O(N__50556),
            .I(N__50552));
    InMux I__8972 (
            .O(N__50555),
            .I(N__50549));
    InMux I__8971 (
            .O(N__50552),
            .I(N__50546));
    LocalMux I__8970 (
            .O(N__50549),
            .I(N__50543));
    LocalMux I__8969 (
            .O(N__50546),
            .I(\ppm_encoder_1.elevatorZ0Z_6 ));
    Odrv12 I__8968 (
            .O(N__50543),
            .I(\ppm_encoder_1.elevatorZ0Z_6 ));
    InMux I__8967 (
            .O(N__50538),
            .I(N__50535));
    LocalMux I__8966 (
            .O(N__50535),
            .I(\ppm_encoder_1.un1_aileron_cry_5_THRU_CO ));
    InMux I__8965 (
            .O(N__50532),
            .I(N__50529));
    LocalMux I__8964 (
            .O(N__50529),
            .I(\ppm_encoder_1.un1_aileron_cry_6_THRU_CO ));
    InMux I__8963 (
            .O(N__50526),
            .I(N__50523));
    LocalMux I__8962 (
            .O(N__50523),
            .I(N__50518));
    InMux I__8961 (
            .O(N__50522),
            .I(N__50515));
    InMux I__8960 (
            .O(N__50521),
            .I(N__50512));
    Odrv4 I__8959 (
            .O(N__50518),
            .I(\uart_drone.un1_state_4_0 ));
    LocalMux I__8958 (
            .O(N__50515),
            .I(\uart_drone.un1_state_4_0 ));
    LocalMux I__8957 (
            .O(N__50512),
            .I(\uart_drone.un1_state_4_0 ));
    CascadeMux I__8956 (
            .O(N__50505),
            .I(\ppm_encoder_1.pulses2count_9_0_3_1_11_cascade_ ));
    InMux I__8955 (
            .O(N__50502),
            .I(N__50499));
    LocalMux I__8954 (
            .O(N__50499),
            .I(N__50495));
    InMux I__8953 (
            .O(N__50498),
            .I(N__50492));
    Span4Mux_h I__8952 (
            .O(N__50495),
            .I(N__50489));
    LocalMux I__8951 (
            .O(N__50492),
            .I(\ppm_encoder_1.elevatorZ0Z_13 ));
    Odrv4 I__8950 (
            .O(N__50489),
            .I(\ppm_encoder_1.elevatorZ0Z_13 ));
    InMux I__8949 (
            .O(N__50484),
            .I(N__50480));
    CascadeMux I__8948 (
            .O(N__50483),
            .I(N__50477));
    LocalMux I__8947 (
            .O(N__50480),
            .I(N__50474));
    InMux I__8946 (
            .O(N__50477),
            .I(N__50470));
    Span4Mux_v I__8945 (
            .O(N__50474),
            .I(N__50467));
    InMux I__8944 (
            .O(N__50473),
            .I(N__50464));
    LocalMux I__8943 (
            .O(N__50470),
            .I(\ppm_encoder_1.rudderZ0Z_12 ));
    Odrv4 I__8942 (
            .O(N__50467),
            .I(\ppm_encoder_1.rudderZ0Z_12 ));
    LocalMux I__8941 (
            .O(N__50464),
            .I(\ppm_encoder_1.rudderZ0Z_12 ));
    InMux I__8940 (
            .O(N__50457),
            .I(N__50454));
    LocalMux I__8939 (
            .O(N__50454),
            .I(\ppm_encoder_1.pulses2count_9_0_3_1_12 ));
    CascadeMux I__8938 (
            .O(N__50451),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_12_cascade_ ));
    InMux I__8937 (
            .O(N__50448),
            .I(N__50445));
    LocalMux I__8936 (
            .O(N__50445),
            .I(N__50440));
    InMux I__8935 (
            .O(N__50444),
            .I(N__50437));
    InMux I__8934 (
            .O(N__50443),
            .I(N__50433));
    Span4Mux_v I__8933 (
            .O(N__50440),
            .I(N__50428));
    LocalMux I__8932 (
            .O(N__50437),
            .I(N__50428));
    CascadeMux I__8931 (
            .O(N__50436),
            .I(N__50425));
    LocalMux I__8930 (
            .O(N__50433),
            .I(N__50422));
    Span4Mux_v I__8929 (
            .O(N__50428),
            .I(N__50419));
    InMux I__8928 (
            .O(N__50425),
            .I(N__50416));
    Span4Mux_v I__8927 (
            .O(N__50422),
            .I(N__50413));
    Span4Mux_s0_v I__8926 (
            .O(N__50419),
            .I(N__50408));
    LocalMux I__8925 (
            .O(N__50416),
            .I(N__50408));
    Odrv4 I__8924 (
            .O(N__50413),
            .I(\ppm_encoder_1.init_pulsesZ0Z_12 ));
    Odrv4 I__8923 (
            .O(N__50408),
            .I(\ppm_encoder_1.init_pulsesZ0Z_12 ));
    InMux I__8922 (
            .O(N__50403),
            .I(N__50400));
    LocalMux I__8921 (
            .O(N__50400),
            .I(N__50397));
    Odrv4 I__8920 (
            .O(N__50397),
            .I(\uart_drone.data_Auxce_0_1 ));
    InMux I__8919 (
            .O(N__50394),
            .I(N__50391));
    LocalMux I__8918 (
            .O(N__50391),
            .I(N__50388));
    Span4Mux_h I__8917 (
            .O(N__50388),
            .I(N__50385));
    Odrv4 I__8916 (
            .O(N__50385),
            .I(\uart_drone.data_Auxce_0_0_2 ));
    InMux I__8915 (
            .O(N__50382),
            .I(N__50379));
    LocalMux I__8914 (
            .O(N__50379),
            .I(\ppm_encoder_1.elevator_RNIOEGEZ0Z_10 ));
    InMux I__8913 (
            .O(N__50376),
            .I(N__50373));
    LocalMux I__8912 (
            .O(N__50373),
            .I(\ppm_encoder_1.un2_throttle_iv_0_2_10 ));
    CascadeMux I__8911 (
            .O(N__50370),
            .I(N__50367));
    InMux I__8910 (
            .O(N__50367),
            .I(N__50364));
    LocalMux I__8909 (
            .O(N__50364),
            .I(N__50361));
    Span4Mux_h I__8908 (
            .O(N__50361),
            .I(N__50357));
    InMux I__8907 (
            .O(N__50360),
            .I(N__50354));
    Odrv4 I__8906 (
            .O(N__50357),
            .I(\ppm_encoder_1.N_255_i_i ));
    LocalMux I__8905 (
            .O(N__50354),
            .I(\ppm_encoder_1.N_255_i_i ));
    InMux I__8904 (
            .O(N__50349),
            .I(N__50346));
    LocalMux I__8903 (
            .O(N__50346),
            .I(N__50343));
    Span4Mux_v I__8902 (
            .O(N__50343),
            .I(N__50340));
    Odrv4 I__8901 (
            .O(N__50340),
            .I(\ppm_encoder_1.un1_aileron_cry_0_THRU_CO ));
    InMux I__8900 (
            .O(N__50337),
            .I(N__50334));
    LocalMux I__8899 (
            .O(N__50334),
            .I(N__50331));
    Span4Mux_h I__8898 (
            .O(N__50331),
            .I(N__50328));
    Odrv4 I__8897 (
            .O(N__50328),
            .I(\ppm_encoder_1.un1_throttle_cry_0_THRU_CO ));
    CascadeMux I__8896 (
            .O(N__50325),
            .I(N__50322));
    InMux I__8895 (
            .O(N__50322),
            .I(N__50319));
    LocalMux I__8894 (
            .O(N__50319),
            .I(N__50316));
    Span4Mux_v I__8893 (
            .O(N__50316),
            .I(N__50312));
    InMux I__8892 (
            .O(N__50315),
            .I(N__50309));
    Span4Mux_h I__8891 (
            .O(N__50312),
            .I(N__50304));
    LocalMux I__8890 (
            .O(N__50309),
            .I(N__50304));
    Span4Mux_v I__8889 (
            .O(N__50304),
            .I(N__50301));
    Odrv4 I__8888 (
            .O(N__50301),
            .I(throttle_order_1));
    InMux I__8887 (
            .O(N__50298),
            .I(N__50295));
    LocalMux I__8886 (
            .O(N__50295),
            .I(N__50292));
    Span4Mux_h I__8885 (
            .O(N__50292),
            .I(N__50289));
    Span4Mux_v I__8884 (
            .O(N__50289),
            .I(N__50286));
    Odrv4 I__8883 (
            .O(N__50286),
            .I(\ppm_encoder_1.un1_elevator_cry_6_THRU_CO ));
    InMux I__8882 (
            .O(N__50283),
            .I(N__50280));
    LocalMux I__8881 (
            .O(N__50280),
            .I(N__50277));
    Span4Mux_h I__8880 (
            .O(N__50277),
            .I(N__50273));
    InMux I__8879 (
            .O(N__50276),
            .I(N__50270));
    Span4Mux_v I__8878 (
            .O(N__50273),
            .I(N__50265));
    LocalMux I__8877 (
            .O(N__50270),
            .I(N__50265));
    Odrv4 I__8876 (
            .O(N__50265),
            .I(front_order_7));
    InMux I__8875 (
            .O(N__50262),
            .I(N__50256));
    InMux I__8874 (
            .O(N__50261),
            .I(N__50256));
    LocalMux I__8873 (
            .O(N__50256),
            .I(\ppm_encoder_1.elevatorZ0Z_7 ));
    InMux I__8872 (
            .O(N__50253),
            .I(N__50250));
    LocalMux I__8871 (
            .O(N__50250),
            .I(\ppm_encoder_1.un2_throttle_iv_0_0_6 ));
    CascadeMux I__8870 (
            .O(N__50247),
            .I(\ppm_encoder_1.un2_throttle_iv_0_1_6_cascade_ ));
    CascadeMux I__8869 (
            .O(N__50244),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_6_cascade_ ));
    CascadeMux I__8868 (
            .O(N__50241),
            .I(N__50237));
    InMux I__8867 (
            .O(N__50240),
            .I(N__50234));
    InMux I__8866 (
            .O(N__50237),
            .I(N__50231));
    LocalMux I__8865 (
            .O(N__50234),
            .I(N__50226));
    LocalMux I__8864 (
            .O(N__50231),
            .I(N__50223));
    InMux I__8863 (
            .O(N__50230),
            .I(N__50220));
    InMux I__8862 (
            .O(N__50229),
            .I(N__50217));
    Odrv4 I__8861 (
            .O(N__50226),
            .I(\ppm_encoder_1.N_262_i_i ));
    Odrv4 I__8860 (
            .O(N__50223),
            .I(\ppm_encoder_1.N_262_i_i ));
    LocalMux I__8859 (
            .O(N__50220),
            .I(\ppm_encoder_1.N_262_i_i ));
    LocalMux I__8858 (
            .O(N__50217),
            .I(\ppm_encoder_1.N_262_i_i ));
    InMux I__8857 (
            .O(N__50208),
            .I(N__50205));
    LocalMux I__8856 (
            .O(N__50205),
            .I(N__50202));
    Odrv4 I__8855 (
            .O(N__50202),
            .I(\ppm_encoder_1.init_pulses_RNIPOJU5Z0Z_6 ));
    InMux I__8854 (
            .O(N__50199),
            .I(N__50196));
    LocalMux I__8853 (
            .O(N__50196),
            .I(\ppm_encoder_1.elevator_RNIB86OZ0Z_4 ));
    InMux I__8852 (
            .O(N__50193),
            .I(N__50190));
    LocalMux I__8851 (
            .O(N__50190),
            .I(N__50187));
    Odrv12 I__8850 (
            .O(N__50187),
            .I(\ppm_encoder_1.un2_throttle_iv_0_2_4 ));
    InMux I__8849 (
            .O(N__50184),
            .I(N__50181));
    LocalMux I__8848 (
            .O(N__50181),
            .I(N__50178));
    Span4Mux_v I__8847 (
            .O(N__50178),
            .I(N__50174));
    CascadeMux I__8846 (
            .O(N__50177),
            .I(N__50171));
    Span4Mux_v I__8845 (
            .O(N__50174),
            .I(N__50168));
    InMux I__8844 (
            .O(N__50171),
            .I(N__50165));
    Odrv4 I__8843 (
            .O(N__50168),
            .I(scaler_4_data_4));
    LocalMux I__8842 (
            .O(N__50165),
            .I(scaler_4_data_4));
    CEMux I__8841 (
            .O(N__50160),
            .I(N__50155));
    CEMux I__8840 (
            .O(N__50159),
            .I(N__50150));
    CEMux I__8839 (
            .O(N__50158),
            .I(N__50147));
    LocalMux I__8838 (
            .O(N__50155),
            .I(N__50143));
    CEMux I__8837 (
            .O(N__50154),
            .I(N__50140));
    CEMux I__8836 (
            .O(N__50153),
            .I(N__50137));
    LocalMux I__8835 (
            .O(N__50150),
            .I(N__50134));
    LocalMux I__8834 (
            .O(N__50147),
            .I(N__50131));
    CEMux I__8833 (
            .O(N__50146),
            .I(N__50128));
    Span4Mux_s3_v I__8832 (
            .O(N__50143),
            .I(N__50125));
    LocalMux I__8831 (
            .O(N__50140),
            .I(N__50122));
    LocalMux I__8830 (
            .O(N__50137),
            .I(N__50119));
    Span4Mux_h I__8829 (
            .O(N__50134),
            .I(N__50116));
    Span4Mux_v I__8828 (
            .O(N__50131),
            .I(N__50113));
    LocalMux I__8827 (
            .O(N__50128),
            .I(N__50108));
    Span4Mux_h I__8826 (
            .O(N__50125),
            .I(N__50108));
    Span4Mux_h I__8825 (
            .O(N__50122),
            .I(N__50103));
    Span4Mux_v I__8824 (
            .O(N__50119),
            .I(N__50103));
    Span4Mux_h I__8823 (
            .O(N__50116),
            .I(N__50100));
    Span4Mux_h I__8822 (
            .O(N__50113),
            .I(N__50095));
    Span4Mux_h I__8821 (
            .O(N__50108),
            .I(N__50095));
    Span4Mux_h I__8820 (
            .O(N__50103),
            .I(N__50092));
    Odrv4 I__8819 (
            .O(N__50100),
            .I(\ppm_encoder_1.pid_altitude_dv_0 ));
    Odrv4 I__8818 (
            .O(N__50095),
            .I(\ppm_encoder_1.pid_altitude_dv_0 ));
    Odrv4 I__8817 (
            .O(N__50092),
            .I(\ppm_encoder_1.pid_altitude_dv_0 ));
    CascadeMux I__8816 (
            .O(N__50085),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_10_cascade_ ));
    InMux I__8815 (
            .O(N__50082),
            .I(N__50079));
    LocalMux I__8814 (
            .O(N__50079),
            .I(N__50076));
    Span4Mux_v I__8813 (
            .O(N__50076),
            .I(N__50073));
    Odrv4 I__8812 (
            .O(N__50073),
            .I(\ppm_encoder_1.init_pulses_RNIUCPF5Z0Z_10 ));
    InMux I__8811 (
            .O(N__50070),
            .I(N__50067));
    LocalMux I__8810 (
            .O(N__50067),
            .I(\ppm_encoder_1.elevator_RNIGD6OZ0Z_9 ));
    InMux I__8809 (
            .O(N__50064),
            .I(N__50061));
    LocalMux I__8808 (
            .O(N__50061),
            .I(\ppm_encoder_1.un2_throttle_iv_0_2_9 ));
    CascadeMux I__8807 (
            .O(N__50058),
            .I(\ppm_encoder_1.N_56_cascade_ ));
    CascadeMux I__8806 (
            .O(N__50055),
            .I(N__50052));
    InMux I__8805 (
            .O(N__50052),
            .I(N__50049));
    LocalMux I__8804 (
            .O(N__50049),
            .I(\ppm_encoder_1.init_pulses_RNIV9203Z0Z_6 ));
    InMux I__8803 (
            .O(N__50046),
            .I(N__50043));
    LocalMux I__8802 (
            .O(N__50043),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_12 ));
    CascadeMux I__8801 (
            .O(N__50040),
            .I(N__50037));
    InMux I__8800 (
            .O(N__50037),
            .I(N__50034));
    LocalMux I__8799 (
            .O(N__50034),
            .I(N__50031));
    Span4Mux_h I__8798 (
            .O(N__50031),
            .I(N__50028));
    Odrv4 I__8797 (
            .O(N__50028),
            .I(\ppm_encoder_1.N_254_i_i ));
    CascadeMux I__8796 (
            .O(N__50025),
            .I(\ppm_encoder_1.N_254_i_i_cascade_ ));
    InMux I__8795 (
            .O(N__50022),
            .I(N__50019));
    LocalMux I__8794 (
            .O(N__50019),
            .I(N__50016));
    Span4Mux_h I__8793 (
            .O(N__50016),
            .I(N__50013));
    Odrv4 I__8792 (
            .O(N__50013),
            .I(\ppm_encoder_1.init_pulses_RNI82G01Z0Z_15 ));
    CascadeMux I__8791 (
            .O(N__50010),
            .I(\ppm_encoder_1.N_268_i_i_cascade_ ));
    CascadeMux I__8790 (
            .O(N__50007),
            .I(N__50004));
    InMux I__8789 (
            .O(N__50004),
            .I(N__50001));
    LocalMux I__8788 (
            .O(N__50001),
            .I(\ppm_encoder_1.init_pulses_RNITIRP2Z0Z_13 ));
    InMux I__8787 (
            .O(N__49998),
            .I(N__49995));
    LocalMux I__8786 (
            .O(N__49995),
            .I(\pid_front.un10lto27_10 ));
    InMux I__8785 (
            .O(N__49992),
            .I(N__49988));
    InMux I__8784 (
            .O(N__49991),
            .I(N__49985));
    LocalMux I__8783 (
            .O(N__49988),
            .I(\pid_front.error_i_acumm_preregZ0Z_19 ));
    LocalMux I__8782 (
            .O(N__49985),
            .I(\pid_front.error_i_acumm_preregZ0Z_19 ));
    InMux I__8781 (
            .O(N__49980),
            .I(N__49976));
    InMux I__8780 (
            .O(N__49979),
            .I(N__49973));
    LocalMux I__8779 (
            .O(N__49976),
            .I(\pid_front.error_i_acumm_preregZ0Z_18 ));
    LocalMux I__8778 (
            .O(N__49973),
            .I(\pid_front.error_i_acumm_preregZ0Z_18 ));
    InMux I__8777 (
            .O(N__49968),
            .I(N__49962));
    InMux I__8776 (
            .O(N__49967),
            .I(N__49962));
    LocalMux I__8775 (
            .O(N__49962),
            .I(\pid_front.error_i_acumm_preregZ0Z_14 ));
    CascadeMux I__8774 (
            .O(N__49959),
            .I(N__49956));
    InMux I__8773 (
            .O(N__49956),
            .I(N__49950));
    InMux I__8772 (
            .O(N__49955),
            .I(N__49950));
    LocalMux I__8771 (
            .O(N__49950),
            .I(\pid_front.error_i_acumm_preregZ0Z_15 ));
    InMux I__8770 (
            .O(N__49947),
            .I(N__49944));
    LocalMux I__8769 (
            .O(N__49944),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_1 ));
    CascadeMux I__8768 (
            .O(N__49941),
            .I(N__49938));
    InMux I__8767 (
            .O(N__49938),
            .I(N__49935));
    LocalMux I__8766 (
            .O(N__49935),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_3 ));
    InMux I__8765 (
            .O(N__49932),
            .I(N__49929));
    LocalMux I__8764 (
            .O(N__49929),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_10 ));
    InMux I__8763 (
            .O(N__49926),
            .I(N__49923));
    LocalMux I__8762 (
            .O(N__49923),
            .I(N__49920));
    Span12Mux_s11_v I__8761 (
            .O(N__49920),
            .I(N__49917));
    Odrv12 I__8760 (
            .O(N__49917),
            .I(\ppm_encoder_1.elevatorZ0Z_14 ));
    CascadeMux I__8759 (
            .O(N__49914),
            .I(N__49911));
    InMux I__8758 (
            .O(N__49911),
            .I(N__49908));
    LocalMux I__8757 (
            .O(N__49908),
            .I(N__49905));
    Span4Mux_s2_v I__8756 (
            .O(N__49905),
            .I(N__49902));
    Span4Mux_v I__8755 (
            .O(N__49902),
            .I(N__49899));
    Odrv4 I__8754 (
            .O(N__49899),
            .I(\ppm_encoder_1.rudderZ0Z_14 ));
    CascadeMux I__8753 (
            .O(N__49896),
            .I(\pid_front.error_i_acumm_prereg_esr_RNIRU7IZ0Z_10_cascade_ ));
    InMux I__8752 (
            .O(N__49893),
            .I(N__49890));
    LocalMux I__8751 (
            .O(N__49890),
            .I(\pid_front.un10lt11_0 ));
    InMux I__8750 (
            .O(N__49887),
            .I(N__49884));
    LocalMux I__8749 (
            .O(N__49884),
            .I(N__49881));
    Span12Mux_h I__8748 (
            .O(N__49881),
            .I(N__49878));
    Span12Mux_h I__8747 (
            .O(N__49878),
            .I(N__49875));
    Odrv12 I__8746 (
            .O(N__49875),
            .I(\pid_front.O_2 ));
    CascadeMux I__8745 (
            .O(N__49872),
            .I(\pid_front.un10lto27_9_cascade_ ));
    InMux I__8744 (
            .O(N__49869),
            .I(N__49866));
    LocalMux I__8743 (
            .O(N__49866),
            .I(\pid_front.error_i_acumm_prereg_esr_RNI18694_0Z0Z_14 ));
    CascadeMux I__8742 (
            .O(N__49863),
            .I(N__49860));
    InMux I__8741 (
            .O(N__49860),
            .I(N__49857));
    LocalMux I__8740 (
            .O(N__49857),
            .I(\pid_front.un10lt9_1 ));
    CascadeMux I__8739 (
            .O(N__49854),
            .I(\pid_front.error_i_acumm16lt9_0_cascade_ ));
    InMux I__8738 (
            .O(N__49851),
            .I(N__49848));
    LocalMux I__8737 (
            .O(N__49848),
            .I(\pid_front.error_i_acumm_prereg_esr_RNISDO3Z0Z_7 ));
    InMux I__8736 (
            .O(N__49845),
            .I(N__49842));
    LocalMux I__8735 (
            .O(N__49842),
            .I(N__49839));
    Sp12to4 I__8734 (
            .O(N__49839),
            .I(N__49836));
    Span12Mux_v I__8733 (
            .O(N__49836),
            .I(N__49833));
    Odrv12 I__8732 (
            .O(N__49833),
            .I(\pid_front.O_0_4 ));
    CascadeMux I__8731 (
            .O(N__49830),
            .I(\pid_front.un1_pid_prereg_9_0_cascade_ ));
    InMux I__8730 (
            .O(N__49827),
            .I(N__49824));
    LocalMux I__8729 (
            .O(N__49824),
            .I(N__49821));
    Span4Mux_h I__8728 (
            .O(N__49821),
            .I(N__49818));
    Span4Mux_v I__8727 (
            .O(N__49818),
            .I(N__49815));
    Odrv4 I__8726 (
            .O(N__49815),
            .I(\pid_front.error_d_reg_prev_esr_RNIMRLTZ0Z_0 ));
    InMux I__8725 (
            .O(N__49812),
            .I(N__49809));
    LocalMux I__8724 (
            .O(N__49809),
            .I(N__49806));
    Span4Mux_v I__8723 (
            .O(N__49806),
            .I(N__49803));
    Span4Mux_h I__8722 (
            .O(N__49803),
            .I(N__49800));
    Span4Mux_h I__8721 (
            .O(N__49800),
            .I(N__49797));
    Span4Mux_h I__8720 (
            .O(N__49797),
            .I(N__49794));
    Odrv4 I__8719 (
            .O(N__49794),
            .I(\pid_front.O_3 ));
    InMux I__8718 (
            .O(N__49791),
            .I(N__49788));
    LocalMux I__8717 (
            .O(N__49788),
            .I(N__49785));
    Span12Mux_s11_h I__8716 (
            .O(N__49785),
            .I(N__49782));
    Odrv12 I__8715 (
            .O(N__49782),
            .I(\pid_front.error_d_reg_prev_esr_RNIAHDKZ0Z_0 ));
    InMux I__8714 (
            .O(N__49779),
            .I(N__49771));
    InMux I__8713 (
            .O(N__49778),
            .I(N__49771));
    InMux I__8712 (
            .O(N__49777),
            .I(N__49766));
    InMux I__8711 (
            .O(N__49776),
            .I(N__49766));
    LocalMux I__8710 (
            .O(N__49771),
            .I(N__49763));
    LocalMux I__8709 (
            .O(N__49766),
            .I(N__49760));
    Span4Mux_v I__8708 (
            .O(N__49763),
            .I(N__49757));
    Odrv12 I__8707 (
            .O(N__49760),
            .I(\pid_front.error_d_regZ0Z_6 ));
    Odrv4 I__8706 (
            .O(N__49757),
            .I(\pid_front.error_d_regZ0Z_6 ));
    InMux I__8705 (
            .O(N__49752),
            .I(N__49749));
    LocalMux I__8704 (
            .O(N__49749),
            .I(N__49746));
    Span4Mux_v I__8703 (
            .O(N__49746),
            .I(N__49743));
    Span4Mux_h I__8702 (
            .O(N__49743),
            .I(N__49740));
    Span4Mux_h I__8701 (
            .O(N__49740),
            .I(N__49737));
    Span4Mux_h I__8700 (
            .O(N__49737),
            .I(N__49734));
    Odrv4 I__8699 (
            .O(N__49734),
            .I(\pid_front.O_9 ));
    InMux I__8698 (
            .O(N__49731),
            .I(N__49725));
    InMux I__8697 (
            .O(N__49730),
            .I(N__49718));
    InMux I__8696 (
            .O(N__49729),
            .I(N__49718));
    InMux I__8695 (
            .O(N__49728),
            .I(N__49718));
    LocalMux I__8694 (
            .O(N__49725),
            .I(N__49713));
    LocalMux I__8693 (
            .O(N__49718),
            .I(N__49713));
    Odrv12 I__8692 (
            .O(N__49713),
            .I(\pid_front.error_d_regZ0Z_7 ));
    InMux I__8691 (
            .O(N__49710),
            .I(N__49707));
    LocalMux I__8690 (
            .O(N__49707),
            .I(N__49704));
    Span4Mux_h I__8689 (
            .O(N__49704),
            .I(N__49701));
    Span4Mux_h I__8688 (
            .O(N__49701),
            .I(N__49698));
    Span4Mux_h I__8687 (
            .O(N__49698),
            .I(N__49695));
    Span4Mux_h I__8686 (
            .O(N__49695),
            .I(N__49692));
    Odrv4 I__8685 (
            .O(N__49692),
            .I(\pid_front.O_10 ));
    InMux I__8684 (
            .O(N__49689),
            .I(N__49683));
    InMux I__8683 (
            .O(N__49688),
            .I(N__49678));
    InMux I__8682 (
            .O(N__49687),
            .I(N__49678));
    InMux I__8681 (
            .O(N__49686),
            .I(N__49675));
    LocalMux I__8680 (
            .O(N__49683),
            .I(N__49670));
    LocalMux I__8679 (
            .O(N__49678),
            .I(N__49670));
    LocalMux I__8678 (
            .O(N__49675),
            .I(N__49667));
    Span4Mux_v I__8677 (
            .O(N__49670),
            .I(N__49664));
    Sp12to4 I__8676 (
            .O(N__49667),
            .I(N__49661));
    Odrv4 I__8675 (
            .O(N__49664),
            .I(\pid_front.error_d_regZ0Z_8 ));
    Odrv12 I__8674 (
            .O(N__49661),
            .I(\pid_front.error_d_regZ0Z_8 ));
    InMux I__8673 (
            .O(N__49656),
            .I(N__49653));
    LocalMux I__8672 (
            .O(N__49653),
            .I(N__49649));
    InMux I__8671 (
            .O(N__49652),
            .I(N__49646));
    Sp12to4 I__8670 (
            .O(N__49649),
            .I(N__49643));
    LocalMux I__8669 (
            .O(N__49646),
            .I(N__49640));
    Span12Mux_s6_v I__8668 (
            .O(N__49643),
            .I(N__49635));
    Span12Mux_v I__8667 (
            .O(N__49640),
            .I(N__49635));
    Span12Mux_h I__8666 (
            .O(N__49635),
            .I(N__49632));
    Odrv12 I__8665 (
            .O(N__49632),
            .I(\pid_front.O_14 ));
    InMux I__8664 (
            .O(N__49629),
            .I(N__49616));
    InMux I__8663 (
            .O(N__49628),
            .I(N__49616));
    InMux I__8662 (
            .O(N__49627),
            .I(N__49611));
    InMux I__8661 (
            .O(N__49626),
            .I(N__49611));
    InMux I__8660 (
            .O(N__49625),
            .I(N__49608));
    InMux I__8659 (
            .O(N__49624),
            .I(N__49604));
    InMux I__8658 (
            .O(N__49623),
            .I(N__49597));
    InMux I__8657 (
            .O(N__49622),
            .I(N__49597));
    InMux I__8656 (
            .O(N__49621),
            .I(N__49597));
    LocalMux I__8655 (
            .O(N__49616),
            .I(N__49592));
    LocalMux I__8654 (
            .O(N__49611),
            .I(N__49592));
    LocalMux I__8653 (
            .O(N__49608),
            .I(N__49589));
    InMux I__8652 (
            .O(N__49607),
            .I(N__49586));
    LocalMux I__8651 (
            .O(N__49604),
            .I(N__49581));
    LocalMux I__8650 (
            .O(N__49597),
            .I(N__49581));
    Span4Mux_v I__8649 (
            .O(N__49592),
            .I(N__49576));
    Span4Mux_h I__8648 (
            .O(N__49589),
            .I(N__49576));
    LocalMux I__8647 (
            .O(N__49586),
            .I(\pid_front.error_d_regZ0Z_12 ));
    Odrv4 I__8646 (
            .O(N__49581),
            .I(\pid_front.error_d_regZ0Z_12 ));
    Odrv4 I__8645 (
            .O(N__49576),
            .I(\pid_front.error_d_regZ0Z_12 ));
    InMux I__8644 (
            .O(N__49569),
            .I(N__49566));
    LocalMux I__8643 (
            .O(N__49566),
            .I(N__49563));
    Span4Mux_v I__8642 (
            .O(N__49563),
            .I(N__49560));
    Sp12to4 I__8641 (
            .O(N__49560),
            .I(N__49557));
    Span12Mux_h I__8640 (
            .O(N__49557),
            .I(N__49554));
    Odrv12 I__8639 (
            .O(N__49554),
            .I(\pid_front.O_0_3 ));
    CascadeMux I__8638 (
            .O(N__49551),
            .I(N__49548));
    InMux I__8637 (
            .O(N__49548),
            .I(N__49544));
    InMux I__8636 (
            .O(N__49547),
            .I(N__49541));
    LocalMux I__8635 (
            .O(N__49544),
            .I(N__49536));
    LocalMux I__8634 (
            .O(N__49541),
            .I(N__49536));
    Span4Mux_h I__8633 (
            .O(N__49536),
            .I(N__49533));
    Span4Mux_v I__8632 (
            .O(N__49533),
            .I(N__49530));
    Odrv4 I__8631 (
            .O(N__49530),
            .I(\pid_front.error_p_regZ0Z_0 ));
    InMux I__8630 (
            .O(N__49527),
            .I(N__49524));
    LocalMux I__8629 (
            .O(N__49524),
            .I(N__49521));
    Span12Mux_v I__8628 (
            .O(N__49521),
            .I(N__49518));
    Odrv12 I__8627 (
            .O(N__49518),
            .I(\pid_front.O_0_13 ));
    InMux I__8626 (
            .O(N__49515),
            .I(N__49512));
    LocalMux I__8625 (
            .O(N__49512),
            .I(N__49508));
    CascadeMux I__8624 (
            .O(N__49511),
            .I(N__49504));
    Span4Mux_v I__8623 (
            .O(N__49508),
            .I(N__49501));
    InMux I__8622 (
            .O(N__49507),
            .I(N__49496));
    InMux I__8621 (
            .O(N__49504),
            .I(N__49496));
    Odrv4 I__8620 (
            .O(N__49501),
            .I(\pid_front.error_p_regZ0Z_10 ));
    LocalMux I__8619 (
            .O(N__49496),
            .I(\pid_front.error_p_regZ0Z_10 ));
    CascadeMux I__8618 (
            .O(N__49491),
            .I(\pid_front.un10lt9_1_cascade_ ));
    CascadeMux I__8617 (
            .O(N__49488),
            .I(\pid_front.un10lt9_cascade_ ));
    InMux I__8616 (
            .O(N__49485),
            .I(N__49482));
    LocalMux I__8615 (
            .O(N__49482),
            .I(N__49479));
    Span4Mux_v I__8614 (
            .O(N__49479),
            .I(N__49475));
    InMux I__8613 (
            .O(N__49478),
            .I(N__49471));
    Span4Mux_h I__8612 (
            .O(N__49475),
            .I(N__49468));
    InMux I__8611 (
            .O(N__49474),
            .I(N__49465));
    LocalMux I__8610 (
            .O(N__49471),
            .I(N__49461));
    Sp12to4 I__8609 (
            .O(N__49468),
            .I(N__49456));
    LocalMux I__8608 (
            .O(N__49465),
            .I(N__49456));
    InMux I__8607 (
            .O(N__49464),
            .I(N__49453));
    Span4Mux_h I__8606 (
            .O(N__49461),
            .I(N__49450));
    Odrv12 I__8605 (
            .O(N__49456),
            .I(\pid_alt.error_i_acumm_preregZ0Z_21 ));
    LocalMux I__8604 (
            .O(N__49453),
            .I(\pid_alt.error_i_acumm_preregZ0Z_21 ));
    Odrv4 I__8603 (
            .O(N__49450),
            .I(\pid_alt.error_i_acumm_preregZ0Z_21 ));
    InMux I__8602 (
            .O(N__49443),
            .I(N__49440));
    LocalMux I__8601 (
            .O(N__49440),
            .I(N__49435));
    InMux I__8600 (
            .O(N__49439),
            .I(N__49432));
    InMux I__8599 (
            .O(N__49438),
            .I(N__49429));
    Odrv12 I__8598 (
            .O(N__49435),
            .I(\pid_alt.error_i_acumm7lto13 ));
    LocalMux I__8597 (
            .O(N__49432),
            .I(\pid_alt.error_i_acumm7lto13 ));
    LocalMux I__8596 (
            .O(N__49429),
            .I(\pid_alt.error_i_acumm7lto13 ));
    InMux I__8595 (
            .O(N__49422),
            .I(N__49419));
    LocalMux I__8594 (
            .O(N__49419),
            .I(N__49416));
    Span4Mux_h I__8593 (
            .O(N__49416),
            .I(N__49412));
    InMux I__8592 (
            .O(N__49415),
            .I(N__49409));
    Span4Mux_h I__8591 (
            .O(N__49412),
            .I(N__49404));
    LocalMux I__8590 (
            .O(N__49409),
            .I(N__49404));
    Odrv4 I__8589 (
            .O(N__49404),
            .I(\pid_alt.N_545 ));
    InMux I__8588 (
            .O(N__49401),
            .I(N__49398));
    LocalMux I__8587 (
            .O(N__49398),
            .I(N__49395));
    Span4Mux_s3_h I__8586 (
            .O(N__49395),
            .I(N__49392));
    Span4Mux_h I__8585 (
            .O(N__49392),
            .I(N__49389));
    Span4Mux_h I__8584 (
            .O(N__49389),
            .I(N__49386));
    Odrv4 I__8583 (
            .O(N__49386),
            .I(\pid_alt.error_i_acummZ0Z_13 ));
    CEMux I__8582 (
            .O(N__49383),
            .I(N__49380));
    LocalMux I__8581 (
            .O(N__49380),
            .I(N__49377));
    Span4Mux_h I__8580 (
            .O(N__49377),
            .I(N__49373));
    CEMux I__8579 (
            .O(N__49376),
            .I(N__49370));
    Span4Mux_h I__8578 (
            .O(N__49373),
            .I(N__49367));
    LocalMux I__8577 (
            .O(N__49370),
            .I(N__49364));
    Odrv4 I__8576 (
            .O(N__49367),
            .I(\pid_alt.N_72_i_0 ));
    Odrv4 I__8575 (
            .O(N__49364),
            .I(\pid_alt.N_72_i_0 ));
    SRMux I__8574 (
            .O(N__49359),
            .I(N__49355));
    SRMux I__8573 (
            .O(N__49358),
            .I(N__49352));
    LocalMux I__8572 (
            .O(N__49355),
            .I(N__49348));
    LocalMux I__8571 (
            .O(N__49352),
            .I(N__49345));
    SRMux I__8570 (
            .O(N__49351),
            .I(N__49342));
    Span4Mux_h I__8569 (
            .O(N__49348),
            .I(N__49338));
    Span4Mux_h I__8568 (
            .O(N__49345),
            .I(N__49335));
    LocalMux I__8567 (
            .O(N__49342),
            .I(N__49332));
    SRMux I__8566 (
            .O(N__49341),
            .I(N__49329));
    Span4Mux_h I__8565 (
            .O(N__49338),
            .I(N__49325));
    Span4Mux_h I__8564 (
            .O(N__49335),
            .I(N__49322));
    Span4Mux_v I__8563 (
            .O(N__49332),
            .I(N__49319));
    LocalMux I__8562 (
            .O(N__49329),
            .I(N__49316));
    InMux I__8561 (
            .O(N__49328),
            .I(N__49313));
    Odrv4 I__8560 (
            .O(N__49325),
            .I(\pid_alt.un1_reset_1_0_i ));
    Odrv4 I__8559 (
            .O(N__49322),
            .I(\pid_alt.un1_reset_1_0_i ));
    Odrv4 I__8558 (
            .O(N__49319),
            .I(\pid_alt.un1_reset_1_0_i ));
    Odrv12 I__8557 (
            .O(N__49316),
            .I(\pid_alt.un1_reset_1_0_i ));
    LocalMux I__8556 (
            .O(N__49313),
            .I(\pid_alt.un1_reset_1_0_i ));
    CascadeMux I__8555 (
            .O(N__49302),
            .I(N__49299));
    InMux I__8554 (
            .O(N__49299),
            .I(N__49293));
    InMux I__8553 (
            .O(N__49298),
            .I(N__49293));
    LocalMux I__8552 (
            .O(N__49293),
            .I(N__49290));
    Odrv4 I__8551 (
            .O(N__49290),
            .I(\pid_front.error_d_reg_prevZ0Z_19 ));
    InMux I__8550 (
            .O(N__49287),
            .I(N__49281));
    InMux I__8549 (
            .O(N__49286),
            .I(N__49281));
    LocalMux I__8548 (
            .O(N__49281),
            .I(N__49278));
    Span4Mux_v I__8547 (
            .O(N__49278),
            .I(N__49275));
    Span4Mux_h I__8546 (
            .O(N__49275),
            .I(N__49272));
    Span4Mux_h I__8545 (
            .O(N__49272),
            .I(N__49269));
    Span4Mux_v I__8544 (
            .O(N__49269),
            .I(N__49266));
    Odrv4 I__8543 (
            .O(N__49266),
            .I(\pid_front.error_p_regZ0Z_19 ));
    InMux I__8542 (
            .O(N__49263),
            .I(N__49257));
    InMux I__8541 (
            .O(N__49262),
            .I(N__49257));
    LocalMux I__8540 (
            .O(N__49257),
            .I(N__49254));
    Span4Mux_v I__8539 (
            .O(N__49254),
            .I(N__49251));
    Odrv4 I__8538 (
            .O(N__49251),
            .I(\pid_front.error_p_reg_esr_RNI0GC61Z0Z_19 ));
    InMux I__8537 (
            .O(N__49248),
            .I(N__49240));
    InMux I__8536 (
            .O(N__49247),
            .I(N__49240));
    InMux I__8535 (
            .O(N__49246),
            .I(N__49237));
    InMux I__8534 (
            .O(N__49245),
            .I(N__49234));
    LocalMux I__8533 (
            .O(N__49240),
            .I(N__49231));
    LocalMux I__8532 (
            .O(N__49237),
            .I(\pid_front.un1_pid_prereg_135_0 ));
    LocalMux I__8531 (
            .O(N__49234),
            .I(\pid_front.un1_pid_prereg_135_0 ));
    Odrv4 I__8530 (
            .O(N__49231),
            .I(\pid_front.un1_pid_prereg_135_0 ));
    InMux I__8529 (
            .O(N__49224),
            .I(N__49220));
    InMux I__8528 (
            .O(N__49223),
            .I(N__49217));
    LocalMux I__8527 (
            .O(N__49220),
            .I(N__49212));
    LocalMux I__8526 (
            .O(N__49217),
            .I(N__49209));
    InMux I__8525 (
            .O(N__49216),
            .I(N__49204));
    InMux I__8524 (
            .O(N__49215),
            .I(N__49204));
    Span4Mux_v I__8523 (
            .O(N__49212),
            .I(N__49200));
    Span4Mux_h I__8522 (
            .O(N__49209),
            .I(N__49197));
    LocalMux I__8521 (
            .O(N__49204),
            .I(N__49194));
    InMux I__8520 (
            .O(N__49203),
            .I(N__49191));
    Odrv4 I__8519 (
            .O(N__49200),
            .I(\pid_front.error_d_reg_prevZ0Z_11 ));
    Odrv4 I__8518 (
            .O(N__49197),
            .I(\pid_front.error_d_reg_prevZ0Z_11 ));
    Odrv4 I__8517 (
            .O(N__49194),
            .I(\pid_front.error_d_reg_prevZ0Z_11 ));
    LocalMux I__8516 (
            .O(N__49191),
            .I(\pid_front.error_d_reg_prevZ0Z_11 ));
    InMux I__8515 (
            .O(N__49182),
            .I(N__49178));
    InMux I__8514 (
            .O(N__49181),
            .I(N__49174));
    LocalMux I__8513 (
            .O(N__49178),
            .I(N__49171));
    InMux I__8512 (
            .O(N__49177),
            .I(N__49168));
    LocalMux I__8511 (
            .O(N__49174),
            .I(N__49164));
    Span4Mux_h I__8510 (
            .O(N__49171),
            .I(N__49161));
    LocalMux I__8509 (
            .O(N__49168),
            .I(N__49158));
    CascadeMux I__8508 (
            .O(N__49167),
            .I(N__49155));
    Span4Mux_h I__8507 (
            .O(N__49164),
            .I(N__49147));
    Span4Mux_v I__8506 (
            .O(N__49161),
            .I(N__49147));
    Span4Mux_h I__8505 (
            .O(N__49158),
            .I(N__49147));
    InMux I__8504 (
            .O(N__49155),
            .I(N__49142));
    InMux I__8503 (
            .O(N__49154),
            .I(N__49142));
    Odrv4 I__8502 (
            .O(N__49147),
            .I(\pid_front.error_d_regZ0Z_11 ));
    LocalMux I__8501 (
            .O(N__49142),
            .I(\pid_front.error_d_regZ0Z_11 ));
    InMux I__8500 (
            .O(N__49137),
            .I(N__49133));
    CascadeMux I__8499 (
            .O(N__49136),
            .I(N__49130));
    LocalMux I__8498 (
            .O(N__49133),
            .I(N__49125));
    InMux I__8497 (
            .O(N__49130),
            .I(N__49122));
    InMux I__8496 (
            .O(N__49129),
            .I(N__49119));
    InMux I__8495 (
            .O(N__49128),
            .I(N__49115));
    Span4Mux_h I__8494 (
            .O(N__49125),
            .I(N__49108));
    LocalMux I__8493 (
            .O(N__49122),
            .I(N__49108));
    LocalMux I__8492 (
            .O(N__49119),
            .I(N__49108));
    InMux I__8491 (
            .O(N__49118),
            .I(N__49105));
    LocalMux I__8490 (
            .O(N__49115),
            .I(N__49102));
    Span4Mux_v I__8489 (
            .O(N__49108),
            .I(N__49099));
    LocalMux I__8488 (
            .O(N__49105),
            .I(N__49096));
    Span4Mux_v I__8487 (
            .O(N__49102),
            .I(N__49091));
    Span4Mux_h I__8486 (
            .O(N__49099),
            .I(N__49091));
    Sp12to4 I__8485 (
            .O(N__49096),
            .I(N__49088));
    Span4Mux_h I__8484 (
            .O(N__49091),
            .I(N__49085));
    Span12Mux_v I__8483 (
            .O(N__49088),
            .I(N__49082));
    Span4Mux_v I__8482 (
            .O(N__49085),
            .I(N__49079));
    Odrv12 I__8481 (
            .O(N__49082),
            .I(\pid_front.error_p_regZ0Z_11 ));
    Odrv4 I__8480 (
            .O(N__49079),
            .I(\pid_front.error_p_regZ0Z_11 ));
    InMux I__8479 (
            .O(N__49074),
            .I(N__49071));
    LocalMux I__8478 (
            .O(N__49071),
            .I(N__49068));
    Odrv4 I__8477 (
            .O(N__49068),
            .I(\pid_front.g0_1_0 ));
    InMux I__8476 (
            .O(N__49065),
            .I(N__49062));
    LocalMux I__8475 (
            .O(N__49062),
            .I(N__49059));
    Span12Mux_h I__8474 (
            .O(N__49059),
            .I(N__49056));
    Odrv12 I__8473 (
            .O(N__49056),
            .I(\pid_front.O_6 ));
    InMux I__8472 (
            .O(N__49053),
            .I(N__49044));
    InMux I__8471 (
            .O(N__49052),
            .I(N__49044));
    InMux I__8470 (
            .O(N__49051),
            .I(N__49044));
    LocalMux I__8469 (
            .O(N__49044),
            .I(N__49041));
    Span4Mux_v I__8468 (
            .O(N__49041),
            .I(N__49038));
    Odrv4 I__8467 (
            .O(N__49038),
            .I(\pid_front.error_d_regZ0Z_4 ));
    InMux I__8466 (
            .O(N__49035),
            .I(N__49032));
    LocalMux I__8465 (
            .O(N__49032),
            .I(N__49029));
    Span12Mux_h I__8464 (
            .O(N__49029),
            .I(N__49026));
    Odrv12 I__8463 (
            .O(N__49026),
            .I(\pid_front.O_7 ));
    InMux I__8462 (
            .O(N__49023),
            .I(N__49016));
    InMux I__8461 (
            .O(N__49022),
            .I(N__49009));
    InMux I__8460 (
            .O(N__49021),
            .I(N__49009));
    InMux I__8459 (
            .O(N__49020),
            .I(N__49009));
    InMux I__8458 (
            .O(N__49019),
            .I(N__49006));
    LocalMux I__8457 (
            .O(N__49016),
            .I(N__49001));
    LocalMux I__8456 (
            .O(N__49009),
            .I(N__49001));
    LocalMux I__8455 (
            .O(N__49006),
            .I(N__48996));
    Span4Mux_v I__8454 (
            .O(N__49001),
            .I(N__48996));
    Odrv4 I__8453 (
            .O(N__48996),
            .I(\pid_front.error_d_regZ0Z_5 ));
    InMux I__8452 (
            .O(N__48993),
            .I(N__48990));
    LocalMux I__8451 (
            .O(N__48990),
            .I(N__48987));
    Span4Mux_v I__8450 (
            .O(N__48987),
            .I(N__48984));
    Span4Mux_h I__8449 (
            .O(N__48984),
            .I(N__48981));
    Span4Mux_h I__8448 (
            .O(N__48981),
            .I(N__48978));
    Span4Mux_h I__8447 (
            .O(N__48978),
            .I(N__48975));
    Odrv4 I__8446 (
            .O(N__48975),
            .I(\pid_front.O_8 ));
    CascadeMux I__8445 (
            .O(N__48972),
            .I(N__48964));
    InMux I__8444 (
            .O(N__48971),
            .I(N__48960));
    InMux I__8443 (
            .O(N__48970),
            .I(N__48955));
    InMux I__8442 (
            .O(N__48969),
            .I(N__48955));
    InMux I__8441 (
            .O(N__48968),
            .I(N__48950));
    InMux I__8440 (
            .O(N__48967),
            .I(N__48950));
    InMux I__8439 (
            .O(N__48964),
            .I(N__48945));
    InMux I__8438 (
            .O(N__48963),
            .I(N__48945));
    LocalMux I__8437 (
            .O(N__48960),
            .I(N__48942));
    LocalMux I__8436 (
            .O(N__48955),
            .I(N__48939));
    LocalMux I__8435 (
            .O(N__48950),
            .I(N__48934));
    LocalMux I__8434 (
            .O(N__48945),
            .I(N__48934));
    Span4Mux_h I__8433 (
            .O(N__48942),
            .I(N__48931));
    Span4Mux_v I__8432 (
            .O(N__48939),
            .I(N__48926));
    Span4Mux_v I__8431 (
            .O(N__48934),
            .I(N__48926));
    Sp12to4 I__8430 (
            .O(N__48931),
            .I(N__48923));
    Span4Mux_v I__8429 (
            .O(N__48926),
            .I(N__48920));
    Span12Mux_v I__8428 (
            .O(N__48923),
            .I(N__48915));
    Sp12to4 I__8427 (
            .O(N__48920),
            .I(N__48915));
    Odrv12 I__8426 (
            .O(N__48915),
            .I(\pid_front.error_p_regZ0Z_12 ));
    CascadeMux I__8425 (
            .O(N__48912),
            .I(\pid_front.N_3_i_1_1_cascade_ ));
    InMux I__8424 (
            .O(N__48909),
            .I(N__48903));
    InMux I__8423 (
            .O(N__48908),
            .I(N__48900));
    InMux I__8422 (
            .O(N__48907),
            .I(N__48897));
    InMux I__8421 (
            .O(N__48906),
            .I(N__48894));
    LocalMux I__8420 (
            .O(N__48903),
            .I(\pid_front.un1_pid_prereg_79 ));
    LocalMux I__8419 (
            .O(N__48900),
            .I(\pid_front.un1_pid_prereg_79 ));
    LocalMux I__8418 (
            .O(N__48897),
            .I(\pid_front.un1_pid_prereg_79 ));
    LocalMux I__8417 (
            .O(N__48894),
            .I(\pid_front.un1_pid_prereg_79 ));
    InMux I__8416 (
            .O(N__48885),
            .I(N__48876));
    InMux I__8415 (
            .O(N__48884),
            .I(N__48869));
    InMux I__8414 (
            .O(N__48883),
            .I(N__48869));
    InMux I__8413 (
            .O(N__48882),
            .I(N__48869));
    InMux I__8412 (
            .O(N__48881),
            .I(N__48866));
    InMux I__8411 (
            .O(N__48880),
            .I(N__48861));
    InMux I__8410 (
            .O(N__48879),
            .I(N__48861));
    LocalMux I__8409 (
            .O(N__48876),
            .I(N__48858));
    LocalMux I__8408 (
            .O(N__48869),
            .I(N__48853));
    LocalMux I__8407 (
            .O(N__48866),
            .I(N__48853));
    LocalMux I__8406 (
            .O(N__48861),
            .I(N__48850));
    Span4Mux_v I__8405 (
            .O(N__48858),
            .I(N__48845));
    Span4Mux_h I__8404 (
            .O(N__48853),
            .I(N__48845));
    Span4Mux_v I__8403 (
            .O(N__48850),
            .I(N__48842));
    Span4Mux_h I__8402 (
            .O(N__48845),
            .I(N__48839));
    Span4Mux_h I__8401 (
            .O(N__48842),
            .I(N__48836));
    Span4Mux_h I__8400 (
            .O(N__48839),
            .I(N__48833));
    Span4Mux_h I__8399 (
            .O(N__48836),
            .I(N__48830));
    Span4Mux_v I__8398 (
            .O(N__48833),
            .I(N__48827));
    Odrv4 I__8397 (
            .O(N__48830),
            .I(\pid_front.error_p_regZ0Z_13 ));
    Odrv4 I__8396 (
            .O(N__48827),
            .I(\pid_front.error_p_regZ0Z_13 ));
    CascadeMux I__8395 (
            .O(N__48822),
            .I(N__48817));
    InMux I__8394 (
            .O(N__48821),
            .I(N__48809));
    InMux I__8393 (
            .O(N__48820),
            .I(N__48809));
    InMux I__8392 (
            .O(N__48817),
            .I(N__48802));
    InMux I__8391 (
            .O(N__48816),
            .I(N__48802));
    InMux I__8390 (
            .O(N__48815),
            .I(N__48802));
    InMux I__8389 (
            .O(N__48814),
            .I(N__48799));
    LocalMux I__8388 (
            .O(N__48809),
            .I(N__48796));
    LocalMux I__8387 (
            .O(N__48802),
            .I(N__48790));
    LocalMux I__8386 (
            .O(N__48799),
            .I(N__48790));
    Span4Mux_h I__8385 (
            .O(N__48796),
            .I(N__48787));
    InMux I__8384 (
            .O(N__48795),
            .I(N__48784));
    Span4Mux_h I__8383 (
            .O(N__48790),
            .I(N__48781));
    Odrv4 I__8382 (
            .O(N__48787),
            .I(\pid_front.error_d_reg_prevZ0Z_13 ));
    LocalMux I__8381 (
            .O(N__48784),
            .I(\pid_front.error_d_reg_prevZ0Z_13 ));
    Odrv4 I__8380 (
            .O(N__48781),
            .I(\pid_front.error_d_reg_prevZ0Z_13 ));
    InMux I__8379 (
            .O(N__48774),
            .I(N__48762));
    InMux I__8378 (
            .O(N__48773),
            .I(N__48762));
    InMux I__8377 (
            .O(N__48772),
            .I(N__48755));
    InMux I__8376 (
            .O(N__48771),
            .I(N__48755));
    InMux I__8375 (
            .O(N__48770),
            .I(N__48755));
    InMux I__8374 (
            .O(N__48769),
            .I(N__48752));
    InMux I__8373 (
            .O(N__48768),
            .I(N__48747));
    InMux I__8372 (
            .O(N__48767),
            .I(N__48747));
    LocalMux I__8371 (
            .O(N__48762),
            .I(N__48740));
    LocalMux I__8370 (
            .O(N__48755),
            .I(N__48740));
    LocalMux I__8369 (
            .O(N__48752),
            .I(N__48740));
    LocalMux I__8368 (
            .O(N__48747),
            .I(\pid_front.error_d_regZ0Z_13 ));
    Odrv4 I__8367 (
            .O(N__48740),
            .I(\pid_front.error_d_regZ0Z_13 ));
    CascadeMux I__8366 (
            .O(N__48735),
            .I(\pid_front.N_2198_0_cascade_ ));
    InMux I__8365 (
            .O(N__48732),
            .I(N__48729));
    LocalMux I__8364 (
            .O(N__48729),
            .I(\pid_front.N_5_0 ));
    InMux I__8363 (
            .O(N__48726),
            .I(N__48723));
    LocalMux I__8362 (
            .O(N__48723),
            .I(\pid_front.N_5_0_0 ));
    CascadeMux I__8361 (
            .O(N__48720),
            .I(\pid_front.g0_2_cascade_ ));
    InMux I__8360 (
            .O(N__48717),
            .I(N__48714));
    LocalMux I__8359 (
            .O(N__48714),
            .I(N__48711));
    Odrv4 I__8358 (
            .O(N__48711),
            .I(\pid_front.N_3_i_1 ));
    CascadeMux I__8357 (
            .O(N__48708),
            .I(\pid_front.error_p_reg_esr_RNI6D5L7Z0Z_12_cascade_ ));
    InMux I__8356 (
            .O(N__48705),
            .I(N__48702));
    LocalMux I__8355 (
            .O(N__48702),
            .I(\pid_front.error_d_reg_prev_esr_RNI6J3B5Z0Z_12 ));
    InMux I__8354 (
            .O(N__48699),
            .I(N__48696));
    LocalMux I__8353 (
            .O(N__48696),
            .I(N__48692));
    InMux I__8352 (
            .O(N__48695),
            .I(N__48689));
    Span4Mux_h I__8351 (
            .O(N__48692),
            .I(N__48686));
    LocalMux I__8350 (
            .O(N__48689),
            .I(N__48683));
    Span4Mux_v I__8349 (
            .O(N__48686),
            .I(N__48680));
    Span4Mux_h I__8348 (
            .O(N__48683),
            .I(N__48677));
    Odrv4 I__8347 (
            .O(N__48680),
            .I(\pid_front.un1_pid_prereg_0_axb_14 ));
    Odrv4 I__8346 (
            .O(N__48677),
            .I(\pid_front.un1_pid_prereg_0_axb_14 ));
    CascadeMux I__8345 (
            .O(N__48672),
            .I(N__48668));
    InMux I__8344 (
            .O(N__48671),
            .I(N__48664));
    InMux I__8343 (
            .O(N__48668),
            .I(N__48659));
    InMux I__8342 (
            .O(N__48667),
            .I(N__48659));
    LocalMux I__8341 (
            .O(N__48664),
            .I(N__48654));
    LocalMux I__8340 (
            .O(N__48659),
            .I(N__48649));
    CascadeMux I__8339 (
            .O(N__48658),
            .I(N__48646));
    InMux I__8338 (
            .O(N__48657),
            .I(N__48642));
    Span4Mux_v I__8337 (
            .O(N__48654),
            .I(N__48639));
    InMux I__8336 (
            .O(N__48653),
            .I(N__48634));
    InMux I__8335 (
            .O(N__48652),
            .I(N__48634));
    Span4Mux_h I__8334 (
            .O(N__48649),
            .I(N__48631));
    InMux I__8333 (
            .O(N__48646),
            .I(N__48626));
    InMux I__8332 (
            .O(N__48645),
            .I(N__48626));
    LocalMux I__8331 (
            .O(N__48642),
            .I(\pid_front.error_d_reg_prevZ0Z_12 ));
    Odrv4 I__8330 (
            .O(N__48639),
            .I(\pid_front.error_d_reg_prevZ0Z_12 ));
    LocalMux I__8329 (
            .O(N__48634),
            .I(\pid_front.error_d_reg_prevZ0Z_12 ));
    Odrv4 I__8328 (
            .O(N__48631),
            .I(\pid_front.error_d_reg_prevZ0Z_12 ));
    LocalMux I__8327 (
            .O(N__48626),
            .I(\pid_front.error_d_reg_prevZ0Z_12 ));
    InMux I__8326 (
            .O(N__48615),
            .I(N__48611));
    InMux I__8325 (
            .O(N__48614),
            .I(N__48608));
    LocalMux I__8324 (
            .O(N__48611),
            .I(N__48605));
    LocalMux I__8323 (
            .O(N__48608),
            .I(\pid_front.error_d_reg_fast_esr_RNIQSG63Z0Z_12 ));
    Odrv4 I__8322 (
            .O(N__48605),
            .I(\pid_front.error_d_reg_fast_esr_RNIQSG63Z0Z_12 ));
    InMux I__8321 (
            .O(N__48600),
            .I(N__48597));
    LocalMux I__8320 (
            .O(N__48597),
            .I(\pid_front.N_5 ));
    InMux I__8319 (
            .O(N__48594),
            .I(N__48588));
    InMux I__8318 (
            .O(N__48593),
            .I(N__48588));
    LocalMux I__8317 (
            .O(N__48588),
            .I(\pid_front.error_d_reg_prevZ0Z_20 ));
    CascadeMux I__8316 (
            .O(N__48585),
            .I(N__48582));
    InMux I__8315 (
            .O(N__48582),
            .I(N__48576));
    InMux I__8314 (
            .O(N__48581),
            .I(N__48576));
    LocalMux I__8313 (
            .O(N__48576),
            .I(\pid_front.error_d_reg_prevZ0Z_21 ));
    InMux I__8312 (
            .O(N__48573),
            .I(N__48570));
    LocalMux I__8311 (
            .O(N__48570),
            .I(N__48564));
    InMux I__8310 (
            .O(N__48569),
            .I(N__48557));
    InMux I__8309 (
            .O(N__48568),
            .I(N__48557));
    InMux I__8308 (
            .O(N__48567),
            .I(N__48557));
    Span4Mux_h I__8307 (
            .O(N__48564),
            .I(N__48552));
    LocalMux I__8306 (
            .O(N__48557),
            .I(N__48552));
    Odrv4 I__8305 (
            .O(N__48552),
            .I(\pid_front.error_d_reg_prevZ0Z_5 ));
    InMux I__8304 (
            .O(N__48549),
            .I(N__48542));
    InMux I__8303 (
            .O(N__48548),
            .I(N__48542));
    InMux I__8302 (
            .O(N__48547),
            .I(N__48539));
    LocalMux I__8301 (
            .O(N__48542),
            .I(N__48536));
    LocalMux I__8300 (
            .O(N__48539),
            .I(N__48533));
    Odrv4 I__8299 (
            .O(N__48536),
            .I(\pid_front.error_d_reg_prevZ0Z_8 ));
    Odrv12 I__8298 (
            .O(N__48533),
            .I(\pid_front.error_d_reg_prevZ0Z_8 ));
    InMux I__8297 (
            .O(N__48528),
            .I(N__48525));
    LocalMux I__8296 (
            .O(N__48525),
            .I(N__48519));
    InMux I__8295 (
            .O(N__48524),
            .I(N__48514));
    InMux I__8294 (
            .O(N__48523),
            .I(N__48514));
    InMux I__8293 (
            .O(N__48522),
            .I(N__48511));
    Span4Mux_h I__8292 (
            .O(N__48519),
            .I(N__48508));
    LocalMux I__8291 (
            .O(N__48514),
            .I(N__48505));
    LocalMux I__8290 (
            .O(N__48511),
            .I(\pid_front.error_d_reg_prev_fastZ0Z_12 ));
    Odrv4 I__8289 (
            .O(N__48508),
            .I(\pid_front.error_d_reg_prev_fastZ0Z_12 ));
    Odrv4 I__8288 (
            .O(N__48505),
            .I(\pid_front.error_d_reg_prev_fastZ0Z_12 ));
    InMux I__8287 (
            .O(N__48498),
            .I(N__48495));
    LocalMux I__8286 (
            .O(N__48495),
            .I(N__48492));
    Odrv12 I__8285 (
            .O(N__48492),
            .I(\dron_frame_decoder_1.drone_H_disp_side_8 ));
    InMux I__8284 (
            .O(N__48489),
            .I(N__48486));
    LocalMux I__8283 (
            .O(N__48486),
            .I(N__48483));
    Odrv12 I__8282 (
            .O(N__48483),
            .I(\dron_frame_decoder_1.drone_H_disp_side_9 ));
    CEMux I__8281 (
            .O(N__48480),
            .I(N__48477));
    LocalMux I__8280 (
            .O(N__48477),
            .I(N__48474));
    Span4Mux_v I__8279 (
            .O(N__48474),
            .I(N__48471));
    Odrv4 I__8278 (
            .O(N__48471),
            .I(\dron_frame_decoder_1.N_716_0 ));
    CascadeMux I__8277 (
            .O(N__48468),
            .I(N__48465));
    InMux I__8276 (
            .O(N__48465),
            .I(N__48462));
    LocalMux I__8275 (
            .O(N__48462),
            .I(N__48459));
    Span4Mux_h I__8274 (
            .O(N__48459),
            .I(N__48454));
    InMux I__8273 (
            .O(N__48458),
            .I(N__48449));
    InMux I__8272 (
            .O(N__48457),
            .I(N__48449));
    Span4Mux_h I__8271 (
            .O(N__48454),
            .I(N__48443));
    LocalMux I__8270 (
            .O(N__48449),
            .I(N__48443));
    InMux I__8269 (
            .O(N__48448),
            .I(N__48440));
    Odrv4 I__8268 (
            .O(N__48443),
            .I(\pid_alt.error_i_acumm7lto5 ));
    LocalMux I__8267 (
            .O(N__48440),
            .I(\pid_alt.error_i_acumm7lto5 ));
    InMux I__8266 (
            .O(N__48435),
            .I(N__48432));
    LocalMux I__8265 (
            .O(N__48432),
            .I(N__48429));
    Span12Mux_h I__8264 (
            .O(N__48429),
            .I(N__48421));
    InMux I__8263 (
            .O(N__48428),
            .I(N__48410));
    InMux I__8262 (
            .O(N__48427),
            .I(N__48410));
    InMux I__8261 (
            .O(N__48426),
            .I(N__48410));
    InMux I__8260 (
            .O(N__48425),
            .I(N__48410));
    InMux I__8259 (
            .O(N__48424),
            .I(N__48410));
    Odrv12 I__8258 (
            .O(N__48421),
            .I(\pid_alt.N_62_mux ));
    LocalMux I__8257 (
            .O(N__48410),
            .I(\pid_alt.N_62_mux ));
    InMux I__8256 (
            .O(N__48405),
            .I(N__48402));
    LocalMux I__8255 (
            .O(N__48402),
            .I(N__48399));
    Span4Mux_v I__8254 (
            .O(N__48399),
            .I(N__48395));
    InMux I__8253 (
            .O(N__48398),
            .I(N__48392));
    Span4Mux_h I__8252 (
            .O(N__48395),
            .I(N__48389));
    LocalMux I__8251 (
            .O(N__48392),
            .I(N__48384));
    Span4Mux_h I__8250 (
            .O(N__48389),
            .I(N__48384));
    Odrv4 I__8249 (
            .O(N__48384),
            .I(\pid_alt.error_i_acummZ0Z_5 ));
    InMux I__8248 (
            .O(N__48381),
            .I(N__48378));
    LocalMux I__8247 (
            .O(N__48378),
            .I(N__48375));
    Odrv12 I__8246 (
            .O(N__48375),
            .I(\pid_front.error_d_reg_prev_esr_RNIBTE61_0Z0Z_21 ));
    CascadeMux I__8245 (
            .O(N__48372),
            .I(\pid_front.error_d_reg_prev_esr_RNIBTE61_0Z0Z_21_cascade_ ));
    InMux I__8244 (
            .O(N__48369),
            .I(N__48364));
    InMux I__8243 (
            .O(N__48368),
            .I(N__48359));
    InMux I__8242 (
            .O(N__48367),
            .I(N__48359));
    LocalMux I__8241 (
            .O(N__48364),
            .I(\pid_front.un1_pid_prereg_0_12 ));
    LocalMux I__8240 (
            .O(N__48359),
            .I(\pid_front.un1_pid_prereg_0_12 ));
    InMux I__8239 (
            .O(N__48354),
            .I(N__48351));
    LocalMux I__8238 (
            .O(N__48351),
            .I(N__48347));
    InMux I__8237 (
            .O(N__48350),
            .I(N__48344));
    Odrv4 I__8236 (
            .O(N__48347),
            .I(\pid_front.error_p_reg_esr_RNI8QE61Z0Z_20 ));
    LocalMux I__8235 (
            .O(N__48344),
            .I(\pid_front.error_p_reg_esr_RNI8QE61Z0Z_20 ));
    InMux I__8234 (
            .O(N__48339),
            .I(N__48327));
    InMux I__8233 (
            .O(N__48338),
            .I(N__48327));
    InMux I__8232 (
            .O(N__48337),
            .I(N__48327));
    InMux I__8231 (
            .O(N__48336),
            .I(N__48324));
    CascadeMux I__8230 (
            .O(N__48335),
            .I(N__48321));
    CascadeMux I__8229 (
            .O(N__48334),
            .I(N__48315));
    LocalMux I__8228 (
            .O(N__48327),
            .I(N__48304));
    LocalMux I__8227 (
            .O(N__48324),
            .I(N__48304));
    InMux I__8226 (
            .O(N__48321),
            .I(N__48295));
    InMux I__8225 (
            .O(N__48320),
            .I(N__48295));
    InMux I__8224 (
            .O(N__48319),
            .I(N__48295));
    InMux I__8223 (
            .O(N__48318),
            .I(N__48295));
    InMux I__8222 (
            .O(N__48315),
            .I(N__48288));
    InMux I__8221 (
            .O(N__48314),
            .I(N__48288));
    InMux I__8220 (
            .O(N__48313),
            .I(N__48288));
    InMux I__8219 (
            .O(N__48312),
            .I(N__48283));
    InMux I__8218 (
            .O(N__48311),
            .I(N__48283));
    InMux I__8217 (
            .O(N__48310),
            .I(N__48278));
    InMux I__8216 (
            .O(N__48309),
            .I(N__48278));
    Span4Mux_v I__8215 (
            .O(N__48304),
            .I(N__48275));
    LocalMux I__8214 (
            .O(N__48295),
            .I(N__48270));
    LocalMux I__8213 (
            .O(N__48288),
            .I(N__48270));
    LocalMux I__8212 (
            .O(N__48283),
            .I(N__48265));
    LocalMux I__8211 (
            .O(N__48278),
            .I(N__48265));
    Span4Mux_h I__8210 (
            .O(N__48275),
            .I(N__48262));
    Span4Mux_v I__8209 (
            .O(N__48270),
            .I(N__48257));
    Span4Mux_h I__8208 (
            .O(N__48265),
            .I(N__48257));
    Span4Mux_h I__8207 (
            .O(N__48262),
            .I(N__48254));
    Span4Mux_h I__8206 (
            .O(N__48257),
            .I(N__48251));
    Span4Mux_v I__8205 (
            .O(N__48254),
            .I(N__48248));
    Span4Mux_v I__8204 (
            .O(N__48251),
            .I(N__48245));
    Odrv4 I__8203 (
            .O(N__48248),
            .I(\pid_front.error_p_regZ0Z_21 ));
    Odrv4 I__8202 (
            .O(N__48245),
            .I(\pid_front.error_p_regZ0Z_21 ));
    CascadeMux I__8201 (
            .O(N__48240),
            .I(N__48237));
    InMux I__8200 (
            .O(N__48237),
            .I(N__48231));
    InMux I__8199 (
            .O(N__48236),
            .I(N__48231));
    LocalMux I__8198 (
            .O(N__48231),
            .I(\pid_front.error_d_reg_prev_esr_RNIBTE61Z0Z_21 ));
    InMux I__8197 (
            .O(N__48228),
            .I(N__48222));
    InMux I__8196 (
            .O(N__48227),
            .I(N__48222));
    LocalMux I__8195 (
            .O(N__48222),
            .I(N__48219));
    Span4Mux_h I__8194 (
            .O(N__48219),
            .I(N__48216));
    Span4Mux_h I__8193 (
            .O(N__48216),
            .I(N__48213));
    Span4Mux_v I__8192 (
            .O(N__48213),
            .I(N__48210));
    Odrv4 I__8191 (
            .O(N__48210),
            .I(\pid_front.error_p_regZ0Z_20 ));
    InMux I__8190 (
            .O(N__48207),
            .I(N__48201));
    InMux I__8189 (
            .O(N__48206),
            .I(N__48201));
    LocalMux I__8188 (
            .O(N__48201),
            .I(N__48198));
    Odrv4 I__8187 (
            .O(N__48198),
            .I(\pid_front.error_p_reg_esr_RNI8QE61_0Z0Z_20 ));
    InMux I__8186 (
            .O(N__48195),
            .I(N__48192));
    LocalMux I__8185 (
            .O(N__48192),
            .I(N__48189));
    Span4Mux_h I__8184 (
            .O(N__48189),
            .I(N__48186));
    Odrv4 I__8183 (
            .O(N__48186),
            .I(\dron_frame_decoder_1.drone_H_disp_side_10 ));
    InMux I__8182 (
            .O(N__48183),
            .I(N__48180));
    LocalMux I__8181 (
            .O(N__48180),
            .I(\pid_front.error_p_reg_esr_RNIBG6FZ0Z_7 ));
    InMux I__8180 (
            .O(N__48177),
            .I(N__48171));
    InMux I__8179 (
            .O(N__48176),
            .I(N__48171));
    LocalMux I__8178 (
            .O(N__48171),
            .I(\pid_front.error_p_reg_esr_RNIGL6F_0Z0Z_8 ));
    InMux I__8177 (
            .O(N__48168),
            .I(N__48164));
    CascadeMux I__8176 (
            .O(N__48167),
            .I(N__48161));
    LocalMux I__8175 (
            .O(N__48164),
            .I(N__48158));
    InMux I__8174 (
            .O(N__48161),
            .I(N__48155));
    Span4Mux_h I__8173 (
            .O(N__48158),
            .I(N__48150));
    LocalMux I__8172 (
            .O(N__48155),
            .I(N__48150));
    Span4Mux_v I__8171 (
            .O(N__48150),
            .I(N__48147));
    Odrv4 I__8170 (
            .O(N__48147),
            .I(\pid_front.error_p_reg_esr_RNICU3D1Z0Z_6 ));
    CascadeMux I__8169 (
            .O(N__48144),
            .I(\pid_front.error_p_reg_esr_RNIBG6FZ0Z_7_cascade_ ));
    InMux I__8168 (
            .O(N__48141),
            .I(N__48138));
    LocalMux I__8167 (
            .O(N__48138),
            .I(N__48135));
    Span4Mux_v I__8166 (
            .O(N__48135),
            .I(N__48132));
    Odrv4 I__8165 (
            .O(N__48132),
            .I(\pid_front.error_p_reg_esr_RNI5B9Q2Z0Z_7 ));
    InMux I__8164 (
            .O(N__48129),
            .I(N__48126));
    LocalMux I__8163 (
            .O(N__48126),
            .I(\pid_front.N_2161_i ));
    CascadeMux I__8162 (
            .O(N__48123),
            .I(N__48120));
    InMux I__8161 (
            .O(N__48120),
            .I(N__48114));
    InMux I__8160 (
            .O(N__48119),
            .I(N__48114));
    LocalMux I__8159 (
            .O(N__48114),
            .I(N__48111));
    Span4Mux_v I__8158 (
            .O(N__48111),
            .I(N__48108));
    Sp12to4 I__8157 (
            .O(N__48108),
            .I(N__48105));
    Odrv12 I__8156 (
            .O(N__48105),
            .I(\pid_front.error_p_regZ0Z_7 ));
    InMux I__8155 (
            .O(N__48102),
            .I(N__48095));
    InMux I__8154 (
            .O(N__48101),
            .I(N__48095));
    InMux I__8153 (
            .O(N__48100),
            .I(N__48092));
    LocalMux I__8152 (
            .O(N__48095),
            .I(\pid_front.error_d_reg_prevZ0Z_6 ));
    LocalMux I__8151 (
            .O(N__48092),
            .I(\pid_front.error_d_reg_prevZ0Z_6 ));
    CascadeMux I__8150 (
            .O(N__48087),
            .I(\pid_front.N_2161_i_cascade_ ));
    InMux I__8149 (
            .O(N__48084),
            .I(N__48078));
    InMux I__8148 (
            .O(N__48083),
            .I(N__48078));
    LocalMux I__8147 (
            .O(N__48078),
            .I(N__48075));
    Span4Mux_v I__8146 (
            .O(N__48075),
            .I(N__48072));
    Odrv4 I__8145 (
            .O(N__48072),
            .I(\pid_front.error_p_reg_esr_RNIBG6F_0Z0Z_7 ));
    InMux I__8144 (
            .O(N__48069),
            .I(N__48066));
    LocalMux I__8143 (
            .O(N__48066),
            .I(N__48063));
    Span4Mux_v I__8142 (
            .O(N__48063),
            .I(N__48060));
    Span4Mux_h I__8141 (
            .O(N__48060),
            .I(N__48056));
    InMux I__8140 (
            .O(N__48059),
            .I(N__48053));
    Span4Mux_h I__8139 (
            .O(N__48056),
            .I(N__48050));
    LocalMux I__8138 (
            .O(N__48053),
            .I(N__48047));
    Odrv4 I__8137 (
            .O(N__48050),
            .I(\pid_front.error_p_regZ0Z_8 ));
    Odrv12 I__8136 (
            .O(N__48047),
            .I(\pid_front.error_p_regZ0Z_8 ));
    CascadeMux I__8135 (
            .O(N__48042),
            .I(N__48038));
    InMux I__8134 (
            .O(N__48041),
            .I(N__48034));
    InMux I__8133 (
            .O(N__48038),
            .I(N__48029));
    InMux I__8132 (
            .O(N__48037),
            .I(N__48029));
    LocalMux I__8131 (
            .O(N__48034),
            .I(\pid_front.error_d_reg_prevZ0Z_7 ));
    LocalMux I__8130 (
            .O(N__48029),
            .I(\pid_front.error_d_reg_prevZ0Z_7 ));
    InMux I__8129 (
            .O(N__48024),
            .I(N__48021));
    LocalMux I__8128 (
            .O(N__48021),
            .I(\pid_front.N_2167_i ));
    InMux I__8127 (
            .O(N__48018),
            .I(N__48014));
    InMux I__8126 (
            .O(N__48017),
            .I(N__48011));
    LocalMux I__8125 (
            .O(N__48014),
            .I(N__48008));
    LocalMux I__8124 (
            .O(N__48011),
            .I(N__48005));
    Span4Mux_h I__8123 (
            .O(N__48008),
            .I(N__48002));
    Odrv4 I__8122 (
            .O(N__48005),
            .I(\pid_front.error_p_reg_esr_RNIGL6FZ0Z_8 ));
    Odrv4 I__8121 (
            .O(N__48002),
            .I(\pid_front.error_p_reg_esr_RNIGL6FZ0Z_8 ));
    IoInMux I__8120 (
            .O(N__47997),
            .I(N__47993));
    CascadeMux I__8119 (
            .O(N__47996),
            .I(N__47983));
    LocalMux I__8118 (
            .O(N__47993),
            .I(N__47979));
    InMux I__8117 (
            .O(N__47992),
            .I(N__47961));
    InMux I__8116 (
            .O(N__47991),
            .I(N__47961));
    InMux I__8115 (
            .O(N__47990),
            .I(N__47961));
    InMux I__8114 (
            .O(N__47989),
            .I(N__47961));
    InMux I__8113 (
            .O(N__47988),
            .I(N__47961));
    InMux I__8112 (
            .O(N__47987),
            .I(N__47961));
    InMux I__8111 (
            .O(N__47986),
            .I(N__47961));
    InMux I__8110 (
            .O(N__47983),
            .I(N__47961));
    InMux I__8109 (
            .O(N__47982),
            .I(N__47958));
    IoSpan4Mux I__8108 (
            .O(N__47979),
            .I(N__47955));
    CascadeMux I__8107 (
            .O(N__47978),
            .I(N__47952));
    LocalMux I__8106 (
            .O(N__47961),
            .I(N__47947));
    LocalMux I__8105 (
            .O(N__47958),
            .I(N__47944));
    Span4Mux_s1_v I__8104 (
            .O(N__47955),
            .I(N__47940));
    InMux I__8103 (
            .O(N__47952),
            .I(N__47935));
    InMux I__8102 (
            .O(N__47951),
            .I(N__47935));
    InMux I__8101 (
            .O(N__47950),
            .I(N__47932));
    Span4Mux_v I__8100 (
            .O(N__47947),
            .I(N__47929));
    Span4Mux_h I__8099 (
            .O(N__47944),
            .I(N__47926));
    InMux I__8098 (
            .O(N__47943),
            .I(N__47923));
    Span4Mux_h I__8097 (
            .O(N__47940),
            .I(N__47920));
    LocalMux I__8096 (
            .O(N__47935),
            .I(N__47909));
    LocalMux I__8095 (
            .O(N__47932),
            .I(N__47909));
    Span4Mux_h I__8094 (
            .O(N__47929),
            .I(N__47909));
    Span4Mux_v I__8093 (
            .O(N__47926),
            .I(N__47909));
    LocalMux I__8092 (
            .O(N__47923),
            .I(N__47909));
    Span4Mux_v I__8091 (
            .O(N__47920),
            .I(N__47904));
    Span4Mux_v I__8090 (
            .O(N__47909),
            .I(N__47904));
    Odrv4 I__8089 (
            .O(N__47904),
            .I(debug_CH0_16A_c));
    InMux I__8088 (
            .O(N__47901),
            .I(N__47898));
    LocalMux I__8087 (
            .O(N__47898),
            .I(N__47895));
    Span4Mux_v I__8086 (
            .O(N__47895),
            .I(N__47890));
    InMux I__8085 (
            .O(N__47894),
            .I(N__47885));
    InMux I__8084 (
            .O(N__47893),
            .I(N__47885));
    Odrv4 I__8083 (
            .O(N__47890),
            .I(\uart_drone.data_rdyc_1 ));
    LocalMux I__8082 (
            .O(N__47885),
            .I(\uart_drone.data_rdyc_1 ));
    CascadeMux I__8081 (
            .O(N__47880),
            .I(N__47877));
    InMux I__8080 (
            .O(N__47877),
            .I(N__47865));
    InMux I__8079 (
            .O(N__47876),
            .I(N__47865));
    InMux I__8078 (
            .O(N__47875),
            .I(N__47865));
    InMux I__8077 (
            .O(N__47874),
            .I(N__47865));
    LocalMux I__8076 (
            .O(N__47865),
            .I(\dron_frame_decoder_1.stateZ0Z_5 ));
    CascadeMux I__8075 (
            .O(N__47862),
            .I(N__47857));
    CascadeMux I__8074 (
            .O(N__47861),
            .I(N__47854));
    CascadeMux I__8073 (
            .O(N__47860),
            .I(N__47851));
    InMux I__8072 (
            .O(N__47857),
            .I(N__47846));
    InMux I__8071 (
            .O(N__47854),
            .I(N__47839));
    InMux I__8070 (
            .O(N__47851),
            .I(N__47839));
    InMux I__8069 (
            .O(N__47850),
            .I(N__47839));
    InMux I__8068 (
            .O(N__47849),
            .I(N__47836));
    LocalMux I__8067 (
            .O(N__47846),
            .I(\dron_frame_decoder_1.stateZ0Z_4 ));
    LocalMux I__8066 (
            .O(N__47839),
            .I(\dron_frame_decoder_1.stateZ0Z_4 ));
    LocalMux I__8065 (
            .O(N__47836),
            .I(\dron_frame_decoder_1.stateZ0Z_4 ));
    CascadeMux I__8064 (
            .O(N__47829),
            .I(\dron_frame_decoder_1.state_RNI6P6KZ0Z_4_cascade_ ));
    CascadeMux I__8063 (
            .O(N__47826),
            .I(\pid_front.N_2167_i_cascade_ ));
    InMux I__8062 (
            .O(N__47823),
            .I(N__47817));
    InMux I__8061 (
            .O(N__47822),
            .I(N__47817));
    LocalMux I__8060 (
            .O(N__47817),
            .I(N__47813));
    InMux I__8059 (
            .O(N__47816),
            .I(N__47810));
    Span4Mux_v I__8058 (
            .O(N__47813),
            .I(N__47805));
    LocalMux I__8057 (
            .O(N__47810),
            .I(N__47805));
    Span4Mux_h I__8056 (
            .O(N__47805),
            .I(N__47802));
    Odrv4 I__8055 (
            .O(N__47802),
            .I(\dron_frame_decoder_1.stateZ0Z_2 ));
    CascadeMux I__8054 (
            .O(N__47799),
            .I(N__47795));
    CascadeMux I__8053 (
            .O(N__47798),
            .I(N__47792));
    InMux I__8052 (
            .O(N__47795),
            .I(N__47789));
    InMux I__8051 (
            .O(N__47792),
            .I(N__47786));
    LocalMux I__8050 (
            .O(N__47789),
            .I(N__47781));
    LocalMux I__8049 (
            .O(N__47786),
            .I(N__47781));
    Span4Mux_h I__8048 (
            .O(N__47781),
            .I(N__47778));
    Odrv4 I__8047 (
            .O(N__47778),
            .I(\pid_front.error_p_reg_esr_RNIPC5D1Z0Z_7 ));
    CascadeMux I__8046 (
            .O(N__47775),
            .I(\dron_frame_decoder_1.state_ns_i_a2_1_1Z0Z_0_cascade_ ));
    InMux I__8045 (
            .O(N__47772),
            .I(N__47769));
    LocalMux I__8044 (
            .O(N__47769),
            .I(\dron_frame_decoder_1.N_220 ));
    InMux I__8043 (
            .O(N__47766),
            .I(N__47763));
    LocalMux I__8042 (
            .O(N__47763),
            .I(\dron_frame_decoder_1.N_224 ));
    CascadeMux I__8041 (
            .O(N__47760),
            .I(\dron_frame_decoder_1.N_220_cascade_ ));
    InMux I__8040 (
            .O(N__47757),
            .I(N__47754));
    LocalMux I__8039 (
            .O(N__47754),
            .I(\dron_frame_decoder_1.N_198 ));
    InMux I__8038 (
            .O(N__47751),
            .I(N__47748));
    LocalMux I__8037 (
            .O(N__47748),
            .I(\dron_frame_decoder_1.state_ns_i_a2_0_2_0 ));
    InMux I__8036 (
            .O(N__47745),
            .I(N__47742));
    LocalMux I__8035 (
            .O(N__47742),
            .I(\dron_frame_decoder_1.un1_sink_data_valid_5_i_0 ));
    CascadeMux I__8034 (
            .O(N__47739),
            .I(\dron_frame_decoder_1.un1_sink_data_valid_5_i_0_cascade_ ));
    CascadeMux I__8033 (
            .O(N__47736),
            .I(\dron_frame_decoder_1.state_RNI3T3K1Z0Z_7_cascade_ ));
    CEMux I__8032 (
            .O(N__47733),
            .I(N__47730));
    LocalMux I__8031 (
            .O(N__47730),
            .I(N__47727));
    Span4Mux_v I__8030 (
            .O(N__47727),
            .I(N__47724));
    Span4Mux_h I__8029 (
            .O(N__47724),
            .I(N__47721));
    Odrv4 I__8028 (
            .O(N__47721),
            .I(\dron_frame_decoder_1.N_732_0 ));
    CascadeMux I__8027 (
            .O(N__47718),
            .I(N__47714));
    InMux I__8026 (
            .O(N__47717),
            .I(N__47711));
    InMux I__8025 (
            .O(N__47714),
            .I(N__47708));
    LocalMux I__8024 (
            .O(N__47711),
            .I(\uart_drone.data_AuxZ0Z_2 ));
    LocalMux I__8023 (
            .O(N__47708),
            .I(\uart_drone.data_AuxZ0Z_2 ));
    CascadeMux I__8022 (
            .O(N__47703),
            .I(N__47699));
    InMux I__8021 (
            .O(N__47702),
            .I(N__47696));
    InMux I__8020 (
            .O(N__47699),
            .I(N__47693));
    LocalMux I__8019 (
            .O(N__47696),
            .I(\uart_drone.data_AuxZ0Z_3 ));
    LocalMux I__8018 (
            .O(N__47693),
            .I(\uart_drone.data_AuxZ0Z_3 ));
    CascadeMux I__8017 (
            .O(N__47688),
            .I(N__47684));
    InMux I__8016 (
            .O(N__47687),
            .I(N__47681));
    InMux I__8015 (
            .O(N__47684),
            .I(N__47678));
    LocalMux I__8014 (
            .O(N__47681),
            .I(\uart_drone.data_AuxZ0Z_4 ));
    LocalMux I__8013 (
            .O(N__47678),
            .I(\uart_drone.data_AuxZ0Z_4 ));
    CascadeMux I__8012 (
            .O(N__47673),
            .I(N__47669));
    InMux I__8011 (
            .O(N__47672),
            .I(N__47666));
    InMux I__8010 (
            .O(N__47669),
            .I(N__47663));
    LocalMux I__8009 (
            .O(N__47666),
            .I(\uart_drone.data_AuxZ0Z_5 ));
    LocalMux I__8008 (
            .O(N__47663),
            .I(\uart_drone.data_AuxZ0Z_5 ));
    CascadeMux I__8007 (
            .O(N__47658),
            .I(N__47654));
    InMux I__8006 (
            .O(N__47657),
            .I(N__47651));
    InMux I__8005 (
            .O(N__47654),
            .I(N__47648));
    LocalMux I__8004 (
            .O(N__47651),
            .I(\uart_drone.data_AuxZ0Z_6 ));
    LocalMux I__8003 (
            .O(N__47648),
            .I(\uart_drone.data_AuxZ0Z_6 ));
    CascadeMux I__8002 (
            .O(N__47643),
            .I(N__47639));
    InMux I__8001 (
            .O(N__47642),
            .I(N__47636));
    InMux I__8000 (
            .O(N__47639),
            .I(N__47633));
    LocalMux I__7999 (
            .O(N__47636),
            .I(\uart_drone.data_AuxZ0Z_7 ));
    LocalMux I__7998 (
            .O(N__47633),
            .I(\uart_drone.data_AuxZ0Z_7 ));
    CEMux I__7997 (
            .O(N__47628),
            .I(N__47625));
    LocalMux I__7996 (
            .O(N__47625),
            .I(N__47622));
    Span4Mux_h I__7995 (
            .O(N__47622),
            .I(N__47619));
    Odrv4 I__7994 (
            .O(N__47619),
            .I(\uart_drone.data_rdyc_1_0 ));
    SRMux I__7993 (
            .O(N__47616),
            .I(N__47613));
    LocalMux I__7992 (
            .O(N__47613),
            .I(N__47610));
    Span4Mux_v I__7991 (
            .O(N__47610),
            .I(N__47607));
    Span4Mux_h I__7990 (
            .O(N__47607),
            .I(N__47604));
    Odrv4 I__7989 (
            .O(N__47604),
            .I(\uart_drone.timer_Count_RNIES9Q1Z0Z_2 ));
    CascadeMux I__7988 (
            .O(N__47601),
            .I(\dron_frame_decoder_1.N_230_5_cascade_ ));
    CascadeMux I__7987 (
            .O(N__47598),
            .I(\dron_frame_decoder_1.N_224_cascade_ ));
    InMux I__7986 (
            .O(N__47595),
            .I(N__47592));
    LocalMux I__7985 (
            .O(N__47592),
            .I(\uart_drone.data_Auxce_0_3 ));
    InMux I__7984 (
            .O(N__47589),
            .I(N__47565));
    InMux I__7983 (
            .O(N__47588),
            .I(N__47565));
    InMux I__7982 (
            .O(N__47587),
            .I(N__47565));
    InMux I__7981 (
            .O(N__47586),
            .I(N__47565));
    InMux I__7980 (
            .O(N__47585),
            .I(N__47565));
    InMux I__7979 (
            .O(N__47584),
            .I(N__47565));
    InMux I__7978 (
            .O(N__47583),
            .I(N__47565));
    InMux I__7977 (
            .O(N__47582),
            .I(N__47565));
    LocalMux I__7976 (
            .O(N__47565),
            .I(N__47562));
    Span4Mux_h I__7975 (
            .O(N__47562),
            .I(N__47559));
    Odrv4 I__7974 (
            .O(N__47559),
            .I(\uart_drone.un1_state_2_0 ));
    SRMux I__7973 (
            .O(N__47556),
            .I(N__47553));
    LocalMux I__7972 (
            .O(N__47553),
            .I(N__47550));
    Span4Mux_h I__7971 (
            .O(N__47550),
            .I(N__47547));
    Span4Mux_v I__7970 (
            .O(N__47547),
            .I(N__47544));
    Odrv4 I__7969 (
            .O(N__47544),
            .I(\uart_drone.state_RNIOU0NZ0Z_4 ));
    InMux I__7968 (
            .O(N__47541),
            .I(N__47537));
    InMux I__7967 (
            .O(N__47540),
            .I(N__47534));
    LocalMux I__7966 (
            .O(N__47537),
            .I(\uart_drone.data_AuxZ0Z_0 ));
    LocalMux I__7965 (
            .O(N__47534),
            .I(\uart_drone.data_AuxZ0Z_0 ));
    CascadeMux I__7964 (
            .O(N__47529),
            .I(N__47525));
    InMux I__7963 (
            .O(N__47528),
            .I(N__47522));
    InMux I__7962 (
            .O(N__47525),
            .I(N__47519));
    LocalMux I__7961 (
            .O(N__47522),
            .I(\uart_drone.data_AuxZ0Z_1 ));
    LocalMux I__7960 (
            .O(N__47519),
            .I(\uart_drone.data_AuxZ0Z_1 ));
    InMux I__7959 (
            .O(N__47514),
            .I(\ppm_encoder_1.un1_aileron_cry_6 ));
    InMux I__7958 (
            .O(N__47511),
            .I(N__47508));
    LocalMux I__7957 (
            .O(N__47508),
            .I(N__47505));
    Odrv4 I__7956 (
            .O(N__47505),
            .I(\ppm_encoder_1.un1_aileron_cry_7_THRU_CO ));
    InMux I__7955 (
            .O(N__47502),
            .I(bfn_11_10_0_));
    InMux I__7954 (
            .O(N__47499),
            .I(N__47496));
    LocalMux I__7953 (
            .O(N__47496),
            .I(\ppm_encoder_1.un1_aileron_cry_8_THRU_CO ));
    InMux I__7952 (
            .O(N__47493),
            .I(\ppm_encoder_1.un1_aileron_cry_8 ));
    InMux I__7951 (
            .O(N__47490),
            .I(N__47487));
    LocalMux I__7950 (
            .O(N__47487),
            .I(N__47484));
    Span4Mux_h I__7949 (
            .O(N__47484),
            .I(N__47481));
    Odrv4 I__7948 (
            .O(N__47481),
            .I(\ppm_encoder_1.un1_aileron_cry_9_THRU_CO ));
    InMux I__7947 (
            .O(N__47478),
            .I(\ppm_encoder_1.un1_aileron_cry_9 ));
    InMux I__7946 (
            .O(N__47475),
            .I(N__47472));
    LocalMux I__7945 (
            .O(N__47472),
            .I(N__47469));
    Odrv4 I__7944 (
            .O(N__47469),
            .I(\ppm_encoder_1.un1_aileron_cry_10_THRU_CO ));
    InMux I__7943 (
            .O(N__47466),
            .I(\ppm_encoder_1.un1_aileron_cry_10 ));
    InMux I__7942 (
            .O(N__47463),
            .I(\ppm_encoder_1.un1_aileron_cry_11 ));
    InMux I__7941 (
            .O(N__47460),
            .I(N__47457));
    LocalMux I__7940 (
            .O(N__47457),
            .I(N__47454));
    Odrv4 I__7939 (
            .O(N__47454),
            .I(\ppm_encoder_1.un1_aileron_cry_12_THRU_CO ));
    InMux I__7938 (
            .O(N__47451),
            .I(\ppm_encoder_1.un1_aileron_cry_12 ));
    InMux I__7937 (
            .O(N__47448),
            .I(\ppm_encoder_1.un1_aileron_cry_13 ));
    InMux I__7936 (
            .O(N__47445),
            .I(N__47442));
    LocalMux I__7935 (
            .O(N__47442),
            .I(N__47438));
    CascadeMux I__7934 (
            .O(N__47441),
            .I(N__47434));
    Span4Mux_h I__7933 (
            .O(N__47438),
            .I(N__47431));
    InMux I__7932 (
            .O(N__47437),
            .I(N__47428));
    InMux I__7931 (
            .O(N__47434),
            .I(N__47425));
    Span4Mux_v I__7930 (
            .O(N__47431),
            .I(N__47422));
    LocalMux I__7929 (
            .O(N__47428),
            .I(\ppm_encoder_1.aileronZ0Z_8 ));
    LocalMux I__7928 (
            .O(N__47425),
            .I(\ppm_encoder_1.aileronZ0Z_8 ));
    Odrv4 I__7927 (
            .O(N__47422),
            .I(\ppm_encoder_1.aileronZ0Z_8 ));
    InMux I__7926 (
            .O(N__47415),
            .I(N__47411));
    CascadeMux I__7925 (
            .O(N__47414),
            .I(N__47408));
    LocalMux I__7924 (
            .O(N__47411),
            .I(N__47404));
    InMux I__7923 (
            .O(N__47408),
            .I(N__47401));
    InMux I__7922 (
            .O(N__47407),
            .I(N__47398));
    Span4Mux_h I__7921 (
            .O(N__47404),
            .I(N__47395));
    LocalMux I__7920 (
            .O(N__47401),
            .I(\ppm_encoder_1.aileronZ0Z_9 ));
    LocalMux I__7919 (
            .O(N__47398),
            .I(\ppm_encoder_1.aileronZ0Z_9 ));
    Odrv4 I__7918 (
            .O(N__47395),
            .I(\ppm_encoder_1.aileronZ0Z_9 ));
    InMux I__7917 (
            .O(N__47388),
            .I(N__47384));
    CascadeMux I__7916 (
            .O(N__47387),
            .I(N__47380));
    LocalMux I__7915 (
            .O(N__47384),
            .I(N__47377));
    InMux I__7914 (
            .O(N__47383),
            .I(N__47374));
    InMux I__7913 (
            .O(N__47380),
            .I(N__47371));
    Span4Mux_h I__7912 (
            .O(N__47377),
            .I(N__47368));
    LocalMux I__7911 (
            .O(N__47374),
            .I(\ppm_encoder_1.elevatorZ0Z_9 ));
    LocalMux I__7910 (
            .O(N__47371),
            .I(\ppm_encoder_1.elevatorZ0Z_9 ));
    Odrv4 I__7909 (
            .O(N__47368),
            .I(\ppm_encoder_1.elevatorZ0Z_9 ));
    InMux I__7908 (
            .O(N__47361),
            .I(\ppm_encoder_1.un1_aileron_cry_0 ));
    InMux I__7907 (
            .O(N__47358),
            .I(N__47355));
    LocalMux I__7906 (
            .O(N__47355),
            .I(\ppm_encoder_1.un1_aileron_cry_1_THRU_CO ));
    InMux I__7905 (
            .O(N__47352),
            .I(\ppm_encoder_1.un1_aileron_cry_1 ));
    InMux I__7904 (
            .O(N__47349),
            .I(\ppm_encoder_1.un1_aileron_cry_2 ));
    InMux I__7903 (
            .O(N__47346),
            .I(N__47343));
    LocalMux I__7902 (
            .O(N__47343),
            .I(\ppm_encoder_1.un1_aileron_cry_3_THRU_CO ));
    InMux I__7901 (
            .O(N__47340),
            .I(\ppm_encoder_1.un1_aileron_cry_3 ));
    InMux I__7900 (
            .O(N__47337),
            .I(N__47334));
    LocalMux I__7899 (
            .O(N__47334),
            .I(N__47331));
    Span4Mux_v I__7898 (
            .O(N__47331),
            .I(N__47328));
    Odrv4 I__7897 (
            .O(N__47328),
            .I(\ppm_encoder_1.un1_aileron_cry_4_THRU_CO ));
    InMux I__7896 (
            .O(N__47325),
            .I(\ppm_encoder_1.un1_aileron_cry_4 ));
    InMux I__7895 (
            .O(N__47322),
            .I(\ppm_encoder_1.un1_aileron_cry_5 ));
    CascadeMux I__7894 (
            .O(N__47319),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_12_cascade_ ));
    CascadeMux I__7893 (
            .O(N__47316),
            .I(N__47313));
    InMux I__7892 (
            .O(N__47313),
            .I(N__47309));
    InMux I__7891 (
            .O(N__47312),
            .I(N__47306));
    LocalMux I__7890 (
            .O(N__47309),
            .I(N__47301));
    LocalMux I__7889 (
            .O(N__47306),
            .I(N__47301));
    Span4Mux_v I__7888 (
            .O(N__47301),
            .I(N__47298));
    Odrv4 I__7887 (
            .O(N__47298),
            .I(\ppm_encoder_1.N_267_i_i ));
    InMux I__7886 (
            .O(N__47295),
            .I(N__47292));
    LocalMux I__7885 (
            .O(N__47292),
            .I(N__47289));
    Odrv4 I__7884 (
            .O(N__47289),
            .I(\ppm_encoder_1.init_pulses_RNI7OHF5Z0Z_12 ));
    InMux I__7883 (
            .O(N__47286),
            .I(N__47281));
    InMux I__7882 (
            .O(N__47285),
            .I(N__47278));
    InMux I__7881 (
            .O(N__47284),
            .I(N__47275));
    LocalMux I__7880 (
            .O(N__47281),
            .I(N__47272));
    LocalMux I__7879 (
            .O(N__47278),
            .I(\ppm_encoder_1.elevatorZ0Z_12 ));
    LocalMux I__7878 (
            .O(N__47275),
            .I(\ppm_encoder_1.elevatorZ0Z_12 ));
    Odrv4 I__7877 (
            .O(N__47272),
            .I(\ppm_encoder_1.elevatorZ0Z_12 ));
    InMux I__7876 (
            .O(N__47265),
            .I(N__47262));
    LocalMux I__7875 (
            .O(N__47262),
            .I(N__47259));
    Span4Mux_v I__7874 (
            .O(N__47259),
            .I(N__47255));
    InMux I__7873 (
            .O(N__47258),
            .I(N__47252));
    Span4Mux_h I__7872 (
            .O(N__47255),
            .I(N__47249));
    LocalMux I__7871 (
            .O(N__47252),
            .I(N__47246));
    Odrv4 I__7870 (
            .O(N__47249),
            .I(throttle_order_12));
    Odrv12 I__7869 (
            .O(N__47246),
            .I(throttle_order_12));
    InMux I__7868 (
            .O(N__47241),
            .I(N__47238));
    LocalMux I__7867 (
            .O(N__47238),
            .I(N__47235));
    Span4Mux_h I__7866 (
            .O(N__47235),
            .I(N__47232));
    Odrv4 I__7865 (
            .O(N__47232),
            .I(\ppm_encoder_1.un1_throttle_cry_11_THRU_CO ));
    CascadeMux I__7864 (
            .O(N__47229),
            .I(N__47225));
    CascadeMux I__7863 (
            .O(N__47228),
            .I(N__47221));
    InMux I__7862 (
            .O(N__47225),
            .I(N__47218));
    InMux I__7861 (
            .O(N__47224),
            .I(N__47213));
    InMux I__7860 (
            .O(N__47221),
            .I(N__47213));
    LocalMux I__7859 (
            .O(N__47218),
            .I(\ppm_encoder_1.throttleZ0Z_12 ));
    LocalMux I__7858 (
            .O(N__47213),
            .I(\ppm_encoder_1.throttleZ0Z_12 ));
    InMux I__7857 (
            .O(N__47208),
            .I(N__47205));
    LocalMux I__7856 (
            .O(N__47205),
            .I(\ppm_encoder_1.un2_throttle_iv_0_1_12 ));
    InMux I__7855 (
            .O(N__47202),
            .I(N__47199));
    LocalMux I__7854 (
            .O(N__47199),
            .I(N__47196));
    Odrv12 I__7853 (
            .O(N__47196),
            .I(\ppm_encoder_1.un1_throttle_cry_6_THRU_CO ));
    InMux I__7852 (
            .O(N__47193),
            .I(N__47190));
    LocalMux I__7851 (
            .O(N__47190),
            .I(N__47185));
    InMux I__7850 (
            .O(N__47189),
            .I(N__47182));
    CascadeMux I__7849 (
            .O(N__47188),
            .I(N__47179));
    Span4Mux_h I__7848 (
            .O(N__47185),
            .I(N__47174));
    LocalMux I__7847 (
            .O(N__47182),
            .I(N__47174));
    InMux I__7846 (
            .O(N__47179),
            .I(N__47171));
    Span4Mux_h I__7845 (
            .O(N__47174),
            .I(N__47168));
    LocalMux I__7844 (
            .O(N__47171),
            .I(throttle_order_7));
    Odrv4 I__7843 (
            .O(N__47168),
            .I(throttle_order_7));
    InMux I__7842 (
            .O(N__47163),
            .I(N__47160));
    LocalMux I__7841 (
            .O(N__47160),
            .I(N__47155));
    InMux I__7840 (
            .O(N__47159),
            .I(N__47152));
    InMux I__7839 (
            .O(N__47158),
            .I(N__47149));
    Span4Mux_v I__7838 (
            .O(N__47155),
            .I(N__47146));
    LocalMux I__7837 (
            .O(N__47152),
            .I(\ppm_encoder_1.elevatorZ0Z_8 ));
    LocalMux I__7836 (
            .O(N__47149),
            .I(\ppm_encoder_1.elevatorZ0Z_8 ));
    Odrv4 I__7835 (
            .O(N__47146),
            .I(\ppm_encoder_1.elevatorZ0Z_8 ));
    CascadeMux I__7834 (
            .O(N__47139),
            .I(N__47136));
    InMux I__7833 (
            .O(N__47136),
            .I(N__47132));
    InMux I__7832 (
            .O(N__47135),
            .I(N__47129));
    LocalMux I__7831 (
            .O(N__47132),
            .I(\ppm_encoder_1.N_265_i_i ));
    LocalMux I__7830 (
            .O(N__47129),
            .I(\ppm_encoder_1.N_265_i_i ));
    CascadeMux I__7829 (
            .O(N__47124),
            .I(N__47121));
    InMux I__7828 (
            .O(N__47121),
            .I(N__47118));
    LocalMux I__7827 (
            .O(N__47118),
            .I(N__47113));
    InMux I__7826 (
            .O(N__47117),
            .I(N__47108));
    InMux I__7825 (
            .O(N__47116),
            .I(N__47108));
    Span4Mux_h I__7824 (
            .O(N__47113),
            .I(N__47105));
    LocalMux I__7823 (
            .O(N__47108),
            .I(\ppm_encoder_1.throttleZ0Z_9 ));
    Odrv4 I__7822 (
            .O(N__47105),
            .I(\ppm_encoder_1.throttleZ0Z_9 ));
    InMux I__7821 (
            .O(N__47100),
            .I(N__47097));
    LocalMux I__7820 (
            .O(N__47097),
            .I(\ppm_encoder_1.un2_throttle_iv_0_1_9 ));
    InMux I__7819 (
            .O(N__47094),
            .I(N__47089));
    InMux I__7818 (
            .O(N__47093),
            .I(N__47084));
    InMux I__7817 (
            .O(N__47092),
            .I(N__47084));
    LocalMux I__7816 (
            .O(N__47089),
            .I(N__47081));
    LocalMux I__7815 (
            .O(N__47084),
            .I(\ppm_encoder_1.elevatorZ0Z_4 ));
    Odrv4 I__7814 (
            .O(N__47081),
            .I(\ppm_encoder_1.elevatorZ0Z_4 ));
    CascadeMux I__7813 (
            .O(N__47076),
            .I(\ppm_encoder_1.rudder_RNIM1KQZ0Z_12_cascade_ ));
    CascadeMux I__7812 (
            .O(N__47073),
            .I(\ppm_encoder_1.un2_throttle_iv_0_2_12_cascade_ ));
    CascadeMux I__7811 (
            .O(N__47070),
            .I(N__47067));
    InMux I__7810 (
            .O(N__47067),
            .I(N__47064));
    LocalMux I__7809 (
            .O(N__47064),
            .I(\ppm_encoder_1.un1_init_pulses_10_16 ));
    InMux I__7808 (
            .O(N__47061),
            .I(N__47058));
    LocalMux I__7807 (
            .O(N__47058),
            .I(\ppm_encoder_1.un1_init_pulses_11_16 ));
    InMux I__7806 (
            .O(N__47055),
            .I(N__47052));
    LocalMux I__7805 (
            .O(N__47052),
            .I(\ppm_encoder_1.un1_init_pulses_11_17 ));
    InMux I__7804 (
            .O(N__47049),
            .I(N__47046));
    LocalMux I__7803 (
            .O(N__47046),
            .I(\ppm_encoder_1.un1_init_pulses_10_17 ));
    InMux I__7802 (
            .O(N__47043),
            .I(N__47040));
    LocalMux I__7801 (
            .O(N__47040),
            .I(\ppm_encoder_1.un1_init_pulses_11_18 ));
    InMux I__7800 (
            .O(N__47037),
            .I(N__47034));
    LocalMux I__7799 (
            .O(N__47034),
            .I(\ppm_encoder_1.un1_init_pulses_10_18 ));
    InMux I__7798 (
            .O(N__47031),
            .I(N__47028));
    LocalMux I__7797 (
            .O(N__47028),
            .I(\ppm_encoder_1.un1_init_pulses_10_1 ));
    InMux I__7796 (
            .O(N__47025),
            .I(N__47022));
    LocalMux I__7795 (
            .O(N__47022),
            .I(N__47019));
    Odrv12 I__7794 (
            .O(N__47019),
            .I(\ppm_encoder_1.un1_init_pulses_11_1 ));
    CascadeMux I__7793 (
            .O(N__47016),
            .I(N__47013));
    InMux I__7792 (
            .O(N__47013),
            .I(N__47010));
    LocalMux I__7791 (
            .O(N__47010),
            .I(N__47007));
    Odrv4 I__7790 (
            .O(N__47007),
            .I(\ppm_encoder_1.un1_init_pulses_10_10 ));
    InMux I__7789 (
            .O(N__47004),
            .I(N__47001));
    LocalMux I__7788 (
            .O(N__47001),
            .I(N__46998));
    Odrv4 I__7787 (
            .O(N__46998),
            .I(\ppm_encoder_1.un1_init_pulses_11_10 ));
    CascadeMux I__7786 (
            .O(N__46995),
            .I(N__46992));
    InMux I__7785 (
            .O(N__46992),
            .I(N__46989));
    LocalMux I__7784 (
            .O(N__46989),
            .I(N__46986));
    Span4Mux_v I__7783 (
            .O(N__46986),
            .I(N__46983));
    Odrv4 I__7782 (
            .O(N__46983),
            .I(\ppm_encoder_1.un1_init_pulses_11_9 ));
    InMux I__7781 (
            .O(N__46980),
            .I(N__46977));
    LocalMux I__7780 (
            .O(N__46977),
            .I(\ppm_encoder_1.un1_init_pulses_10_9 ));
    CascadeMux I__7779 (
            .O(N__46974),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_9_cascade_ ));
    InMux I__7778 (
            .O(N__46971),
            .I(N__46968));
    LocalMux I__7777 (
            .O(N__46968),
            .I(\ppm_encoder_1.init_pulses_RNIEBKU5Z0Z_9 ));
    InMux I__7776 (
            .O(N__46965),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_14 ));
    InMux I__7775 (
            .O(N__46962),
            .I(bfn_11_3_0_));
    InMux I__7774 (
            .O(N__46959),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_16 ));
    InMux I__7773 (
            .O(N__46956),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_17 ));
    InMux I__7772 (
            .O(N__46953),
            .I(N__46950));
    LocalMux I__7771 (
            .O(N__46950),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_15 ));
    InMux I__7770 (
            .O(N__46947),
            .I(N__46944));
    LocalMux I__7769 (
            .O(N__46944),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_16 ));
    CascadeMux I__7768 (
            .O(N__46941),
            .I(N__46938));
    InMux I__7767 (
            .O(N__46938),
            .I(N__46935));
    LocalMux I__7766 (
            .O(N__46935),
            .I(N__46932));
    Odrv4 I__7765 (
            .O(N__46932),
            .I(\ppm_encoder_1.un1_init_pulses_11_15 ));
    InMux I__7764 (
            .O(N__46929),
            .I(N__46926));
    LocalMux I__7763 (
            .O(N__46926),
            .I(\ppm_encoder_1.un1_init_pulses_10_15 ));
    InMux I__7762 (
            .O(N__46923),
            .I(N__46920));
    LocalMux I__7761 (
            .O(N__46920),
            .I(N__46917));
    Span4Mux_h I__7760 (
            .O(N__46917),
            .I(N__46914));
    Odrv4 I__7759 (
            .O(N__46914),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_7 ));
    InMux I__7758 (
            .O(N__46911),
            .I(N__46908));
    LocalMux I__7757 (
            .O(N__46908),
            .I(\ppm_encoder_1.un1_init_pulses_11_7 ));
    InMux I__7756 (
            .O(N__46905),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_6 ));
    InMux I__7755 (
            .O(N__46902),
            .I(N__46899));
    LocalMux I__7754 (
            .O(N__46899),
            .I(N__46896));
    Span4Mux_s2_v I__7753 (
            .O(N__46896),
            .I(N__46893));
    Odrv4 I__7752 (
            .O(N__46893),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_8 ));
    InMux I__7751 (
            .O(N__46890),
            .I(N__46887));
    LocalMux I__7750 (
            .O(N__46887),
            .I(\ppm_encoder_1.un1_init_pulses_11_8 ));
    InMux I__7749 (
            .O(N__46884),
            .I(bfn_11_2_0_));
    InMux I__7748 (
            .O(N__46881),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_8 ));
    InMux I__7747 (
            .O(N__46878),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_9 ));
    InMux I__7746 (
            .O(N__46875),
            .I(N__46872));
    LocalMux I__7745 (
            .O(N__46872),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_11 ));
    InMux I__7744 (
            .O(N__46869),
            .I(N__46866));
    LocalMux I__7743 (
            .O(N__46866),
            .I(\ppm_encoder_1.un1_init_pulses_11_11 ));
    InMux I__7742 (
            .O(N__46863),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_10 ));
    InMux I__7741 (
            .O(N__46860),
            .I(N__46857));
    LocalMux I__7740 (
            .O(N__46857),
            .I(\ppm_encoder_1.un1_init_pulses_11_12 ));
    InMux I__7739 (
            .O(N__46854),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_11 ));
    InMux I__7738 (
            .O(N__46851),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_12 ));
    InMux I__7737 (
            .O(N__46848),
            .I(N__46845));
    LocalMux I__7736 (
            .O(N__46845),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_14 ));
    InMux I__7735 (
            .O(N__46842),
            .I(N__46839));
    LocalMux I__7734 (
            .O(N__46839),
            .I(\ppm_encoder_1.un1_init_pulses_11_14 ));
    InMux I__7733 (
            .O(N__46836),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_13 ));
    IoInMux I__7732 (
            .O(N__46833),
            .I(N__46830));
    LocalMux I__7731 (
            .O(N__46830),
            .I(N__46827));
    Span4Mux_s0_v I__7730 (
            .O(N__46827),
            .I(N__46824));
    Span4Mux_h I__7729 (
            .O(N__46824),
            .I(N__46821));
    Odrv4 I__7728 (
            .O(N__46821),
            .I(\pid_front.state_RNIPKTDZ0Z_0 ));
    InMux I__7727 (
            .O(N__46818),
            .I(N__46815));
    LocalMux I__7726 (
            .O(N__46815),
            .I(\ppm_encoder_1.N_39_i ));
    InMux I__7725 (
            .O(N__46812),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_0 ));
    InMux I__7724 (
            .O(N__46809),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_1 ));
    InMux I__7723 (
            .O(N__46806),
            .I(N__46803));
    LocalMux I__7722 (
            .O(N__46803),
            .I(\ppm_encoder_1.un1_init_pulses_11_3 ));
    InMux I__7721 (
            .O(N__46800),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_2 ));
    InMux I__7720 (
            .O(N__46797),
            .I(N__46794));
    LocalMux I__7719 (
            .O(N__46794),
            .I(\ppm_encoder_1.un1_init_pulses_11_4 ));
    InMux I__7718 (
            .O(N__46791),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_3 ));
    InMux I__7717 (
            .O(N__46788),
            .I(N__46785));
    LocalMux I__7716 (
            .O(N__46785),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_5 ));
    InMux I__7715 (
            .O(N__46782),
            .I(N__46779));
    LocalMux I__7714 (
            .O(N__46779),
            .I(\ppm_encoder_1.un1_init_pulses_11_5 ));
    InMux I__7713 (
            .O(N__46776),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_4 ));
    InMux I__7712 (
            .O(N__46773),
            .I(N__46770));
    LocalMux I__7711 (
            .O(N__46770),
            .I(\ppm_encoder_1.un1_init_pulses_11_6 ));
    InMux I__7710 (
            .O(N__46767),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_5 ));
    CascadeMux I__7709 (
            .O(N__46764),
            .I(\pid_front.error_d_reg_prev_esr_RNI5JRF4_0Z0Z_10_cascade_ ));
    InMux I__7708 (
            .O(N__46761),
            .I(N__46758));
    LocalMux I__7707 (
            .O(N__46758),
            .I(N__46755));
    Span4Mux_v I__7706 (
            .O(N__46755),
            .I(N__46751));
    InMux I__7705 (
            .O(N__46754),
            .I(N__46748));
    Span4Mux_h I__7704 (
            .O(N__46751),
            .I(N__46743));
    LocalMux I__7703 (
            .O(N__46748),
            .I(N__46743));
    Span4Mux_v I__7702 (
            .O(N__46743),
            .I(N__46740));
    Odrv4 I__7701 (
            .O(N__46740),
            .I(\pid_front.error_d_reg_prev_esr_RNIO00C5_0Z0Z_10 ));
    InMux I__7700 (
            .O(N__46737),
            .I(N__46734));
    LocalMux I__7699 (
            .O(N__46734),
            .I(N__46731));
    Span4Mux_v I__7698 (
            .O(N__46731),
            .I(N__46728));
    Span4Mux_v I__7697 (
            .O(N__46728),
            .I(N__46724));
    InMux I__7696 (
            .O(N__46727),
            .I(N__46721));
    Odrv4 I__7695 (
            .O(N__46724),
            .I(\pid_front.error_d_reg_prev_esr_RNI5JRF4_0Z0Z_10 ));
    LocalMux I__7694 (
            .O(N__46721),
            .I(\pid_front.error_d_reg_prev_esr_RNI5JRF4_0Z0Z_10 ));
    CascadeMux I__7693 (
            .O(N__46716),
            .I(N__46713));
    InMux I__7692 (
            .O(N__46713),
            .I(N__46710));
    LocalMux I__7691 (
            .O(N__46710),
            .I(N__46707));
    Span4Mux_v I__7690 (
            .O(N__46707),
            .I(N__46704));
    Odrv4 I__7689 (
            .O(N__46704),
            .I(\pid_front.error_d_reg_prev_esr_RNIO00C5Z0Z_10 ));
    InMux I__7688 (
            .O(N__46701),
            .I(N__46698));
    LocalMux I__7687 (
            .O(N__46698),
            .I(N__46691));
    InMux I__7686 (
            .O(N__46697),
            .I(N__46682));
    InMux I__7685 (
            .O(N__46696),
            .I(N__46682));
    InMux I__7684 (
            .O(N__46695),
            .I(N__46682));
    InMux I__7683 (
            .O(N__46694),
            .I(N__46682));
    Odrv12 I__7682 (
            .O(N__46691),
            .I(\pid_front.error_d_regZ0Z_9 ));
    LocalMux I__7681 (
            .O(N__46682),
            .I(\pid_front.error_d_regZ0Z_9 ));
    InMux I__7680 (
            .O(N__46677),
            .I(N__46674));
    LocalMux I__7679 (
            .O(N__46674),
            .I(N__46669));
    CascadeMux I__7678 (
            .O(N__46673),
            .I(N__46666));
    CascadeMux I__7677 (
            .O(N__46672),
            .I(N__46663));
    Span4Mux_v I__7676 (
            .O(N__46669),
            .I(N__46659));
    InMux I__7675 (
            .O(N__46666),
            .I(N__46652));
    InMux I__7674 (
            .O(N__46663),
            .I(N__46652));
    InMux I__7673 (
            .O(N__46662),
            .I(N__46652));
    Odrv4 I__7672 (
            .O(N__46659),
            .I(\pid_front.error_d_reg_prevZ0Z_9 ));
    LocalMux I__7671 (
            .O(N__46652),
            .I(\pid_front.error_d_reg_prevZ0Z_9 ));
    CascadeMux I__7670 (
            .O(N__46647),
            .I(N__46644));
    InMux I__7669 (
            .O(N__46644),
            .I(N__46638));
    InMux I__7668 (
            .O(N__46643),
            .I(N__46638));
    LocalMux I__7667 (
            .O(N__46638),
            .I(N__46635));
    Span4Mux_v I__7666 (
            .O(N__46635),
            .I(N__46632));
    Odrv4 I__7665 (
            .O(N__46632),
            .I(\pid_front.N_2173_i ));
    InMux I__7664 (
            .O(N__46629),
            .I(N__46626));
    LocalMux I__7663 (
            .O(N__46626),
            .I(N__46623));
    Span4Mux_h I__7662 (
            .O(N__46623),
            .I(N__46620));
    Span4Mux_h I__7661 (
            .O(N__46620),
            .I(N__46617));
    Span4Mux_h I__7660 (
            .O(N__46617),
            .I(N__46614));
    Span4Mux_h I__7659 (
            .O(N__46614),
            .I(N__46611));
    Odrv4 I__7658 (
            .O(N__46611),
            .I(\pid_front.O_13 ));
    InMux I__7657 (
            .O(N__46608),
            .I(N__46605));
    LocalMux I__7656 (
            .O(N__46605),
            .I(N__46602));
    Span4Mux_h I__7655 (
            .O(N__46602),
            .I(N__46599));
    Span4Mux_h I__7654 (
            .O(N__46599),
            .I(N__46596));
    Span4Mux_h I__7653 (
            .O(N__46596),
            .I(N__46593));
    Span4Mux_h I__7652 (
            .O(N__46593),
            .I(N__46590));
    Odrv4 I__7651 (
            .O(N__46590),
            .I(\pid_front.O_11 ));
    InMux I__7650 (
            .O(N__46587),
            .I(N__46584));
    LocalMux I__7649 (
            .O(N__46584),
            .I(N__46578));
    InMux I__7648 (
            .O(N__46583),
            .I(N__46575));
    InMux I__7647 (
            .O(N__46582),
            .I(N__46570));
    InMux I__7646 (
            .O(N__46581),
            .I(N__46570));
    Odrv4 I__7645 (
            .O(N__46578),
            .I(\pid_front.error_d_reg_fastZ0Z_12 ));
    LocalMux I__7644 (
            .O(N__46575),
            .I(\pid_front.error_d_reg_fastZ0Z_12 ));
    LocalMux I__7643 (
            .O(N__46570),
            .I(\pid_front.error_d_reg_fastZ0Z_12 ));
    InMux I__7642 (
            .O(N__46563),
            .I(N__46560));
    LocalMux I__7641 (
            .O(N__46560),
            .I(N__46557));
    Span12Mux_v I__7640 (
            .O(N__46557),
            .I(N__46554));
    Span12Mux_h I__7639 (
            .O(N__46554),
            .I(N__46551));
    Odrv12 I__7638 (
            .O(N__46551),
            .I(\pid_front.O_15 ));
    CascadeMux I__7637 (
            .O(N__46548),
            .I(\pid_front.error_p_reg_esr_RNIKG5U_0Z0Z_10_cascade_ ));
    InMux I__7636 (
            .O(N__46545),
            .I(N__46542));
    LocalMux I__7635 (
            .O(N__46542),
            .I(\pid_front.error_p_reg_esr_RNIKG5UZ0Z_10 ));
    InMux I__7634 (
            .O(N__46539),
            .I(N__46536));
    LocalMux I__7633 (
            .O(N__46536),
            .I(\pid_front.error_d_reg_prev_esr_RNI379B2Z0Z_10 ));
    InMux I__7632 (
            .O(N__46533),
            .I(N__46528));
    InMux I__7631 (
            .O(N__46532),
            .I(N__46523));
    InMux I__7630 (
            .O(N__46531),
            .I(N__46523));
    LocalMux I__7629 (
            .O(N__46528),
            .I(N__46520));
    LocalMux I__7628 (
            .O(N__46523),
            .I(N__46516));
    Span4Mux_v I__7627 (
            .O(N__46520),
            .I(N__46513));
    InMux I__7626 (
            .O(N__46519),
            .I(N__46510));
    Span4Mux_v I__7625 (
            .O(N__46516),
            .I(N__46507));
    Odrv4 I__7624 (
            .O(N__46513),
            .I(\pid_front.error_d_reg_prevZ0Z_10 ));
    LocalMux I__7623 (
            .O(N__46510),
            .I(\pid_front.error_d_reg_prevZ0Z_10 ));
    Odrv4 I__7622 (
            .O(N__46507),
            .I(\pid_front.error_d_reg_prevZ0Z_10 ));
    CascadeMux I__7621 (
            .O(N__46500),
            .I(N__46497));
    InMux I__7620 (
            .O(N__46497),
            .I(N__46492));
    InMux I__7619 (
            .O(N__46496),
            .I(N__46487));
    InMux I__7618 (
            .O(N__46495),
            .I(N__46487));
    LocalMux I__7617 (
            .O(N__46492),
            .I(N__46481));
    LocalMux I__7616 (
            .O(N__46487),
            .I(N__46478));
    InMux I__7615 (
            .O(N__46486),
            .I(N__46471));
    InMux I__7614 (
            .O(N__46485),
            .I(N__46471));
    InMux I__7613 (
            .O(N__46484),
            .I(N__46471));
    Odrv4 I__7612 (
            .O(N__46481),
            .I(\pid_front.error_d_regZ0Z_10 ));
    Odrv12 I__7611 (
            .O(N__46478),
            .I(\pid_front.error_d_regZ0Z_10 ));
    LocalMux I__7610 (
            .O(N__46471),
            .I(\pid_front.error_d_regZ0Z_10 ));
    CascadeMux I__7609 (
            .O(N__46464),
            .I(\pid_front.error_d_reg_prev_esr_RNI379B2Z0Z_10_cascade_ ));
    InMux I__7608 (
            .O(N__46461),
            .I(N__46457));
    InMux I__7607 (
            .O(N__46460),
            .I(N__46454));
    LocalMux I__7606 (
            .O(N__46457),
            .I(N__46451));
    LocalMux I__7605 (
            .O(N__46454),
            .I(\pid_front.error_p_reg_esr_RNI8NB61_1Z0Z_11 ));
    Odrv4 I__7604 (
            .O(N__46451),
            .I(\pid_front.error_p_reg_esr_RNI8NB61_1Z0Z_11 ));
    CascadeMux I__7603 (
            .O(N__46446),
            .I(\pid_front.error_d_reg_fast_esr_RNID6KB1Z0Z_12_cascade_ ));
    CascadeMux I__7602 (
            .O(N__46443),
            .I(\pid_front.error_d_reg_fast_esr_RNIQSG63Z0Z_12_cascade_ ));
    InMux I__7601 (
            .O(N__46440),
            .I(N__46437));
    LocalMux I__7600 (
            .O(N__46437),
            .I(\pid_front.error_p_reg_esr_RNIETB61_1Z0Z_13 ));
    CascadeMux I__7599 (
            .O(N__46434),
            .I(\pid_front.un1_pid_prereg_97_cascade_ ));
    InMux I__7598 (
            .O(N__46431),
            .I(N__46428));
    LocalMux I__7597 (
            .O(N__46428),
            .I(N__46425));
    Odrv4 I__7596 (
            .O(N__46425),
            .I(\pid_front.un1_pid_prereg_167_0 ));
    InMux I__7595 (
            .O(N__46422),
            .I(N__46419));
    LocalMux I__7594 (
            .O(N__46419),
            .I(N__46416));
    Span4Mux_v I__7593 (
            .O(N__46416),
            .I(N__46412));
    InMux I__7592 (
            .O(N__46415),
            .I(N__46409));
    Odrv4 I__7591 (
            .O(N__46412),
            .I(\pid_front.error_p_reg_esr_RNI8C7GBZ0Z_13 ));
    LocalMux I__7590 (
            .O(N__46409),
            .I(\pid_front.error_p_reg_esr_RNI8C7GBZ0Z_13 ));
    InMux I__7589 (
            .O(N__46404),
            .I(N__46401));
    LocalMux I__7588 (
            .O(N__46401),
            .I(N__46397));
    InMux I__7587 (
            .O(N__46400),
            .I(N__46394));
    Odrv4 I__7586 (
            .O(N__46397),
            .I(\pid_front.error_p_reg_esr_RNIT79QCZ0Z_12 ));
    LocalMux I__7585 (
            .O(N__46394),
            .I(\pid_front.error_p_reg_esr_RNIT79QCZ0Z_12 ));
    CascadeMux I__7584 (
            .O(N__46389),
            .I(\pid_front.error_p_reg_esr_RNI8C7GBZ0Z_13_cascade_ ));
    CascadeMux I__7583 (
            .O(N__46386),
            .I(N__46383));
    InMux I__7582 (
            .O(N__46383),
            .I(N__46380));
    LocalMux I__7581 (
            .O(N__46380),
            .I(N__46375));
    InMux I__7580 (
            .O(N__46379),
            .I(N__46372));
    InMux I__7579 (
            .O(N__46378),
            .I(N__46369));
    Odrv12 I__7578 (
            .O(N__46375),
            .I(\pid_front.error_p_reg_esr_RNIBJ5B3_0Z0Z_14 ));
    LocalMux I__7577 (
            .O(N__46372),
            .I(\pid_front.error_p_reg_esr_RNIBJ5B3_0Z0Z_14 ));
    LocalMux I__7576 (
            .O(N__46369),
            .I(\pid_front.error_p_reg_esr_RNIBJ5B3_0Z0Z_14 ));
    CascadeMux I__7575 (
            .O(N__46362),
            .I(N__46359));
    InMux I__7574 (
            .O(N__46359),
            .I(N__46356));
    LocalMux I__7573 (
            .O(N__46356),
            .I(N__46353));
    Odrv4 I__7572 (
            .O(N__46353),
            .I(\pid_front.error_p_reg_esr_RNIG7MLRZ0Z_12 ));
    InMux I__7571 (
            .O(N__46350),
            .I(N__46347));
    LocalMux I__7570 (
            .O(N__46347),
            .I(\pid_front.error_d_reg_fast_esr_RNI5VGKZ0Z_12 ));
    CascadeMux I__7569 (
            .O(N__46344),
            .I(N__46341));
    InMux I__7568 (
            .O(N__46341),
            .I(N__46328));
    InMux I__7567 (
            .O(N__46340),
            .I(N__46323));
    InMux I__7566 (
            .O(N__46339),
            .I(N__46323));
    CascadeMux I__7565 (
            .O(N__46338),
            .I(N__46319));
    CascadeMux I__7564 (
            .O(N__46337),
            .I(N__46316));
    CascadeMux I__7563 (
            .O(N__46336),
            .I(N__46313));
    CascadeMux I__7562 (
            .O(N__46335),
            .I(N__46309));
    CascadeMux I__7561 (
            .O(N__46334),
            .I(N__46306));
    CascadeMux I__7560 (
            .O(N__46333),
            .I(N__46303));
    CascadeMux I__7559 (
            .O(N__46332),
            .I(N__46300));
    CascadeMux I__7558 (
            .O(N__46331),
            .I(N__46297));
    LocalMux I__7557 (
            .O(N__46328),
            .I(N__46294));
    LocalMux I__7556 (
            .O(N__46323),
            .I(N__46291));
    InMux I__7555 (
            .O(N__46322),
            .I(N__46282));
    InMux I__7554 (
            .O(N__46319),
            .I(N__46282));
    InMux I__7553 (
            .O(N__46316),
            .I(N__46282));
    InMux I__7552 (
            .O(N__46313),
            .I(N__46282));
    InMux I__7551 (
            .O(N__46312),
            .I(N__46275));
    InMux I__7550 (
            .O(N__46309),
            .I(N__46275));
    InMux I__7549 (
            .O(N__46306),
            .I(N__46275));
    InMux I__7548 (
            .O(N__46303),
            .I(N__46268));
    InMux I__7547 (
            .O(N__46300),
            .I(N__46268));
    InMux I__7546 (
            .O(N__46297),
            .I(N__46268));
    Span4Mux_v I__7545 (
            .O(N__46294),
            .I(N__46265));
    Span4Mux_h I__7544 (
            .O(N__46291),
            .I(N__46262));
    LocalMux I__7543 (
            .O(N__46282),
            .I(\pid_front.error_d_reg_prevZ0Z_22 ));
    LocalMux I__7542 (
            .O(N__46275),
            .I(\pid_front.error_d_reg_prevZ0Z_22 ));
    LocalMux I__7541 (
            .O(N__46268),
            .I(\pid_front.error_d_reg_prevZ0Z_22 ));
    Odrv4 I__7540 (
            .O(N__46265),
            .I(\pid_front.error_d_reg_prevZ0Z_22 ));
    Odrv4 I__7539 (
            .O(N__46262),
            .I(\pid_front.error_d_reg_prevZ0Z_22 ));
    InMux I__7538 (
            .O(N__46251),
            .I(N__46242));
    InMux I__7537 (
            .O(N__46250),
            .I(N__46242));
    InMux I__7536 (
            .O(N__46249),
            .I(N__46242));
    LocalMux I__7535 (
            .O(N__46242),
            .I(\pid_front.un1_pid_prereg_0_16 ));
    InMux I__7534 (
            .O(N__46239),
            .I(N__46236));
    LocalMux I__7533 (
            .O(N__46236),
            .I(N__46233));
    Span4Mux_h I__7532 (
            .O(N__46233),
            .I(N__46230));
    Span4Mux_h I__7531 (
            .O(N__46230),
            .I(N__46227));
    Span4Mux_h I__7530 (
            .O(N__46227),
            .I(N__46224));
    Span4Mux_h I__7529 (
            .O(N__46224),
            .I(N__46221));
    Odrv4 I__7528 (
            .O(N__46221),
            .I(\pid_front.O_12 ));
    CascadeMux I__7527 (
            .O(N__46218),
            .I(\pid_front.g0_1_cascade_ ));
    InMux I__7526 (
            .O(N__46215),
            .I(N__46212));
    LocalMux I__7525 (
            .O(N__46212),
            .I(\pid_front.g0_2_0 ));
    CascadeMux I__7524 (
            .O(N__46209),
            .I(\pid_front.error_p_reg_esr_RNIU52U6Z0Z_12_cascade_ ));
    InMux I__7523 (
            .O(N__46206),
            .I(N__46203));
    LocalMux I__7522 (
            .O(N__46203),
            .I(\pid_front.g1_3 ));
    InMux I__7521 (
            .O(N__46200),
            .I(N__46197));
    LocalMux I__7520 (
            .O(N__46197),
            .I(N__46194));
    Odrv4 I__7519 (
            .O(N__46194),
            .I(\pid_front.g1_2_1 ));
    InMux I__7518 (
            .O(N__46191),
            .I(N__46188));
    LocalMux I__7517 (
            .O(N__46188),
            .I(N__46185));
    Span4Mux_h I__7516 (
            .O(N__46185),
            .I(N__46182));
    Odrv4 I__7515 (
            .O(N__46182),
            .I(\pid_front.error_p_reg_esr_RNICU3D1_0Z0Z_6 ));
    CascadeMux I__7514 (
            .O(N__46179),
            .I(N__46176));
    InMux I__7513 (
            .O(N__46176),
            .I(N__46170));
    InMux I__7512 (
            .O(N__46175),
            .I(N__46170));
    LocalMux I__7511 (
            .O(N__46170),
            .I(N__46167));
    Span4Mux_v I__7510 (
            .O(N__46167),
            .I(N__46164));
    Odrv4 I__7509 (
            .O(N__46164),
            .I(\pid_front.error_p_reg_esr_RNI6B6FZ0Z_6 ));
    InMux I__7508 (
            .O(N__46161),
            .I(N__46158));
    LocalMux I__7507 (
            .O(N__46158),
            .I(\pid_front.N_2198_0_0_0 ));
    CascadeMux I__7506 (
            .O(N__46155),
            .I(N__46152));
    InMux I__7505 (
            .O(N__46152),
            .I(N__46149));
    LocalMux I__7504 (
            .O(N__46149),
            .I(N__46145));
    InMux I__7503 (
            .O(N__46148),
            .I(N__46142));
    Odrv4 I__7502 (
            .O(N__46145),
            .I(\pid_front.un1_pid_prereg_0_15 ));
    LocalMux I__7501 (
            .O(N__46142),
            .I(\pid_front.un1_pid_prereg_0_15 ));
    InMux I__7500 (
            .O(N__46137),
            .I(N__46134));
    LocalMux I__7499 (
            .O(N__46134),
            .I(\pid_front.error_d_reg_prev_esr_RNIOS1BCZ0Z_22 ));
    InMux I__7498 (
            .O(N__46131),
            .I(N__46128));
    LocalMux I__7497 (
            .O(N__46128),
            .I(\pid_front.un1_pid_prereg_370_1 ));
    CascadeMux I__7496 (
            .O(N__46125),
            .I(\pid_front.un1_pid_prereg_370_1_cascade_ ));
    InMux I__7495 (
            .O(N__46122),
            .I(N__46116));
    InMux I__7494 (
            .O(N__46121),
            .I(N__46116));
    LocalMux I__7493 (
            .O(N__46116),
            .I(\pid_front.un1_pid_prereg_0_13 ));
    CascadeMux I__7492 (
            .O(N__46113),
            .I(\pid_front.un1_pid_prereg_0_13_cascade_ ));
    CascadeMux I__7491 (
            .O(N__46110),
            .I(N__46107));
    InMux I__7490 (
            .O(N__46107),
            .I(N__46104));
    LocalMux I__7489 (
            .O(N__46104),
            .I(\pid_front.error_p_reg_esr_RNID7NO6Z0Z_20 ));
    CascadeMux I__7488 (
            .O(N__46101),
            .I(\pid_front.g1_1_cascade_ ));
    CascadeMux I__7487 (
            .O(N__46098),
            .I(\pid_front.g0_3_2_cascade_ ));
    CascadeMux I__7486 (
            .O(N__46095),
            .I(N__46092));
    InMux I__7485 (
            .O(N__46092),
            .I(N__46089));
    LocalMux I__7484 (
            .O(N__46089),
            .I(N__46086));
    Span4Mux_v I__7483 (
            .O(N__46086),
            .I(N__46083));
    Odrv4 I__7482 (
            .O(N__46083),
            .I(\pid_front.g0_1_0_1 ));
    InMux I__7481 (
            .O(N__46080),
            .I(N__46077));
    LocalMux I__7480 (
            .O(N__46077),
            .I(\pid_front.N_4_1_1_1 ));
    InMux I__7479 (
            .O(N__46074),
            .I(N__46071));
    LocalMux I__7478 (
            .O(N__46071),
            .I(\pid_front.error_p_reg_esr_RNIFM3D1Z0Z_10 ));
    CascadeMux I__7477 (
            .O(N__46068),
            .I(\pid_front.error_p_reg_esr_RNILQ6FZ0Z_9_cascade_ ));
    CascadeMux I__7476 (
            .O(N__46065),
            .I(N__46062));
    InMux I__7475 (
            .O(N__46062),
            .I(N__46059));
    LocalMux I__7474 (
            .O(N__46059),
            .I(\pid_front.error_p_reg_esr_RNIEB5T7Z0Z_9 ));
    CascadeMux I__7473 (
            .O(N__46056),
            .I(N__46052));
    InMux I__7472 (
            .O(N__46055),
            .I(N__46047));
    InMux I__7471 (
            .O(N__46052),
            .I(N__46047));
    LocalMux I__7470 (
            .O(N__46047),
            .I(N__46044));
    Span4Mux_h I__7469 (
            .O(N__46044),
            .I(N__46041));
    Span4Mux_h I__7468 (
            .O(N__46041),
            .I(N__46038));
    Odrv4 I__7467 (
            .O(N__46038),
            .I(\pid_front.error_p_regZ0Z_9 ));
    InMux I__7466 (
            .O(N__46035),
            .I(N__46032));
    LocalMux I__7465 (
            .O(N__46032),
            .I(N__46029));
    Odrv4 I__7464 (
            .O(N__46029),
            .I(\pid_front.error_p_reg_esr_RNILQ6F_0Z0Z_9 ));
    CascadeMux I__7463 (
            .O(N__46026),
            .I(\pid_front.error_p_reg_esr_RNILQ6F_0Z0Z_9_cascade_ ));
    CascadeMux I__7462 (
            .O(N__46023),
            .I(N__46019));
    InMux I__7461 (
            .O(N__46022),
            .I(N__46016));
    InMux I__7460 (
            .O(N__46019),
            .I(N__46013));
    LocalMux I__7459 (
            .O(N__46016),
            .I(\pid_front.error_p_reg_esr_RNI6R6D1Z0Z_8 ));
    LocalMux I__7458 (
            .O(N__46013),
            .I(\pid_front.error_p_reg_esr_RNI6R6D1Z0Z_8 ));
    CascadeMux I__7457 (
            .O(N__46008),
            .I(\pid_front.un1_pid_prereg_0_15_cascade_ ));
    CascadeMux I__7456 (
            .O(N__46005),
            .I(N__46002));
    InMux I__7455 (
            .O(N__46002),
            .I(N__45999));
    LocalMux I__7454 (
            .O(N__45999),
            .I(\pid_front.error_d_reg_prev_esr_RNIBLAI5Z0Z_22 ));
    InMux I__7453 (
            .O(N__45996),
            .I(N__45993));
    LocalMux I__7452 (
            .O(N__45993),
            .I(N__45989));
    InMux I__7451 (
            .O(N__45992),
            .I(N__45986));
    Odrv12 I__7450 (
            .O(N__45989),
            .I(\pid_front.un1_pid_prereg_0_10 ));
    LocalMux I__7449 (
            .O(N__45986),
            .I(\pid_front.un1_pid_prereg_0_10 ));
    CascadeMux I__7448 (
            .O(N__45981),
            .I(N__45978));
    InMux I__7447 (
            .O(N__45978),
            .I(N__45975));
    LocalMux I__7446 (
            .O(N__45975),
            .I(N__45970));
    InMux I__7445 (
            .O(N__45974),
            .I(N__45965));
    InMux I__7444 (
            .O(N__45973),
            .I(N__45965));
    Odrv4 I__7443 (
            .O(N__45970),
            .I(\pid_front.un1_pid_prereg_0_11 ));
    LocalMux I__7442 (
            .O(N__45965),
            .I(\pid_front.un1_pid_prereg_0_11 ));
    InMux I__7441 (
            .O(N__45960),
            .I(N__45957));
    LocalMux I__7440 (
            .O(N__45957),
            .I(\pid_front.error_p_reg_esr_RNIF7HGDZ0Z_19 ));
    InMux I__7439 (
            .O(N__45954),
            .I(N__45951));
    LocalMux I__7438 (
            .O(N__45951),
            .I(N__45948));
    Span4Mux_v I__7437 (
            .O(N__45948),
            .I(N__45944));
    InMux I__7436 (
            .O(N__45947),
            .I(N__45941));
    Odrv4 I__7435 (
            .O(N__45944),
            .I(\pid_front.un1_pid_prereg_0_14 ));
    LocalMux I__7434 (
            .O(N__45941),
            .I(\pid_front.un1_pid_prereg_0_14 ));
    CascadeMux I__7433 (
            .O(N__45936),
            .I(\pid_front.un1_pid_prereg_0_14_cascade_ ));
    InMux I__7432 (
            .O(N__45933),
            .I(N__45930));
    LocalMux I__7431 (
            .O(N__45930),
            .I(\pid_front.error_p_reg_esr_RNI6B6F_0Z0Z_6 ));
    CascadeMux I__7430 (
            .O(N__45927),
            .I(N__45924));
    InMux I__7429 (
            .O(N__45924),
            .I(N__45921));
    LocalMux I__7428 (
            .O(N__45921),
            .I(\pid_front.error_p_reg_esr_RNIT2PE1Z0Z_5 ));
    CascadeMux I__7427 (
            .O(N__45918),
            .I(N__45915));
    InMux I__7426 (
            .O(N__45915),
            .I(N__45911));
    InMux I__7425 (
            .O(N__45914),
            .I(N__45908));
    LocalMux I__7424 (
            .O(N__45911),
            .I(N__45905));
    LocalMux I__7423 (
            .O(N__45908),
            .I(N__45902));
    Span4Mux_h I__7422 (
            .O(N__45905),
            .I(N__45899));
    Span4Mux_h I__7421 (
            .O(N__45902),
            .I(N__45896));
    Span4Mux_h I__7420 (
            .O(N__45899),
            .I(N__45893));
    Span4Mux_h I__7419 (
            .O(N__45896),
            .I(N__45890));
    Span4Mux_h I__7418 (
            .O(N__45893),
            .I(N__45887));
    Span4Mux_h I__7417 (
            .O(N__45890),
            .I(N__45884));
    Odrv4 I__7416 (
            .O(N__45887),
            .I(\pid_front.error_p_regZ0Z_5 ));
    Odrv4 I__7415 (
            .O(N__45884),
            .I(\pid_front.error_p_regZ0Z_5 ));
    InMux I__7414 (
            .O(N__45879),
            .I(N__45876));
    LocalMux I__7413 (
            .O(N__45876),
            .I(\pid_front.error_p_reg_esr_RNIUAE8Z0Z_4 ));
    InMux I__7412 (
            .O(N__45873),
            .I(N__45867));
    InMux I__7411 (
            .O(N__45872),
            .I(N__45867));
    LocalMux I__7410 (
            .O(N__45867),
            .I(\pid_front.error_p_reg_esr_RNIVOSGZ0Z_5 ));
    InMux I__7409 (
            .O(N__45864),
            .I(N__45861));
    LocalMux I__7408 (
            .O(N__45861),
            .I(\pid_front.N_2155_i ));
    CascadeMux I__7407 (
            .O(N__45858),
            .I(\pid_front.N_2155_i_cascade_ ));
    CascadeMux I__7406 (
            .O(N__45855),
            .I(N__45852));
    InMux I__7405 (
            .O(N__45852),
            .I(N__45848));
    InMux I__7404 (
            .O(N__45851),
            .I(N__45845));
    LocalMux I__7403 (
            .O(N__45848),
            .I(N__45840));
    LocalMux I__7402 (
            .O(N__45845),
            .I(N__45840));
    Span4Mux_v I__7401 (
            .O(N__45840),
            .I(N__45837));
    Sp12to4 I__7400 (
            .O(N__45837),
            .I(N__45834));
    Odrv12 I__7399 (
            .O(N__45834),
            .I(\pid_front.error_p_regZ0Z_6 ));
    CascadeMux I__7398 (
            .O(N__45831),
            .I(\pid_front.N_2179_i_cascade_ ));
    CascadeMux I__7397 (
            .O(N__45828),
            .I(\pid_front.error_p_reg_esr_RNIFM3D1Z0Z_10_cascade_ ));
    InMux I__7396 (
            .O(N__45825),
            .I(N__45822));
    LocalMux I__7395 (
            .O(N__45822),
            .I(\pid_front.error_p_reg_esr_RNIS5CU3Z0Z_9 ));
    InMux I__7394 (
            .O(N__45819),
            .I(N__45816));
    LocalMux I__7393 (
            .O(N__45816),
            .I(\pid_front.error_p_reg_esr_RNILQ6FZ0Z_9 ));
    CascadeMux I__7392 (
            .O(N__45813),
            .I(\pid_front.error_p_reg_esr_RNIUAE8_0Z0Z_4_cascade_ ));
    CascadeMux I__7391 (
            .O(N__45810),
            .I(N__45807));
    InMux I__7390 (
            .O(N__45807),
            .I(N__45804));
    LocalMux I__7389 (
            .O(N__45804),
            .I(\pid_front.error_p_reg_esr_RNIMI772Z0Z_3 ));
    InMux I__7388 (
            .O(N__45801),
            .I(N__45797));
    InMux I__7387 (
            .O(N__45800),
            .I(N__45794));
    LocalMux I__7386 (
            .O(N__45797),
            .I(\pid_front.error_p_reg_esr_RNIB9N71_0Z0Z_5 ));
    LocalMux I__7385 (
            .O(N__45794),
            .I(\pid_front.error_p_reg_esr_RNIB9N71_0Z0Z_5 ));
    InMux I__7384 (
            .O(N__45789),
            .I(N__45783));
    InMux I__7383 (
            .O(N__45788),
            .I(N__45783));
    LocalMux I__7382 (
            .O(N__45783),
            .I(N__45780));
    Span4Mux_v I__7381 (
            .O(N__45780),
            .I(N__45777));
    Sp12to4 I__7380 (
            .O(N__45777),
            .I(N__45774));
    Odrv12 I__7379 (
            .O(N__45774),
            .I(\pid_front.error_p_regZ0Z_4 ));
    InMux I__7378 (
            .O(N__45771),
            .I(N__45765));
    InMux I__7377 (
            .O(N__45770),
            .I(N__45765));
    LocalMux I__7376 (
            .O(N__45765),
            .I(\pid_front.error_d_reg_prevZ0Z_4 ));
    CascadeMux I__7375 (
            .O(N__45762),
            .I(\pid_front.error_p_reg_esr_RNIUAE8Z0Z_4_cascade_ ));
    CascadeMux I__7374 (
            .O(N__45759),
            .I(\pid_front.error_p_reg_esr_RNIVOSG_0Z0Z_5_cascade_ ));
    CascadeMux I__7373 (
            .O(N__45756),
            .I(N__45753));
    InMux I__7372 (
            .O(N__45753),
            .I(N__45750));
    LocalMux I__7371 (
            .O(N__45750),
            .I(\pid_front.error_p_reg_esr_RNIB9N71Z0Z_5 ));
    CascadeMux I__7370 (
            .O(N__45747),
            .I(\pid_front.error_p_reg_esr_RNI6B6F_0Z0Z_6_cascade_ ));
    InMux I__7369 (
            .O(N__45744),
            .I(N__45740));
    InMux I__7368 (
            .O(N__45743),
            .I(N__45737));
    LocalMux I__7367 (
            .O(N__45740),
            .I(\pid_front.error_p_reg_esr_RNIVOSG_0Z0Z_5 ));
    LocalMux I__7366 (
            .O(N__45737),
            .I(\pid_front.error_p_reg_esr_RNIVOSG_0Z0Z_5 ));
    CascadeMux I__7365 (
            .O(N__45732),
            .I(\pid_front.un1_pid_prereg_66_0_cascade_ ));
    InMux I__7364 (
            .O(N__45729),
            .I(N__45726));
    LocalMux I__7363 (
            .O(N__45726),
            .I(\pid_front.error_p_reg_esr_RNI8CGM2Z0Z_5 ));
    InMux I__7362 (
            .O(N__45723),
            .I(\ppm_encoder_1.un1_elevator_cry_13 ));
    InMux I__7361 (
            .O(N__45720),
            .I(N__45717));
    LocalMux I__7360 (
            .O(N__45717),
            .I(N__45714));
    Span4Mux_h I__7359 (
            .O(N__45714),
            .I(N__45710));
    InMux I__7358 (
            .O(N__45713),
            .I(N__45707));
    Odrv4 I__7357 (
            .O(N__45710),
            .I(front_order_13));
    LocalMux I__7356 (
            .O(N__45707),
            .I(front_order_13));
    InMux I__7355 (
            .O(N__45702),
            .I(N__45699));
    LocalMux I__7354 (
            .O(N__45699),
            .I(N__45694));
    InMux I__7353 (
            .O(N__45698),
            .I(N__45691));
    InMux I__7352 (
            .O(N__45697),
            .I(N__45687));
    Span4Mux_h I__7351 (
            .O(N__45694),
            .I(N__45684));
    LocalMux I__7350 (
            .O(N__45691),
            .I(N__45681));
    InMux I__7349 (
            .O(N__45690),
            .I(N__45678));
    LocalMux I__7348 (
            .O(N__45687),
            .I(N__45675));
    Span4Mux_v I__7347 (
            .O(N__45684),
            .I(N__45672));
    Span4Mux_h I__7346 (
            .O(N__45681),
            .I(N__45667));
    LocalMux I__7345 (
            .O(N__45678),
            .I(N__45667));
    Span4Mux_v I__7344 (
            .O(N__45675),
            .I(N__45664));
    Odrv4 I__7343 (
            .O(N__45672),
            .I(\pid_front.N_98 ));
    Odrv4 I__7342 (
            .O(N__45667),
            .I(\pid_front.N_98 ));
    Odrv4 I__7341 (
            .O(N__45664),
            .I(\pid_front.N_98 ));
    InMux I__7340 (
            .O(N__45657),
            .I(N__45650));
    InMux I__7339 (
            .O(N__45656),
            .I(N__45647));
    InMux I__7338 (
            .O(N__45655),
            .I(N__45644));
    InMux I__7337 (
            .O(N__45654),
            .I(N__45639));
    InMux I__7336 (
            .O(N__45653),
            .I(N__45639));
    LocalMux I__7335 (
            .O(N__45650),
            .I(N__45633));
    LocalMux I__7334 (
            .O(N__45647),
            .I(N__45633));
    LocalMux I__7333 (
            .O(N__45644),
            .I(N__45628));
    LocalMux I__7332 (
            .O(N__45639),
            .I(N__45628));
    CascadeMux I__7331 (
            .O(N__45638),
            .I(N__45625));
    Span4Mux_v I__7330 (
            .O(N__45633),
            .I(N__45622));
    Span4Mux_h I__7329 (
            .O(N__45628),
            .I(N__45619));
    InMux I__7328 (
            .O(N__45625),
            .I(N__45616));
    Odrv4 I__7327 (
            .O(N__45622),
            .I(\pid_front.pid_preregZ0Z_13 ));
    Odrv4 I__7326 (
            .O(N__45619),
            .I(\pid_front.pid_preregZ0Z_13 ));
    LocalMux I__7325 (
            .O(N__45616),
            .I(\pid_front.pid_preregZ0Z_13 ));
    CascadeMux I__7324 (
            .O(N__45609),
            .I(N__45605));
    InMux I__7323 (
            .O(N__45608),
            .I(N__45602));
    InMux I__7322 (
            .O(N__45605),
            .I(N__45599));
    LocalMux I__7321 (
            .O(N__45602),
            .I(N__45595));
    LocalMux I__7320 (
            .O(N__45599),
            .I(N__45592));
    InMux I__7319 (
            .O(N__45598),
            .I(N__45589));
    Span4Mux_h I__7318 (
            .O(N__45595),
            .I(N__45584));
    Span4Mux_h I__7317 (
            .O(N__45592),
            .I(N__45579));
    LocalMux I__7316 (
            .O(N__45589),
            .I(N__45579));
    InMux I__7315 (
            .O(N__45588),
            .I(N__45574));
    InMux I__7314 (
            .O(N__45587),
            .I(N__45574));
    Odrv4 I__7313 (
            .O(N__45584),
            .I(\pid_front.pid_preregZ0Z_12 ));
    Odrv4 I__7312 (
            .O(N__45579),
            .I(\pid_front.pid_preregZ0Z_12 ));
    LocalMux I__7311 (
            .O(N__45574),
            .I(\pid_front.pid_preregZ0Z_12 ));
    InMux I__7310 (
            .O(N__45567),
            .I(N__45564));
    LocalMux I__7309 (
            .O(N__45564),
            .I(N__45560));
    InMux I__7308 (
            .O(N__45563),
            .I(N__45557));
    Span4Mux_v I__7307 (
            .O(N__45560),
            .I(N__45552));
    LocalMux I__7306 (
            .O(N__45557),
            .I(N__45552));
    Odrv4 I__7305 (
            .O(N__45552),
            .I(front_order_12));
    InMux I__7304 (
            .O(N__45549),
            .I(N__45545));
    InMux I__7303 (
            .O(N__45548),
            .I(N__45542));
    LocalMux I__7302 (
            .O(N__45545),
            .I(N__45539));
    LocalMux I__7301 (
            .O(N__45542),
            .I(N__45536));
    Span4Mux_h I__7300 (
            .O(N__45539),
            .I(N__45532));
    Span4Mux_h I__7299 (
            .O(N__45536),
            .I(N__45529));
    InMux I__7298 (
            .O(N__45535),
            .I(N__45526));
    Odrv4 I__7297 (
            .O(N__45532),
            .I(\pid_front.pid_preregZ0Z_8 ));
    Odrv4 I__7296 (
            .O(N__45529),
            .I(\pid_front.pid_preregZ0Z_8 ));
    LocalMux I__7295 (
            .O(N__45526),
            .I(\pid_front.pid_preregZ0Z_8 ));
    InMux I__7294 (
            .O(N__45519),
            .I(N__45515));
    InMux I__7293 (
            .O(N__45518),
            .I(N__45512));
    LocalMux I__7292 (
            .O(N__45515),
            .I(N__45509));
    LocalMux I__7291 (
            .O(N__45512),
            .I(N__45506));
    Odrv12 I__7290 (
            .O(N__45509),
            .I(front_order_8));
    Odrv4 I__7289 (
            .O(N__45506),
            .I(front_order_8));
    InMux I__7288 (
            .O(N__45501),
            .I(N__45496));
    CascadeMux I__7287 (
            .O(N__45500),
            .I(N__45493));
    CascadeMux I__7286 (
            .O(N__45499),
            .I(N__45490));
    LocalMux I__7285 (
            .O(N__45496),
            .I(N__45487));
    InMux I__7284 (
            .O(N__45493),
            .I(N__45482));
    InMux I__7283 (
            .O(N__45490),
            .I(N__45482));
    Odrv4 I__7282 (
            .O(N__45487),
            .I(\pid_front.pid_preregZ0Z_11 ));
    LocalMux I__7281 (
            .O(N__45482),
            .I(\pid_front.pid_preregZ0Z_11 ));
    InMux I__7280 (
            .O(N__45477),
            .I(N__45473));
    InMux I__7279 (
            .O(N__45476),
            .I(N__45470));
    LocalMux I__7278 (
            .O(N__45473),
            .I(N__45465));
    LocalMux I__7277 (
            .O(N__45470),
            .I(N__45465));
    Odrv12 I__7276 (
            .O(N__45465),
            .I(front_order_11));
    CascadeMux I__7275 (
            .O(N__45462),
            .I(N__45450));
    CascadeMux I__7274 (
            .O(N__45461),
            .I(N__45447));
    CascadeMux I__7273 (
            .O(N__45460),
            .I(N__45442));
    CascadeMux I__7272 (
            .O(N__45459),
            .I(N__45439));
    InMux I__7271 (
            .O(N__45458),
            .I(N__45436));
    InMux I__7270 (
            .O(N__45457),
            .I(N__45429));
    InMux I__7269 (
            .O(N__45456),
            .I(N__45429));
    InMux I__7268 (
            .O(N__45455),
            .I(N__45429));
    InMux I__7267 (
            .O(N__45454),
            .I(N__45420));
    InMux I__7266 (
            .O(N__45453),
            .I(N__45420));
    InMux I__7265 (
            .O(N__45450),
            .I(N__45420));
    InMux I__7264 (
            .O(N__45447),
            .I(N__45420));
    InMux I__7263 (
            .O(N__45446),
            .I(N__45415));
    InMux I__7262 (
            .O(N__45445),
            .I(N__45415));
    InMux I__7261 (
            .O(N__45442),
            .I(N__45410));
    InMux I__7260 (
            .O(N__45439),
            .I(N__45410));
    LocalMux I__7259 (
            .O(N__45436),
            .I(N__45405));
    LocalMux I__7258 (
            .O(N__45429),
            .I(N__45405));
    LocalMux I__7257 (
            .O(N__45420),
            .I(N__45400));
    LocalMux I__7256 (
            .O(N__45415),
            .I(N__45400));
    LocalMux I__7255 (
            .O(N__45410),
            .I(N__45397));
    Span4Mux_h I__7254 (
            .O(N__45405),
            .I(N__45394));
    Span4Mux_h I__7253 (
            .O(N__45400),
            .I(N__45391));
    Odrv4 I__7252 (
            .O(N__45397),
            .I(\pid_front.N_76 ));
    Odrv4 I__7251 (
            .O(N__45394),
            .I(\pid_front.N_76 ));
    Odrv4 I__7250 (
            .O(N__45391),
            .I(\pid_front.N_76 ));
    InMux I__7249 (
            .O(N__45384),
            .I(N__45370));
    CascadeMux I__7248 (
            .O(N__45383),
            .I(N__45367));
    InMux I__7247 (
            .O(N__45382),
            .I(N__45362));
    CascadeMux I__7246 (
            .O(N__45381),
            .I(N__45359));
    CascadeMux I__7245 (
            .O(N__45380),
            .I(N__45356));
    CascadeMux I__7244 (
            .O(N__45379),
            .I(N__45353));
    InMux I__7243 (
            .O(N__45378),
            .I(N__45344));
    InMux I__7242 (
            .O(N__45377),
            .I(N__45344));
    InMux I__7241 (
            .O(N__45376),
            .I(N__45339));
    InMux I__7240 (
            .O(N__45375),
            .I(N__45339));
    InMux I__7239 (
            .O(N__45374),
            .I(N__45334));
    InMux I__7238 (
            .O(N__45373),
            .I(N__45334));
    LocalMux I__7237 (
            .O(N__45370),
            .I(N__45331));
    InMux I__7236 (
            .O(N__45367),
            .I(N__45328));
    InMux I__7235 (
            .O(N__45366),
            .I(N__45323));
    InMux I__7234 (
            .O(N__45365),
            .I(N__45323));
    LocalMux I__7233 (
            .O(N__45362),
            .I(N__45320));
    InMux I__7232 (
            .O(N__45359),
            .I(N__45313));
    InMux I__7231 (
            .O(N__45356),
            .I(N__45313));
    InMux I__7230 (
            .O(N__45353),
            .I(N__45313));
    InMux I__7229 (
            .O(N__45352),
            .I(N__45304));
    InMux I__7228 (
            .O(N__45351),
            .I(N__45304));
    InMux I__7227 (
            .O(N__45350),
            .I(N__45304));
    InMux I__7226 (
            .O(N__45349),
            .I(N__45304));
    LocalMux I__7225 (
            .O(N__45344),
            .I(N__45299));
    LocalMux I__7224 (
            .O(N__45339),
            .I(N__45299));
    LocalMux I__7223 (
            .O(N__45334),
            .I(N__45296));
    Span4Mux_h I__7222 (
            .O(N__45331),
            .I(N__45293));
    LocalMux I__7221 (
            .O(N__45328),
            .I(N__45290));
    LocalMux I__7220 (
            .O(N__45323),
            .I(N__45281));
    Span4Mux_h I__7219 (
            .O(N__45320),
            .I(N__45281));
    LocalMux I__7218 (
            .O(N__45313),
            .I(N__45281));
    LocalMux I__7217 (
            .O(N__45304),
            .I(N__45281));
    Span4Mux_v I__7216 (
            .O(N__45299),
            .I(N__45278));
    Span12Mux_v I__7215 (
            .O(N__45296),
            .I(N__45275));
    Span4Mux_v I__7214 (
            .O(N__45293),
            .I(N__45272));
    Span4Mux_v I__7213 (
            .O(N__45290),
            .I(N__45267));
    Span4Mux_v I__7212 (
            .O(N__45281),
            .I(N__45267));
    Odrv4 I__7211 (
            .O(N__45278),
            .I(\pid_front.pid_preregZ0Z_30 ));
    Odrv12 I__7210 (
            .O(N__45275),
            .I(\pid_front.pid_preregZ0Z_30 ));
    Odrv4 I__7209 (
            .O(N__45272),
            .I(\pid_front.pid_preregZ0Z_30 ));
    Odrv4 I__7208 (
            .O(N__45267),
            .I(\pid_front.pid_preregZ0Z_30 ));
    InMux I__7207 (
            .O(N__45258),
            .I(N__45255));
    LocalMux I__7206 (
            .O(N__45255),
            .I(N__45250));
    InMux I__7205 (
            .O(N__45254),
            .I(N__45245));
    InMux I__7204 (
            .O(N__45253),
            .I(N__45245));
    Odrv4 I__7203 (
            .O(N__45250),
            .I(\pid_front.pid_preregZ0Z_10 ));
    LocalMux I__7202 (
            .O(N__45245),
            .I(\pid_front.pid_preregZ0Z_10 ));
    InMux I__7201 (
            .O(N__45240),
            .I(N__45237));
    LocalMux I__7200 (
            .O(N__45237),
            .I(N__45233));
    InMux I__7199 (
            .O(N__45236),
            .I(N__45230));
    Span12Mux_s9_v I__7198 (
            .O(N__45233),
            .I(N__45225));
    LocalMux I__7197 (
            .O(N__45230),
            .I(N__45225));
    Odrv12 I__7196 (
            .O(N__45225),
            .I(front_order_10));
    CEMux I__7195 (
            .O(N__45222),
            .I(N__45219));
    LocalMux I__7194 (
            .O(N__45219),
            .I(N__45216));
    Span4Mux_v I__7193 (
            .O(N__45216),
            .I(N__45208));
    CEMux I__7192 (
            .O(N__45215),
            .I(N__45205));
    CEMux I__7191 (
            .O(N__45214),
            .I(N__45202));
    CEMux I__7190 (
            .O(N__45213),
            .I(N__45199));
    CEMux I__7189 (
            .O(N__45212),
            .I(N__45196));
    CEMux I__7188 (
            .O(N__45211),
            .I(N__45193));
    Odrv4 I__7187 (
            .O(N__45208),
            .I(\pid_front.state_0_1 ));
    LocalMux I__7186 (
            .O(N__45205),
            .I(\pid_front.state_0_1 ));
    LocalMux I__7185 (
            .O(N__45202),
            .I(\pid_front.state_0_1 ));
    LocalMux I__7184 (
            .O(N__45199),
            .I(\pid_front.state_0_1 ));
    LocalMux I__7183 (
            .O(N__45196),
            .I(\pid_front.state_0_1 ));
    LocalMux I__7182 (
            .O(N__45193),
            .I(\pid_front.state_0_1 ));
    SRMux I__7181 (
            .O(N__45180),
            .I(N__45177));
    LocalMux I__7180 (
            .O(N__45177),
            .I(N__45173));
    SRMux I__7179 (
            .O(N__45176),
            .I(N__45170));
    Span4Mux_v I__7178 (
            .O(N__45173),
            .I(N__45161));
    LocalMux I__7177 (
            .O(N__45170),
            .I(N__45161));
    SRMux I__7176 (
            .O(N__45169),
            .I(N__45158));
    SRMux I__7175 (
            .O(N__45168),
            .I(N__45155));
    SRMux I__7174 (
            .O(N__45167),
            .I(N__45152));
    SRMux I__7173 (
            .O(N__45166),
            .I(N__45149));
    Span4Mux_v I__7172 (
            .O(N__45161),
            .I(N__45144));
    LocalMux I__7171 (
            .O(N__45158),
            .I(N__45144));
    LocalMux I__7170 (
            .O(N__45155),
            .I(N__45141));
    LocalMux I__7169 (
            .O(N__45152),
            .I(N__45138));
    LocalMux I__7168 (
            .O(N__45149),
            .I(N__45133));
    Span4Mux_h I__7167 (
            .O(N__45144),
            .I(N__45133));
    Odrv4 I__7166 (
            .O(N__45141),
            .I(\pid_front.un1_reset_0_i ));
    Odrv4 I__7165 (
            .O(N__45138),
            .I(\pid_front.un1_reset_0_i ));
    Odrv4 I__7164 (
            .O(N__45133),
            .I(\pid_front.un1_reset_0_i ));
    InMux I__7163 (
            .O(N__45126),
            .I(N__45123));
    LocalMux I__7162 (
            .O(N__45123),
            .I(\pid_front.error_p_reg_esr_RNID8VU1Z0Z_3 ));
    CascadeMux I__7161 (
            .O(N__45120),
            .I(N__45117));
    InMux I__7160 (
            .O(N__45117),
            .I(N__45114));
    LocalMux I__7159 (
            .O(N__45114),
            .I(\pid_front.error_p_reg_esr_RNIUAE8_0Z0Z_4 ));
    InMux I__7158 (
            .O(N__45111),
            .I(N__45107));
    InMux I__7157 (
            .O(N__45110),
            .I(N__45104));
    LocalMux I__7156 (
            .O(N__45107),
            .I(N__45101));
    LocalMux I__7155 (
            .O(N__45104),
            .I(N__45098));
    Span12Mux_s7_v I__7154 (
            .O(N__45101),
            .I(N__45095));
    Span4Mux_h I__7153 (
            .O(N__45098),
            .I(N__45092));
    Odrv12 I__7152 (
            .O(N__45095),
            .I(front_order_5));
    Odrv4 I__7151 (
            .O(N__45092),
            .I(front_order_5));
    InMux I__7150 (
            .O(N__45087),
            .I(N__45084));
    LocalMux I__7149 (
            .O(N__45084),
            .I(N__45081));
    Span12Mux_s10_v I__7148 (
            .O(N__45081),
            .I(N__45078));
    Odrv12 I__7147 (
            .O(N__45078),
            .I(\ppm_encoder_1.un1_elevator_cry_4_THRU_CO ));
    InMux I__7146 (
            .O(N__45075),
            .I(\ppm_encoder_1.un1_elevator_cry_4 ));
    InMux I__7145 (
            .O(N__45072),
            .I(\ppm_encoder_1.un1_elevator_cry_5 ));
    InMux I__7144 (
            .O(N__45069),
            .I(\ppm_encoder_1.un1_elevator_cry_6 ));
    InMux I__7143 (
            .O(N__45066),
            .I(N__45063));
    LocalMux I__7142 (
            .O(N__45063),
            .I(N__45060));
    Odrv4 I__7141 (
            .O(N__45060),
            .I(\ppm_encoder_1.un1_elevator_cry_7_THRU_CO ));
    InMux I__7140 (
            .O(N__45057),
            .I(bfn_10_12_0_));
    InMux I__7139 (
            .O(N__45054),
            .I(N__45051));
    LocalMux I__7138 (
            .O(N__45051),
            .I(N__45047));
    InMux I__7137 (
            .O(N__45050),
            .I(N__45044));
    Span4Mux_v I__7136 (
            .O(N__45047),
            .I(N__45039));
    LocalMux I__7135 (
            .O(N__45044),
            .I(N__45039));
    Odrv4 I__7134 (
            .O(N__45039),
            .I(front_order_9));
    InMux I__7133 (
            .O(N__45036),
            .I(N__45033));
    LocalMux I__7132 (
            .O(N__45033),
            .I(N__45030));
    Odrv4 I__7131 (
            .O(N__45030),
            .I(\ppm_encoder_1.un1_elevator_cry_8_THRU_CO ));
    InMux I__7130 (
            .O(N__45027),
            .I(\ppm_encoder_1.un1_elevator_cry_8 ));
    InMux I__7129 (
            .O(N__45024),
            .I(N__45021));
    LocalMux I__7128 (
            .O(N__45021),
            .I(N__45018));
    Odrv4 I__7127 (
            .O(N__45018),
            .I(\ppm_encoder_1.un1_elevator_cry_9_THRU_CO ));
    InMux I__7126 (
            .O(N__45015),
            .I(\ppm_encoder_1.un1_elevator_cry_9 ));
    InMux I__7125 (
            .O(N__45012),
            .I(N__45009));
    LocalMux I__7124 (
            .O(N__45009),
            .I(N__45006));
    Odrv12 I__7123 (
            .O(N__45006),
            .I(\ppm_encoder_1.un1_elevator_cry_10_THRU_CO ));
    InMux I__7122 (
            .O(N__45003),
            .I(\ppm_encoder_1.un1_elevator_cry_10 ));
    InMux I__7121 (
            .O(N__45000),
            .I(N__44997));
    LocalMux I__7120 (
            .O(N__44997),
            .I(N__44994));
    Odrv12 I__7119 (
            .O(N__44994),
            .I(\ppm_encoder_1.un1_elevator_cry_11_THRU_CO ));
    InMux I__7118 (
            .O(N__44991),
            .I(\ppm_encoder_1.un1_elevator_cry_11 ));
    InMux I__7117 (
            .O(N__44988),
            .I(N__44985));
    LocalMux I__7116 (
            .O(N__44985),
            .I(N__44982));
    Odrv4 I__7115 (
            .O(N__44982),
            .I(\ppm_encoder_1.un1_elevator_cry_12_THRU_CO ));
    InMux I__7114 (
            .O(N__44979),
            .I(\ppm_encoder_1.un1_elevator_cry_12 ));
    CascadeMux I__7113 (
            .O(N__44976),
            .I(N__44973));
    InMux I__7112 (
            .O(N__44973),
            .I(N__44967));
    InMux I__7111 (
            .O(N__44972),
            .I(N__44967));
    LocalMux I__7110 (
            .O(N__44967),
            .I(N__44960));
    InMux I__7109 (
            .O(N__44966),
            .I(N__44955));
    InMux I__7108 (
            .O(N__44965),
            .I(N__44955));
    CascadeMux I__7107 (
            .O(N__44964),
            .I(N__44950));
    InMux I__7106 (
            .O(N__44963),
            .I(N__44947));
    Span4Mux_h I__7105 (
            .O(N__44960),
            .I(N__44944));
    LocalMux I__7104 (
            .O(N__44955),
            .I(N__44941));
    InMux I__7103 (
            .O(N__44954),
            .I(N__44934));
    InMux I__7102 (
            .O(N__44953),
            .I(N__44934));
    InMux I__7101 (
            .O(N__44950),
            .I(N__44934));
    LocalMux I__7100 (
            .O(N__44947),
            .I(\uart_drone.stateZ0Z_3 ));
    Odrv4 I__7099 (
            .O(N__44944),
            .I(\uart_drone.stateZ0Z_3 ));
    Odrv12 I__7098 (
            .O(N__44941),
            .I(\uart_drone.stateZ0Z_3 ));
    LocalMux I__7097 (
            .O(N__44934),
            .I(\uart_drone.stateZ0Z_3 ));
    CascadeMux I__7096 (
            .O(N__44925),
            .I(\uart_drone.N_152_cascade_ ));
    CascadeMux I__7095 (
            .O(N__44922),
            .I(N__44919));
    InMux I__7094 (
            .O(N__44919),
            .I(N__44916));
    LocalMux I__7093 (
            .O(N__44916),
            .I(N__44912));
    InMux I__7092 (
            .O(N__44915),
            .I(N__44909));
    Span4Mux_h I__7091 (
            .O(N__44912),
            .I(N__44904));
    LocalMux I__7090 (
            .O(N__44909),
            .I(N__44904));
    Span4Mux_v I__7089 (
            .O(N__44904),
            .I(N__44901));
    Odrv4 I__7088 (
            .O(N__44901),
            .I(front_order_1));
    InMux I__7087 (
            .O(N__44898),
            .I(N__44895));
    LocalMux I__7086 (
            .O(N__44895),
            .I(N__44892));
    Odrv4 I__7085 (
            .O(N__44892),
            .I(\ppm_encoder_1.un1_elevator_cry_0_THRU_CO ));
    InMux I__7084 (
            .O(N__44889),
            .I(\ppm_encoder_1.un1_elevator_cry_0 ));
    InMux I__7083 (
            .O(N__44886),
            .I(N__44883));
    LocalMux I__7082 (
            .O(N__44883),
            .I(N__44879));
    InMux I__7081 (
            .O(N__44882),
            .I(N__44876));
    Span4Mux_v I__7080 (
            .O(N__44879),
            .I(N__44871));
    LocalMux I__7079 (
            .O(N__44876),
            .I(N__44871));
    Span4Mux_v I__7078 (
            .O(N__44871),
            .I(N__44868));
    Odrv4 I__7077 (
            .O(N__44868),
            .I(front_order_2));
    InMux I__7076 (
            .O(N__44865),
            .I(N__44862));
    LocalMux I__7075 (
            .O(N__44862),
            .I(N__44859));
    Odrv12 I__7074 (
            .O(N__44859),
            .I(\ppm_encoder_1.un1_elevator_cry_1_THRU_CO ));
    InMux I__7073 (
            .O(N__44856),
            .I(\ppm_encoder_1.un1_elevator_cry_1 ));
    InMux I__7072 (
            .O(N__44853),
            .I(N__44850));
    LocalMux I__7071 (
            .O(N__44850),
            .I(N__44846));
    InMux I__7070 (
            .O(N__44849),
            .I(N__44843));
    Span4Mux_v I__7069 (
            .O(N__44846),
            .I(N__44840));
    LocalMux I__7068 (
            .O(N__44843),
            .I(N__44837));
    Span4Mux_v I__7067 (
            .O(N__44840),
            .I(N__44834));
    Span4Mux_v I__7066 (
            .O(N__44837),
            .I(N__44831));
    Odrv4 I__7065 (
            .O(N__44834),
            .I(front_order_3));
    Odrv4 I__7064 (
            .O(N__44831),
            .I(front_order_3));
    InMux I__7063 (
            .O(N__44826),
            .I(N__44823));
    LocalMux I__7062 (
            .O(N__44823),
            .I(N__44820));
    Odrv4 I__7061 (
            .O(N__44820),
            .I(\ppm_encoder_1.un1_elevator_cry_2_THRU_CO ));
    InMux I__7060 (
            .O(N__44817),
            .I(\ppm_encoder_1.un1_elevator_cry_2 ));
    InMux I__7059 (
            .O(N__44814),
            .I(N__44810));
    InMux I__7058 (
            .O(N__44813),
            .I(N__44807));
    LocalMux I__7057 (
            .O(N__44810),
            .I(N__44804));
    LocalMux I__7056 (
            .O(N__44807),
            .I(N__44801));
    Span12Mux_s6_v I__7055 (
            .O(N__44804),
            .I(N__44798));
    Span4Mux_h I__7054 (
            .O(N__44801),
            .I(N__44795));
    Odrv12 I__7053 (
            .O(N__44798),
            .I(front_order_4));
    Odrv4 I__7052 (
            .O(N__44795),
            .I(front_order_4));
    InMux I__7051 (
            .O(N__44790),
            .I(N__44787));
    LocalMux I__7050 (
            .O(N__44787),
            .I(N__44784));
    Span4Mux_v I__7049 (
            .O(N__44784),
            .I(N__44781));
    Odrv4 I__7048 (
            .O(N__44781),
            .I(\ppm_encoder_1.un1_elevator_cry_3_THRU_CO ));
    InMux I__7047 (
            .O(N__44778),
            .I(\ppm_encoder_1.un1_elevator_cry_3 ));
    CascadeMux I__7046 (
            .O(N__44775),
            .I(N__44770));
    InMux I__7045 (
            .O(N__44774),
            .I(N__44765));
    InMux I__7044 (
            .O(N__44773),
            .I(N__44765));
    InMux I__7043 (
            .O(N__44770),
            .I(N__44762));
    LocalMux I__7042 (
            .O(N__44765),
            .I(N__44759));
    LocalMux I__7041 (
            .O(N__44762),
            .I(N__44754));
    Span4Mux_h I__7040 (
            .O(N__44759),
            .I(N__44754));
    Odrv4 I__7039 (
            .O(N__44754),
            .I(\ppm_encoder_1.aileronZ0Z_4 ));
    CascadeMux I__7038 (
            .O(N__44751),
            .I(N__44747));
    InMux I__7037 (
            .O(N__44750),
            .I(N__44744));
    InMux I__7036 (
            .O(N__44747),
            .I(N__44741));
    LocalMux I__7035 (
            .O(N__44744),
            .I(N__44734));
    LocalMux I__7034 (
            .O(N__44741),
            .I(N__44734));
    CascadeMux I__7033 (
            .O(N__44740),
            .I(N__44731));
    InMux I__7032 (
            .O(N__44739),
            .I(N__44728));
    Span4Mux_h I__7031 (
            .O(N__44734),
            .I(N__44725));
    InMux I__7030 (
            .O(N__44731),
            .I(N__44722));
    LocalMux I__7029 (
            .O(N__44728),
            .I(\uart_drone.stateZ0Z_2 ));
    Odrv4 I__7028 (
            .O(N__44725),
            .I(\uart_drone.stateZ0Z_2 ));
    LocalMux I__7027 (
            .O(N__44722),
            .I(\uart_drone.stateZ0Z_2 ));
    CascadeMux I__7026 (
            .O(N__44715),
            .I(\uart_drone.N_145_cascade_ ));
    InMux I__7025 (
            .O(N__44712),
            .I(N__44703));
    InMux I__7024 (
            .O(N__44711),
            .I(N__44703));
    InMux I__7023 (
            .O(N__44710),
            .I(N__44700));
    InMux I__7022 (
            .O(N__44709),
            .I(N__44694));
    InMux I__7021 (
            .O(N__44708),
            .I(N__44694));
    LocalMux I__7020 (
            .O(N__44703),
            .I(N__44691));
    LocalMux I__7019 (
            .O(N__44700),
            .I(N__44688));
    InMux I__7018 (
            .O(N__44699),
            .I(N__44685));
    LocalMux I__7017 (
            .O(N__44694),
            .I(\uart_drone.stateZ0Z_4 ));
    Odrv4 I__7016 (
            .O(N__44691),
            .I(\uart_drone.stateZ0Z_4 ));
    Odrv4 I__7015 (
            .O(N__44688),
            .I(\uart_drone.stateZ0Z_4 ));
    LocalMux I__7014 (
            .O(N__44685),
            .I(\uart_drone.stateZ0Z_4 ));
    CascadeMux I__7013 (
            .O(N__44676),
            .I(\uart_drone.un1_state_4_0_cascade_ ));
    InMux I__7012 (
            .O(N__44673),
            .I(N__44670));
    LocalMux I__7011 (
            .O(N__44670),
            .I(N__44667));
    Span4Mux_v I__7010 (
            .O(N__44667),
            .I(N__44664));
    Odrv4 I__7009 (
            .O(N__44664),
            .I(\ppm_encoder_1.un1_throttle_cry_9_THRU_CO ));
    InMux I__7008 (
            .O(N__44661),
            .I(N__44658));
    LocalMux I__7007 (
            .O(N__44658),
            .I(N__44653));
    InMux I__7006 (
            .O(N__44657),
            .I(N__44650));
    CascadeMux I__7005 (
            .O(N__44656),
            .I(N__44647));
    Span4Mux_h I__7004 (
            .O(N__44653),
            .I(N__44644));
    LocalMux I__7003 (
            .O(N__44650),
            .I(N__44641));
    InMux I__7002 (
            .O(N__44647),
            .I(N__44638));
    Span4Mux_h I__7001 (
            .O(N__44644),
            .I(N__44635));
    Span4Mux_v I__7000 (
            .O(N__44641),
            .I(N__44632));
    LocalMux I__6999 (
            .O(N__44638),
            .I(throttle_order_10));
    Odrv4 I__6998 (
            .O(N__44635),
            .I(throttle_order_10));
    Odrv4 I__6997 (
            .O(N__44632),
            .I(throttle_order_10));
    InMux I__6996 (
            .O(N__44625),
            .I(N__44622));
    LocalMux I__6995 (
            .O(N__44622),
            .I(N__44618));
    InMux I__6994 (
            .O(N__44621),
            .I(N__44615));
    Span4Mux_h I__6993 (
            .O(N__44618),
            .I(N__44612));
    LocalMux I__6992 (
            .O(N__44615),
            .I(N__44609));
    Span4Mux_h I__6991 (
            .O(N__44612),
            .I(N__44606));
    Span4Mux_h I__6990 (
            .O(N__44609),
            .I(N__44603));
    Odrv4 I__6989 (
            .O(N__44606),
            .I(throttle_order_13));
    Odrv4 I__6988 (
            .O(N__44603),
            .I(throttle_order_13));
    InMux I__6987 (
            .O(N__44598),
            .I(N__44595));
    LocalMux I__6986 (
            .O(N__44595),
            .I(N__44592));
    Span4Mux_h I__6985 (
            .O(N__44592),
            .I(N__44589));
    Odrv4 I__6984 (
            .O(N__44589),
            .I(\ppm_encoder_1.un1_throttle_cry_12_THRU_CO ));
    InMux I__6983 (
            .O(N__44586),
            .I(N__44583));
    LocalMux I__6982 (
            .O(N__44583),
            .I(N__44580));
    Span4Mux_h I__6981 (
            .O(N__44580),
            .I(N__44577));
    Odrv4 I__6980 (
            .O(N__44577),
            .I(\ppm_encoder_1.un1_throttle_cry_1_THRU_CO ));
    InMux I__6979 (
            .O(N__44574),
            .I(N__44571));
    LocalMux I__6978 (
            .O(N__44571),
            .I(N__44567));
    InMux I__6977 (
            .O(N__44570),
            .I(N__44564));
    Span4Mux_h I__6976 (
            .O(N__44567),
            .I(N__44559));
    LocalMux I__6975 (
            .O(N__44564),
            .I(N__44559));
    Span4Mux_v I__6974 (
            .O(N__44559),
            .I(N__44556));
    Odrv4 I__6973 (
            .O(N__44556),
            .I(throttle_order_2));
    CascadeMux I__6972 (
            .O(N__44553),
            .I(N__44548));
    InMux I__6971 (
            .O(N__44552),
            .I(N__44545));
    CascadeMux I__6970 (
            .O(N__44551),
            .I(N__44542));
    InMux I__6969 (
            .O(N__44548),
            .I(N__44539));
    LocalMux I__6968 (
            .O(N__44545),
            .I(N__44536));
    InMux I__6967 (
            .O(N__44542),
            .I(N__44533));
    LocalMux I__6966 (
            .O(N__44539),
            .I(N__44530));
    Span4Mux_s2_v I__6965 (
            .O(N__44536),
            .I(N__44527));
    LocalMux I__6964 (
            .O(N__44533),
            .I(\ppm_encoder_1.aileronZ0Z_5 ));
    Odrv4 I__6963 (
            .O(N__44530),
            .I(\ppm_encoder_1.aileronZ0Z_5 ));
    Odrv4 I__6962 (
            .O(N__44527),
            .I(\ppm_encoder_1.aileronZ0Z_5 ));
    InMux I__6961 (
            .O(N__44520),
            .I(N__44517));
    LocalMux I__6960 (
            .O(N__44517),
            .I(\ppm_encoder_1.un1_rudder_cry_9_THRU_CO ));
    CascadeMux I__6959 (
            .O(N__44514),
            .I(N__44511));
    InMux I__6958 (
            .O(N__44511),
            .I(N__44507));
    InMux I__6957 (
            .O(N__44510),
            .I(N__44504));
    LocalMux I__6956 (
            .O(N__44507),
            .I(N__44499));
    LocalMux I__6955 (
            .O(N__44504),
            .I(N__44499));
    Odrv4 I__6954 (
            .O(N__44499),
            .I(scaler_4_data_10));
    InMux I__6953 (
            .O(N__44496),
            .I(N__44493));
    LocalMux I__6952 (
            .O(N__44493),
            .I(\ppm_encoder_1.un1_rudder_cry_11_THRU_CO ));
    InMux I__6951 (
            .O(N__44490),
            .I(N__44486));
    CascadeMux I__6950 (
            .O(N__44489),
            .I(N__44483));
    LocalMux I__6949 (
            .O(N__44486),
            .I(N__44480));
    InMux I__6948 (
            .O(N__44483),
            .I(N__44477));
    Span4Mux_h I__6947 (
            .O(N__44480),
            .I(N__44474));
    LocalMux I__6946 (
            .O(N__44477),
            .I(N__44471));
    Odrv4 I__6945 (
            .O(N__44474),
            .I(scaler_4_data_12));
    Odrv4 I__6944 (
            .O(N__44471),
            .I(scaler_4_data_12));
    InMux I__6943 (
            .O(N__44466),
            .I(N__44463));
    LocalMux I__6942 (
            .O(N__44463),
            .I(\ppm_encoder_1.un1_rudder_cry_6_THRU_CO ));
    InMux I__6941 (
            .O(N__44460),
            .I(N__44456));
    InMux I__6940 (
            .O(N__44459),
            .I(N__44453));
    LocalMux I__6939 (
            .O(N__44456),
            .I(N__44450));
    LocalMux I__6938 (
            .O(N__44453),
            .I(N__44447));
    Odrv4 I__6937 (
            .O(N__44450),
            .I(scaler_4_data_7));
    Odrv4 I__6936 (
            .O(N__44447),
            .I(scaler_4_data_7));
    InMux I__6935 (
            .O(N__44442),
            .I(N__44439));
    LocalMux I__6934 (
            .O(N__44439),
            .I(\ppm_encoder_1.un1_rudder_cry_7_THRU_CO ));
    InMux I__6933 (
            .O(N__44436),
            .I(N__44433));
    LocalMux I__6932 (
            .O(N__44433),
            .I(N__44429));
    InMux I__6931 (
            .O(N__44432),
            .I(N__44426));
    Span4Mux_v I__6930 (
            .O(N__44429),
            .I(N__44423));
    LocalMux I__6929 (
            .O(N__44426),
            .I(N__44420));
    Odrv4 I__6928 (
            .O(N__44423),
            .I(scaler_4_data_8));
    Odrv4 I__6927 (
            .O(N__44420),
            .I(scaler_4_data_8));
    InMux I__6926 (
            .O(N__44415),
            .I(N__44411));
    InMux I__6925 (
            .O(N__44414),
            .I(N__44408));
    LocalMux I__6924 (
            .O(N__44411),
            .I(N__44405));
    LocalMux I__6923 (
            .O(N__44408),
            .I(scaler_4_data_9));
    Odrv4 I__6922 (
            .O(N__44405),
            .I(scaler_4_data_9));
    InMux I__6921 (
            .O(N__44400),
            .I(N__44397));
    LocalMux I__6920 (
            .O(N__44397),
            .I(\ppm_encoder_1.un1_rudder_cry_8_THRU_CO ));
    CascadeMux I__6919 (
            .O(N__44394),
            .I(\ppm_encoder_1.counter24_0_I_57_c_RNIJMMDZ0_cascade_ ));
    IoInMux I__6918 (
            .O(N__44391),
            .I(N__44388));
    LocalMux I__6917 (
            .O(N__44388),
            .I(N__44385));
    IoSpan4Mux I__6916 (
            .O(N__44385),
            .I(N__44382));
    Span4Mux_s2_v I__6915 (
            .O(N__44382),
            .I(N__44378));
    InMux I__6914 (
            .O(N__44381),
            .I(N__44375));
    Odrv4 I__6913 (
            .O(N__44378),
            .I(ppm_output_c));
    LocalMux I__6912 (
            .O(N__44375),
            .I(ppm_output_c));
    InMux I__6911 (
            .O(N__44370),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_12 ));
    InMux I__6910 (
            .O(N__44367),
            .I(N__44364));
    LocalMux I__6909 (
            .O(N__44364),
            .I(N__44361));
    Span4Mux_s1_v I__6908 (
            .O(N__44361),
            .I(N__44358));
    Odrv4 I__6907 (
            .O(N__44358),
            .I(\ppm_encoder_1.un1_init_pulses_10_14 ));
    InMux I__6906 (
            .O(N__44355),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_13 ));
    InMux I__6905 (
            .O(N__44352),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_14 ));
    InMux I__6904 (
            .O(N__44349),
            .I(bfn_10_5_0_));
    InMux I__6903 (
            .O(N__44346),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_16 ));
    InMux I__6902 (
            .O(N__44343),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_17 ));
    CascadeMux I__6901 (
            .O(N__44340),
            .I(N__44337));
    InMux I__6900 (
            .O(N__44337),
            .I(N__44334));
    LocalMux I__6899 (
            .O(N__44334),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_16 ));
    InMux I__6898 (
            .O(N__44331),
            .I(N__44328));
    LocalMux I__6897 (
            .O(N__44328),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_17 ));
    InMux I__6896 (
            .O(N__44325),
            .I(N__44322));
    LocalMux I__6895 (
            .O(N__44322),
            .I(\ppm_encoder_1.un2_throttle_iv_0_1_3 ));
    InMux I__6894 (
            .O(N__44319),
            .I(N__44316));
    LocalMux I__6893 (
            .O(N__44316),
            .I(\ppm_encoder_1.init_pulses_RNISKNT5Z0Z_5 ));
    CascadeMux I__6892 (
            .O(N__44313),
            .I(N__44310));
    InMux I__6891 (
            .O(N__44310),
            .I(N__44306));
    InMux I__6890 (
            .O(N__44309),
            .I(N__44303));
    LocalMux I__6889 (
            .O(N__44306),
            .I(\ppm_encoder_1.N_261_i_i ));
    LocalMux I__6888 (
            .O(N__44303),
            .I(\ppm_encoder_1.N_261_i_i ));
    InMux I__6887 (
            .O(N__44298),
            .I(N__44295));
    LocalMux I__6886 (
            .O(N__44295),
            .I(N__44292));
    Odrv4 I__6885 (
            .O(N__44292),
            .I(\ppm_encoder_1.un1_init_pulses_10_5 ));
    InMux I__6884 (
            .O(N__44289),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_4 ));
    InMux I__6883 (
            .O(N__44286),
            .I(N__44283));
    LocalMux I__6882 (
            .O(N__44283),
            .I(\ppm_encoder_1.un1_init_pulses_10_6 ));
    InMux I__6881 (
            .O(N__44280),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_5 ));
    InMux I__6880 (
            .O(N__44277),
            .I(N__44274));
    LocalMux I__6879 (
            .O(N__44274),
            .I(\ppm_encoder_1.un1_init_pulses_10_7 ));
    InMux I__6878 (
            .O(N__44271),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_6 ));
    InMux I__6877 (
            .O(N__44268),
            .I(N__44265));
    LocalMux I__6876 (
            .O(N__44265),
            .I(\ppm_encoder_1.init_pulses_RNI85KU5Z0Z_8 ));
    CascadeMux I__6875 (
            .O(N__44262),
            .I(N__44259));
    InMux I__6874 (
            .O(N__44259),
            .I(N__44255));
    InMux I__6873 (
            .O(N__44258),
            .I(N__44252));
    LocalMux I__6872 (
            .O(N__44255),
            .I(\ppm_encoder_1.N_264_i_i ));
    LocalMux I__6871 (
            .O(N__44252),
            .I(\ppm_encoder_1.N_264_i_i ));
    InMux I__6870 (
            .O(N__44247),
            .I(N__44244));
    LocalMux I__6869 (
            .O(N__44244),
            .I(N__44241));
    Odrv4 I__6868 (
            .O(N__44241),
            .I(\ppm_encoder_1.un1_init_pulses_10_8 ));
    InMux I__6867 (
            .O(N__44238),
            .I(bfn_10_4_0_));
    InMux I__6866 (
            .O(N__44235),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_8 ));
    InMux I__6865 (
            .O(N__44232),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_9 ));
    InMux I__6864 (
            .O(N__44229),
            .I(N__44226));
    LocalMux I__6863 (
            .O(N__44226),
            .I(N__44223));
    Odrv4 I__6862 (
            .O(N__44223),
            .I(\ppm_encoder_1.un1_init_pulses_10_11 ));
    InMux I__6861 (
            .O(N__44220),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_10 ));
    InMux I__6860 (
            .O(N__44217),
            .I(N__44214));
    LocalMux I__6859 (
            .O(N__44214),
            .I(N__44211));
    Odrv4 I__6858 (
            .O(N__44211),
            .I(\ppm_encoder_1.un1_init_pulses_10_12 ));
    InMux I__6857 (
            .O(N__44208),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_11 ));
    InMux I__6856 (
            .O(N__44205),
            .I(N__44201));
    CascadeMux I__6855 (
            .O(N__44204),
            .I(N__44198));
    LocalMux I__6854 (
            .O(N__44201),
            .I(N__44195));
    InMux I__6853 (
            .O(N__44198),
            .I(N__44192));
    Span4Mux_v I__6852 (
            .O(N__44195),
            .I(N__44187));
    LocalMux I__6851 (
            .O(N__44192),
            .I(N__44187));
    Odrv4 I__6850 (
            .O(N__44187),
            .I(scaler_4_data_11));
    InMux I__6849 (
            .O(N__44184),
            .I(N__44181));
    LocalMux I__6848 (
            .O(N__44181),
            .I(N__44178));
    Span4Mux_s1_v I__6847 (
            .O(N__44178),
            .I(N__44175));
    Odrv4 I__6846 (
            .O(N__44175),
            .I(\ppm_encoder_1.un1_rudder_cry_10_THRU_CO ));
    InMux I__6845 (
            .O(N__44172),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_0 ));
    InMux I__6844 (
            .O(N__44169),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_1 ));
    InMux I__6843 (
            .O(N__44166),
            .I(N__44163));
    LocalMux I__6842 (
            .O(N__44163),
            .I(\ppm_encoder_1.init_pulses_RNIALAI5Z0Z_3 ));
    CascadeMux I__6841 (
            .O(N__44160),
            .I(N__44157));
    InMux I__6840 (
            .O(N__44157),
            .I(N__44153));
    InMux I__6839 (
            .O(N__44156),
            .I(N__44150));
    LocalMux I__6838 (
            .O(N__44153),
            .I(\ppm_encoder_1.N_256_i_i ));
    LocalMux I__6837 (
            .O(N__44150),
            .I(\ppm_encoder_1.N_256_i_i ));
    InMux I__6836 (
            .O(N__44145),
            .I(N__44142));
    LocalMux I__6835 (
            .O(N__44142),
            .I(\ppm_encoder_1.un1_init_pulses_10_3 ));
    InMux I__6834 (
            .O(N__44139),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_2 ));
    InMux I__6833 (
            .O(N__44136),
            .I(N__44133));
    LocalMux I__6832 (
            .O(N__44133),
            .I(\ppm_encoder_1.init_pulses_RNIMENT5Z0Z_4 ));
    CascadeMux I__6831 (
            .O(N__44130),
            .I(N__44127));
    InMux I__6830 (
            .O(N__44127),
            .I(N__44123));
    InMux I__6829 (
            .O(N__44126),
            .I(N__44120));
    LocalMux I__6828 (
            .O(N__44123),
            .I(\ppm_encoder_1.N_260_i_i ));
    LocalMux I__6827 (
            .O(N__44120),
            .I(\ppm_encoder_1.N_260_i_i ));
    InMux I__6826 (
            .O(N__44115),
            .I(N__44112));
    LocalMux I__6825 (
            .O(N__44112),
            .I(\ppm_encoder_1.un1_init_pulses_10_4 ));
    InMux I__6824 (
            .O(N__44109),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_3 ));
    InMux I__6823 (
            .O(N__44106),
            .I(N__44100));
    InMux I__6822 (
            .O(N__44105),
            .I(N__44100));
    LocalMux I__6821 (
            .O(N__44100),
            .I(N__44097));
    Span4Mux_v I__6820 (
            .O(N__44097),
            .I(N__44094));
    Span4Mux_h I__6819 (
            .O(N__44094),
            .I(N__44091));
    Span4Mux_h I__6818 (
            .O(N__44091),
            .I(N__44088));
    Span4Mux_v I__6817 (
            .O(N__44088),
            .I(N__44085));
    Odrv4 I__6816 (
            .O(N__44085),
            .I(\pid_front.error_p_regZ0Z_16 ));
    InMux I__6815 (
            .O(N__44082),
            .I(N__44076));
    InMux I__6814 (
            .O(N__44081),
            .I(N__44076));
    LocalMux I__6813 (
            .O(N__44076),
            .I(\pid_front.error_d_reg_prevZ0Z_16 ));
    InMux I__6812 (
            .O(N__44073),
            .I(N__44070));
    LocalMux I__6811 (
            .O(N__44070),
            .I(N__44065));
    InMux I__6810 (
            .O(N__44069),
            .I(N__44060));
    InMux I__6809 (
            .O(N__44068),
            .I(N__44060));
    Odrv4 I__6808 (
            .O(N__44065),
            .I(\pid_front.un1_pid_prereg_0_0 ));
    LocalMux I__6807 (
            .O(N__44060),
            .I(\pid_front.un1_pid_prereg_0_0 ));
    CascadeMux I__6806 (
            .O(N__44055),
            .I(N__44052));
    InMux I__6805 (
            .O(N__44052),
            .I(N__44049));
    LocalMux I__6804 (
            .O(N__44049),
            .I(N__44045));
    InMux I__6803 (
            .O(N__44048),
            .I(N__44042));
    Odrv12 I__6802 (
            .O(N__44045),
            .I(\pid_front.un1_pid_prereg_0_1 ));
    LocalMux I__6801 (
            .O(N__44042),
            .I(\pid_front.un1_pid_prereg_0_1 ));
    InMux I__6800 (
            .O(N__44037),
            .I(N__44034));
    LocalMux I__6799 (
            .O(N__44034),
            .I(N__44031));
    Span4Mux_v I__6798 (
            .O(N__44031),
            .I(N__44028));
    Odrv4 I__6797 (
            .O(N__44028),
            .I(\pid_front.error_p_reg_esr_RNICIRCDZ0Z_14 ));
    CascadeMux I__6796 (
            .O(N__44025),
            .I(\pid_front.un1_pid_prereg_0_3_cascade_ ));
    CascadeMux I__6795 (
            .O(N__44022),
            .I(N__44019));
    InMux I__6794 (
            .O(N__44019),
            .I(N__44016));
    LocalMux I__6793 (
            .O(N__44016),
            .I(N__44013));
    Span4Mux_v I__6792 (
            .O(N__44013),
            .I(N__44010));
    Odrv4 I__6791 (
            .O(N__44010),
            .I(\pid_front.error_p_reg_esr_RNIE2FM6Z0Z_15 ));
    InMux I__6790 (
            .O(N__44007),
            .I(N__44001));
    InMux I__6789 (
            .O(N__44006),
            .I(N__44001));
    LocalMux I__6788 (
            .O(N__44001),
            .I(\pid_front.error_p_reg_esr_RNIN6C61Z0Z_16 ));
    InMux I__6787 (
            .O(N__43998),
            .I(N__43992));
    InMux I__6786 (
            .O(N__43997),
            .I(N__43992));
    LocalMux I__6785 (
            .O(N__43992),
            .I(\pid_front.un1_pid_prereg_0_3 ));
    CascadeMux I__6784 (
            .O(N__43989),
            .I(\pid_front.un1_pid_prereg_0_4_cascade_ ));
    InMux I__6783 (
            .O(N__43986),
            .I(N__43983));
    LocalMux I__6782 (
            .O(N__43983),
            .I(N__43980));
    Odrv12 I__6781 (
            .O(N__43980),
            .I(\pid_front.error_p_reg_esr_RNICN0DDZ0Z_15 ));
    CascadeMux I__6780 (
            .O(N__43977),
            .I(\pid_front.un1_pid_prereg_0_5_cascade_ ));
    CascadeMux I__6779 (
            .O(N__43974),
            .I(N__43971));
    InMux I__6778 (
            .O(N__43971),
            .I(N__43968));
    LocalMux I__6777 (
            .O(N__43968),
            .I(N__43965));
    Span4Mux_v I__6776 (
            .O(N__43965),
            .I(N__43962));
    Odrv4 I__6775 (
            .O(N__43962),
            .I(\pid_front.error_p_reg_esr_RNIUKHM6Z0Z_16 ));
    InMux I__6774 (
            .O(N__43959),
            .I(N__43955));
    InMux I__6773 (
            .O(N__43958),
            .I(N__43952));
    LocalMux I__6772 (
            .O(N__43955),
            .I(\pid_front.error_p_reg_esr_RNIK3C61Z0Z_15 ));
    LocalMux I__6771 (
            .O(N__43952),
            .I(\pid_front.error_p_reg_esr_RNIK3C61Z0Z_15 ));
    InMux I__6770 (
            .O(N__43947),
            .I(N__43944));
    LocalMux I__6769 (
            .O(N__43944),
            .I(N__43940));
    InMux I__6768 (
            .O(N__43943),
            .I(N__43937));
    Odrv4 I__6767 (
            .O(N__43940),
            .I(\pid_front.error_p_reg_esr_RNIN6C61_0Z0Z_16 ));
    LocalMux I__6766 (
            .O(N__43937),
            .I(\pid_front.error_p_reg_esr_RNIN6C61_0Z0Z_16 ));
    InMux I__6765 (
            .O(N__43932),
            .I(N__43927));
    InMux I__6764 (
            .O(N__43931),
            .I(N__43922));
    InMux I__6763 (
            .O(N__43930),
            .I(N__43922));
    LocalMux I__6762 (
            .O(N__43927),
            .I(\pid_front.un1_pid_prereg_0_2 ));
    LocalMux I__6761 (
            .O(N__43922),
            .I(\pid_front.un1_pid_prereg_0_2 ));
    InMux I__6760 (
            .O(N__43917),
            .I(N__43914));
    LocalMux I__6759 (
            .O(N__43914),
            .I(\pid_front.error_p_reg_esr_RNIH0C61Z0Z_14 ));
    InMux I__6758 (
            .O(N__43911),
            .I(N__43905));
    InMux I__6757 (
            .O(N__43910),
            .I(N__43905));
    LocalMux I__6756 (
            .O(N__43905),
            .I(\pid_front.error_d_reg_prev_esr_RNI5JRF4Z0Z_10 ));
    CascadeMux I__6755 (
            .O(N__43902),
            .I(N__43899));
    InMux I__6754 (
            .O(N__43899),
            .I(N__43893));
    InMux I__6753 (
            .O(N__43898),
            .I(N__43893));
    LocalMux I__6752 (
            .O(N__43893),
            .I(\pid_front.error_p_reg_esr_RNIK3C61_0Z0Z_15 ));
    InMux I__6751 (
            .O(N__43890),
            .I(N__43884));
    InMux I__6750 (
            .O(N__43889),
            .I(N__43884));
    LocalMux I__6749 (
            .O(N__43884),
            .I(N__43881));
    Span4Mux_v I__6748 (
            .O(N__43881),
            .I(N__43878));
    Span4Mux_h I__6747 (
            .O(N__43878),
            .I(N__43875));
    Span4Mux_h I__6746 (
            .O(N__43875),
            .I(N__43872));
    Span4Mux_v I__6745 (
            .O(N__43872),
            .I(N__43869));
    Odrv4 I__6744 (
            .O(N__43869),
            .I(\pid_front.error_p_regZ0Z_15 ));
    InMux I__6743 (
            .O(N__43866),
            .I(N__43860));
    InMux I__6742 (
            .O(N__43865),
            .I(N__43860));
    LocalMux I__6741 (
            .O(N__43860),
            .I(\pid_front.error_d_reg_prevZ0Z_15 ));
    CascadeMux I__6740 (
            .O(N__43857),
            .I(\pid_front.un1_pid_prereg_153_0_cascade_ ));
    InMux I__6739 (
            .O(N__43854),
            .I(N__43851));
    LocalMux I__6738 (
            .O(N__43851),
            .I(N__43848));
    Span4Mux_h I__6737 (
            .O(N__43848),
            .I(N__43845));
    Odrv4 I__6736 (
            .O(N__43845),
            .I(\pid_front.error_d_reg_prev_esr_RNIHM5CDZ0Z_10 ));
    CascadeMux I__6735 (
            .O(N__43842),
            .I(N__43839));
    InMux I__6734 (
            .O(N__43839),
            .I(N__43836));
    LocalMux I__6733 (
            .O(N__43836),
            .I(\pid_front.N_2191_i ));
    CascadeMux I__6732 (
            .O(N__43833),
            .I(\pid_front.N_2191_i_cascade_ ));
    InMux I__6731 (
            .O(N__43830),
            .I(N__43824));
    InMux I__6730 (
            .O(N__43829),
            .I(N__43824));
    LocalMux I__6729 (
            .O(N__43824),
            .I(\pid_front.error_p_reg_esr_RNILTVH2Z0Z_12 ));
    InMux I__6728 (
            .O(N__43821),
            .I(N__43818));
    LocalMux I__6727 (
            .O(N__43818),
            .I(N__43815));
    Span4Mux_h I__6726 (
            .O(N__43815),
            .I(N__43812));
    Odrv4 I__6725 (
            .O(N__43812),
            .I(\pid_front.error_p_reg_esr_RNIJVCREZ0Z_13 ));
    CascadeMux I__6724 (
            .O(N__43809),
            .I(N__43806));
    InMux I__6723 (
            .O(N__43806),
            .I(N__43803));
    LocalMux I__6722 (
            .O(N__43803),
            .I(N__43800));
    Odrv12 I__6721 (
            .O(N__43800),
            .I(\pid_front.error_p_reg_esr_RNIHFPHLZ0Z_13 ));
    CascadeMux I__6720 (
            .O(N__43797),
            .I(\pid_front.un1_pid_prereg_0_1_cascade_ ));
    CascadeMux I__6719 (
            .O(N__43794),
            .I(N__43791));
    InMux I__6718 (
            .O(N__43791),
            .I(N__43788));
    LocalMux I__6717 (
            .O(N__43788),
            .I(N__43785));
    Span4Mux_h I__6716 (
            .O(N__43785),
            .I(N__43782));
    Odrv4 I__6715 (
            .O(N__43782),
            .I(\pid_front.error_p_reg_esr_RNIUFCM6Z0Z_14 ));
    CascadeMux I__6714 (
            .O(N__43779),
            .I(\pid_front.error_p_reg_esr_RNIH0C61Z0Z_14_cascade_ ));
    CascadeMux I__6713 (
            .O(N__43776),
            .I(\pid_front.un1_pid_prereg_0_18_cascade_ ));
    InMux I__6712 (
            .O(N__43773),
            .I(N__43770));
    LocalMux I__6711 (
            .O(N__43770),
            .I(\pid_front.error_d_reg_prev_esr_RNIC2UN8Z0Z_22 ));
    InMux I__6710 (
            .O(N__43767),
            .I(N__43764));
    LocalMux I__6709 (
            .O(N__43764),
            .I(N__43760));
    InMux I__6708 (
            .O(N__43763),
            .I(N__43757));
    Odrv4 I__6707 (
            .O(N__43760),
            .I(\pid_front.un1_pid_prereg_0_17 ));
    LocalMux I__6706 (
            .O(N__43757),
            .I(\pid_front.un1_pid_prereg_0_17 ));
    InMux I__6705 (
            .O(N__43752),
            .I(N__43749));
    LocalMux I__6704 (
            .O(N__43749),
            .I(\pid_front.error_d_reg_prev_esr_RNIFJ8U9Z0Z_22 ));
    InMux I__6703 (
            .O(N__43746),
            .I(N__43742));
    InMux I__6702 (
            .O(N__43745),
            .I(N__43739));
    LocalMux I__6701 (
            .O(N__43742),
            .I(\pid_front.un1_pid_prereg_0_19 ));
    LocalMux I__6700 (
            .O(N__43739),
            .I(\pid_front.un1_pid_prereg_0_19 ));
    CascadeMux I__6699 (
            .O(N__43734),
            .I(\pid_front.un1_pid_prereg_0_19_cascade_ ));
    InMux I__6698 (
            .O(N__43731),
            .I(N__43727));
    InMux I__6697 (
            .O(N__43730),
            .I(N__43724));
    LocalMux I__6696 (
            .O(N__43727),
            .I(\pid_front.un1_pid_prereg_0_18 ));
    LocalMux I__6695 (
            .O(N__43724),
            .I(\pid_front.un1_pid_prereg_0_18 ));
    CascadeMux I__6694 (
            .O(N__43719),
            .I(N__43716));
    InMux I__6693 (
            .O(N__43716),
            .I(N__43713));
    LocalMux I__6692 (
            .O(N__43713),
            .I(\pid_front.error_d_reg_prev_esr_RNI840C4Z0Z_22 ));
    CascadeMux I__6691 (
            .O(N__43710),
            .I(N__43707));
    InMux I__6690 (
            .O(N__43707),
            .I(N__43704));
    LocalMux I__6689 (
            .O(N__43704),
            .I(N__43701));
    Odrv12 I__6688 (
            .O(N__43701),
            .I(\pid_front.error_p_reg_esr_RNI1IK9EZ0Z_12 ));
    CascadeMux I__6687 (
            .O(N__43698),
            .I(\pid_front.un1_pid_prereg_167_0_1_cascade_ ));
    InMux I__6686 (
            .O(N__43695),
            .I(N__43692));
    LocalMux I__6685 (
            .O(N__43692),
            .I(N__43689));
    Odrv4 I__6684 (
            .O(N__43689),
            .I(\pid_front.pid_preregZ0Z_25 ));
    InMux I__6683 (
            .O(N__43686),
            .I(\pid_front.un1_pid_prereg_0_cry_24 ));
    InMux I__6682 (
            .O(N__43683),
            .I(N__43680));
    LocalMux I__6681 (
            .O(N__43680),
            .I(\pid_front.error_d_reg_prev_esr_RNIKE2O8Z0Z_22 ));
    InMux I__6680 (
            .O(N__43677),
            .I(N__43674));
    LocalMux I__6679 (
            .O(N__43674),
            .I(N__43671));
    Odrv4 I__6678 (
            .O(N__43671),
            .I(\pid_front.pid_preregZ0Z_26 ));
    InMux I__6677 (
            .O(N__43668),
            .I(\pid_front.un1_pid_prereg_0_cry_25 ));
    InMux I__6676 (
            .O(N__43665),
            .I(N__43662));
    LocalMux I__6675 (
            .O(N__43662),
            .I(\pid_front.error_d_reg_prev_esr_RNISQ6O8Z0Z_22 ));
    CascadeMux I__6674 (
            .O(N__43659),
            .I(N__43656));
    InMux I__6673 (
            .O(N__43656),
            .I(N__43653));
    LocalMux I__6672 (
            .O(N__43653),
            .I(\pid_front.error_d_reg_prev_esr_RNICA2C4Z0Z_22 ));
    CascadeMux I__6671 (
            .O(N__43650),
            .I(N__43647));
    InMux I__6670 (
            .O(N__43647),
            .I(N__43644));
    LocalMux I__6669 (
            .O(N__43644),
            .I(N__43641));
    Odrv4 I__6668 (
            .O(N__43641),
            .I(\pid_front.pid_preregZ0Z_27 ));
    InMux I__6667 (
            .O(N__43638),
            .I(\pid_front.un1_pid_prereg_0_cry_26 ));
    InMux I__6666 (
            .O(N__43635),
            .I(N__43632));
    LocalMux I__6665 (
            .O(N__43632),
            .I(\pid_front.error_d_reg_prev_esr_RNI36BO8Z0Z_22 ));
    CascadeMux I__6664 (
            .O(N__43629),
            .I(N__43626));
    InMux I__6663 (
            .O(N__43626),
            .I(N__43623));
    LocalMux I__6662 (
            .O(N__43623),
            .I(\pid_front.error_d_reg_prev_esr_RNIGG4C4Z0Z_22 ));
    InMux I__6661 (
            .O(N__43620),
            .I(N__43617));
    LocalMux I__6660 (
            .O(N__43617),
            .I(N__43614));
    Odrv12 I__6659 (
            .O(N__43614),
            .I(\pid_front.pid_preregZ0Z_28 ));
    InMux I__6658 (
            .O(N__43611),
            .I(\pid_front.un1_pid_prereg_0_cry_27 ));
    InMux I__6657 (
            .O(N__43608),
            .I(N__43605));
    LocalMux I__6656 (
            .O(N__43605),
            .I(\pid_front.error_d_reg_prev_esr_RNI7DEO8Z0Z_22 ));
    CascadeMux I__6655 (
            .O(N__43602),
            .I(N__43599));
    InMux I__6654 (
            .O(N__43599),
            .I(N__43596));
    LocalMux I__6653 (
            .O(N__43596),
            .I(\pid_front.error_d_reg_prev_esr_RNIJL6C4Z0Z_22 ));
    InMux I__6652 (
            .O(N__43593),
            .I(N__43590));
    LocalMux I__6651 (
            .O(N__43590),
            .I(N__43587));
    Span4Mux_v I__6650 (
            .O(N__43587),
            .I(N__43584));
    Odrv4 I__6649 (
            .O(N__43584),
            .I(\pid_front.pid_preregZ0Z_29 ));
    InMux I__6648 (
            .O(N__43581),
            .I(\pid_front.un1_pid_prereg_0_cry_28 ));
    InMux I__6647 (
            .O(N__43578),
            .I(N__43575));
    LocalMux I__6646 (
            .O(N__43575),
            .I(\pid_front.un1_pid_prereg_0_axb_30 ));
    InMux I__6645 (
            .O(N__43572),
            .I(\pid_front.un1_pid_prereg_0_cry_29 ));
    CascadeMux I__6644 (
            .O(N__43569),
            .I(\pid_front.un1_pid_prereg_0_17_cascade_ ));
    CascadeMux I__6643 (
            .O(N__43566),
            .I(N__43563));
    InMux I__6642 (
            .O(N__43563),
            .I(N__43560));
    LocalMux I__6641 (
            .O(N__43560),
            .I(\pid_front.error_d_reg_prev_esr_RNI4UTB4Z0Z_22 ));
    CascadeMux I__6640 (
            .O(N__43557),
            .I(N__43554));
    InMux I__6639 (
            .O(N__43554),
            .I(N__43551));
    LocalMux I__6638 (
            .O(N__43551),
            .I(N__43548));
    Span4Mux_h I__6637 (
            .O(N__43548),
            .I(N__43545));
    Odrv4 I__6636 (
            .O(N__43545),
            .I(\pid_front.pid_preregZ0Z_17 ));
    InMux I__6635 (
            .O(N__43542),
            .I(\pid_front.un1_pid_prereg_0_cry_16 ));
    InMux I__6634 (
            .O(N__43539),
            .I(N__43536));
    LocalMux I__6633 (
            .O(N__43536),
            .I(N__43533));
    Odrv4 I__6632 (
            .O(N__43533),
            .I(\pid_front.pid_preregZ0Z_18 ));
    InMux I__6631 (
            .O(N__43530),
            .I(\pid_front.un1_pid_prereg_0_cry_17 ));
    InMux I__6630 (
            .O(N__43527),
            .I(N__43524));
    LocalMux I__6629 (
            .O(N__43524),
            .I(N__43521));
    Odrv4 I__6628 (
            .O(N__43521),
            .I(\pid_front.pid_preregZ0Z_19 ));
    InMux I__6627 (
            .O(N__43518),
            .I(\pid_front.un1_pid_prereg_0_cry_18 ));
    InMux I__6626 (
            .O(N__43515),
            .I(N__43512));
    LocalMux I__6625 (
            .O(N__43512),
            .I(\pid_front.error_p_reg_esr_RNI80EDDZ0Z_17 ));
    InMux I__6624 (
            .O(N__43509),
            .I(N__43506));
    LocalMux I__6623 (
            .O(N__43506),
            .I(\pid_front.pid_preregZ0Z_20 ));
    InMux I__6622 (
            .O(N__43503),
            .I(\pid_front.un1_pid_prereg_0_cry_19 ));
    InMux I__6621 (
            .O(N__43500),
            .I(N__43497));
    LocalMux I__6620 (
            .O(N__43497),
            .I(\pid_front.error_p_reg_esr_RNISOJEDZ0Z_18 ));
    CascadeMux I__6619 (
            .O(N__43494),
            .I(N__43491));
    InMux I__6618 (
            .O(N__43491),
            .I(N__43488));
    LocalMux I__6617 (
            .O(N__43488),
            .I(\pid_front.error_p_reg_esr_RNIQOPM6Z0Z_18 ));
    InMux I__6616 (
            .O(N__43485),
            .I(N__43482));
    LocalMux I__6615 (
            .O(N__43482),
            .I(\pid_front.pid_preregZ0Z_21 ));
    InMux I__6614 (
            .O(N__43479),
            .I(\pid_front.un1_pid_prereg_0_cry_20 ));
    CascadeMux I__6613 (
            .O(N__43476),
            .I(N__43473));
    InMux I__6612 (
            .O(N__43473),
            .I(N__43470));
    LocalMux I__6611 (
            .O(N__43470),
            .I(\pid_front.error_p_reg_esr_RNI20QN6Z0Z_19 ));
    InMux I__6610 (
            .O(N__43467),
            .I(N__43464));
    LocalMux I__6609 (
            .O(N__43464),
            .I(\pid_front.pid_preregZ0Z_22 ));
    InMux I__6608 (
            .O(N__43461),
            .I(\pid_front.un1_pid_prereg_0_cry_21 ));
    CascadeMux I__6607 (
            .O(N__43458),
            .I(N__43455));
    InMux I__6606 (
            .O(N__43455),
            .I(N__43452));
    LocalMux I__6605 (
            .O(N__43452),
            .I(N__43449));
    Odrv4 I__6604 (
            .O(N__43449),
            .I(\pid_front.pid_preregZ0Z_23 ));
    InMux I__6603 (
            .O(N__43446),
            .I(bfn_9_20_0_));
    InMux I__6602 (
            .O(N__43443),
            .I(N__43440));
    LocalMux I__6601 (
            .O(N__43440),
            .I(N__43437));
    Odrv4 I__6600 (
            .O(N__43437),
            .I(\pid_front.pid_preregZ0Z_24 ));
    InMux I__6599 (
            .O(N__43434),
            .I(\pid_front.un1_pid_prereg_0_cry_23 ));
    InMux I__6598 (
            .O(N__43431),
            .I(N__43428));
    LocalMux I__6597 (
            .O(N__43428),
            .I(\pid_front.error_p_reg_esr_RNIV7CQ2Z0Z_8 ));
    InMux I__6596 (
            .O(N__43425),
            .I(N__43421));
    InMux I__6595 (
            .O(N__43424),
            .I(N__43418));
    LocalMux I__6594 (
            .O(N__43421),
            .I(N__43415));
    LocalMux I__6593 (
            .O(N__43418),
            .I(N__43411));
    Span4Mux_v I__6592 (
            .O(N__43415),
            .I(N__43408));
    InMux I__6591 (
            .O(N__43414),
            .I(N__43405));
    Odrv12 I__6590 (
            .O(N__43411),
            .I(\pid_front.pid_preregZ0Z_9 ));
    Odrv4 I__6589 (
            .O(N__43408),
            .I(\pid_front.pid_preregZ0Z_9 ));
    LocalMux I__6588 (
            .O(N__43405),
            .I(\pid_front.pid_preregZ0Z_9 ));
    InMux I__6587 (
            .O(N__43398),
            .I(\pid_front.un1_pid_prereg_0_cry_8 ));
    InMux I__6586 (
            .O(N__43395),
            .I(\pid_front.un1_pid_prereg_0_cry_9 ));
    InMux I__6585 (
            .O(N__43392),
            .I(\pid_front.un1_pid_prereg_0_cry_10 ));
    InMux I__6584 (
            .O(N__43389),
            .I(\pid_front.un1_pid_prereg_0_cry_11 ));
    InMux I__6583 (
            .O(N__43386),
            .I(\pid_front.un1_pid_prereg_0_cry_12 ));
    InMux I__6582 (
            .O(N__43383),
            .I(N__43380));
    LocalMux I__6581 (
            .O(N__43380),
            .I(\pid_front.un1_pid_prereg_0_cry_13_THRU_CO ));
    InMux I__6580 (
            .O(N__43377),
            .I(\pid_front.un1_pid_prereg_0_cry_13 ));
    CascadeMux I__6579 (
            .O(N__43374),
            .I(N__43371));
    InMux I__6578 (
            .O(N__43371),
            .I(N__43367));
    InMux I__6577 (
            .O(N__43370),
            .I(N__43364));
    LocalMux I__6576 (
            .O(N__43367),
            .I(N__43359));
    LocalMux I__6575 (
            .O(N__43364),
            .I(N__43359));
    Odrv4 I__6574 (
            .O(N__43359),
            .I(\pid_front.pid_preregZ0Z_15 ));
    InMux I__6573 (
            .O(N__43356),
            .I(bfn_9_19_0_));
    InMux I__6572 (
            .O(N__43353),
            .I(N__43350));
    LocalMux I__6571 (
            .O(N__43350),
            .I(N__43347));
    Odrv4 I__6570 (
            .O(N__43347),
            .I(\pid_front.pid_preregZ0Z_16 ));
    InMux I__6569 (
            .O(N__43344),
            .I(\pid_front.un1_pid_prereg_0_cry_15 ));
    InMux I__6568 (
            .O(N__43341),
            .I(N__43338));
    LocalMux I__6567 (
            .O(N__43338),
            .I(N__43333));
    InMux I__6566 (
            .O(N__43337),
            .I(N__43330));
    InMux I__6565 (
            .O(N__43336),
            .I(N__43327));
    Odrv4 I__6564 (
            .O(N__43333),
            .I(\pid_front.pid_preregZ0Z_0 ));
    LocalMux I__6563 (
            .O(N__43330),
            .I(\pid_front.pid_preregZ0Z_0 ));
    LocalMux I__6562 (
            .O(N__43327),
            .I(\pid_front.pid_preregZ0Z_0 ));
    InMux I__6561 (
            .O(N__43320),
            .I(\pid_front.un1_pid_prereg_0_cry_0_c_THRU_CO ));
    InMux I__6560 (
            .O(N__43317),
            .I(N__43314));
    LocalMux I__6559 (
            .O(N__43314),
            .I(N__43309));
    InMux I__6558 (
            .O(N__43313),
            .I(N__43304));
    InMux I__6557 (
            .O(N__43312),
            .I(N__43304));
    Odrv4 I__6556 (
            .O(N__43309),
            .I(\pid_front.pid_preregZ0Z_1 ));
    LocalMux I__6555 (
            .O(N__43304),
            .I(\pid_front.pid_preregZ0Z_1 ));
    InMux I__6554 (
            .O(N__43299),
            .I(\pid_front.un1_pid_prereg_0_cry_0 ));
    InMux I__6553 (
            .O(N__43296),
            .I(N__43287));
    InMux I__6552 (
            .O(N__43295),
            .I(N__43287));
    InMux I__6551 (
            .O(N__43294),
            .I(N__43287));
    LocalMux I__6550 (
            .O(N__43287),
            .I(\pid_front.pid_preregZ0Z_2 ));
    InMux I__6549 (
            .O(N__43284),
            .I(\pid_front.un1_pid_prereg_0_cry_1 ));
    CascadeMux I__6548 (
            .O(N__43281),
            .I(N__43277));
    CascadeMux I__6547 (
            .O(N__43280),
            .I(N__43273));
    InMux I__6546 (
            .O(N__43277),
            .I(N__43270));
    InMux I__6545 (
            .O(N__43276),
            .I(N__43265));
    InMux I__6544 (
            .O(N__43273),
            .I(N__43265));
    LocalMux I__6543 (
            .O(N__43270),
            .I(\pid_front.pid_preregZ0Z_3 ));
    LocalMux I__6542 (
            .O(N__43265),
            .I(\pid_front.pid_preregZ0Z_3 ));
    InMux I__6541 (
            .O(N__43260),
            .I(\pid_front.un1_pid_prereg_0_cry_2 ));
    InMux I__6540 (
            .O(N__43257),
            .I(N__43253));
    InMux I__6539 (
            .O(N__43256),
            .I(N__43250));
    LocalMux I__6538 (
            .O(N__43253),
            .I(N__43247));
    LocalMux I__6537 (
            .O(N__43250),
            .I(N__43244));
    Span4Mux_v I__6536 (
            .O(N__43247),
            .I(N__43237));
    Span4Mux_h I__6535 (
            .O(N__43244),
            .I(N__43237));
    InMux I__6534 (
            .O(N__43243),
            .I(N__43232));
    InMux I__6533 (
            .O(N__43242),
            .I(N__43232));
    Odrv4 I__6532 (
            .O(N__43237),
            .I(\pid_front.pid_preregZ0Z_4 ));
    LocalMux I__6531 (
            .O(N__43232),
            .I(\pid_front.pid_preregZ0Z_4 ));
    InMux I__6530 (
            .O(N__43227),
            .I(\pid_front.un1_pid_prereg_0_cry_3 ));
    InMux I__6529 (
            .O(N__43224),
            .I(N__43220));
    InMux I__6528 (
            .O(N__43223),
            .I(N__43217));
    LocalMux I__6527 (
            .O(N__43220),
            .I(N__43213));
    LocalMux I__6526 (
            .O(N__43217),
            .I(N__43209));
    InMux I__6525 (
            .O(N__43216),
            .I(N__43206));
    Span4Mux_h I__6524 (
            .O(N__43213),
            .I(N__43203));
    InMux I__6523 (
            .O(N__43212),
            .I(N__43200));
    Odrv4 I__6522 (
            .O(N__43209),
            .I(\pid_front.pid_preregZ0Z_5 ));
    LocalMux I__6521 (
            .O(N__43206),
            .I(\pid_front.pid_preregZ0Z_5 ));
    Odrv4 I__6520 (
            .O(N__43203),
            .I(\pid_front.pid_preregZ0Z_5 ));
    LocalMux I__6519 (
            .O(N__43200),
            .I(\pid_front.pid_preregZ0Z_5 ));
    InMux I__6518 (
            .O(N__43191),
            .I(\pid_front.un1_pid_prereg_0_cry_4 ));
    CascadeMux I__6517 (
            .O(N__43188),
            .I(N__43183));
    InMux I__6516 (
            .O(N__43187),
            .I(N__43180));
    InMux I__6515 (
            .O(N__43186),
            .I(N__43177));
    InMux I__6514 (
            .O(N__43183),
            .I(N__43174));
    LocalMux I__6513 (
            .O(N__43180),
            .I(N__43171));
    LocalMux I__6512 (
            .O(N__43177),
            .I(N__43166));
    LocalMux I__6511 (
            .O(N__43174),
            .I(N__43166));
    Odrv12 I__6510 (
            .O(N__43171),
            .I(\pid_front.pid_preregZ0Z_6 ));
    Odrv4 I__6509 (
            .O(N__43166),
            .I(\pid_front.pid_preregZ0Z_6 ));
    InMux I__6508 (
            .O(N__43161),
            .I(\pid_front.un1_pid_prereg_0_cry_5 ));
    InMux I__6507 (
            .O(N__43158),
            .I(N__43153));
    InMux I__6506 (
            .O(N__43157),
            .I(N__43148));
    InMux I__6505 (
            .O(N__43156),
            .I(N__43148));
    LocalMux I__6504 (
            .O(N__43153),
            .I(N__43145));
    LocalMux I__6503 (
            .O(N__43148),
            .I(N__43142));
    Odrv12 I__6502 (
            .O(N__43145),
            .I(\pid_front.pid_preregZ0Z_7 ));
    Odrv4 I__6501 (
            .O(N__43142),
            .I(\pid_front.pid_preregZ0Z_7 ));
    InMux I__6500 (
            .O(N__43137),
            .I(bfn_9_18_0_));
    InMux I__6499 (
            .O(N__43134),
            .I(\pid_front.un1_pid_prereg_0_cry_7 ));
    InMux I__6498 (
            .O(N__43131),
            .I(N__43128));
    LocalMux I__6497 (
            .O(N__43128),
            .I(N__43124));
    InMux I__6496 (
            .O(N__43127),
            .I(N__43121));
    Span4Mux_h I__6495 (
            .O(N__43124),
            .I(N__43116));
    LocalMux I__6494 (
            .O(N__43121),
            .I(N__43116));
    Odrv4 I__6493 (
            .O(N__43116),
            .I(\pid_front.N_99 ));
    InMux I__6492 (
            .O(N__43113),
            .I(N__43110));
    LocalMux I__6491 (
            .O(N__43110),
            .I(N__43107));
    Odrv4 I__6490 (
            .O(N__43107),
            .I(\pid_front.source_pid_1_sqmuxa_1_0_a4_4 ));
    InMux I__6489 (
            .O(N__43104),
            .I(N__43101));
    LocalMux I__6488 (
            .O(N__43101),
            .I(\pid_front.source_pid10lt4_0 ));
    InMux I__6487 (
            .O(N__43098),
            .I(N__43084));
    InMux I__6486 (
            .O(N__43097),
            .I(N__43084));
    InMux I__6485 (
            .O(N__43096),
            .I(N__43084));
    InMux I__6484 (
            .O(N__43095),
            .I(N__43084));
    InMux I__6483 (
            .O(N__43094),
            .I(N__43079));
    InMux I__6482 (
            .O(N__43093),
            .I(N__43079));
    LocalMux I__6481 (
            .O(N__43084),
            .I(N__43076));
    LocalMux I__6480 (
            .O(N__43079),
            .I(N__43073));
    Span4Mux_h I__6479 (
            .O(N__43076),
            .I(N__43070));
    Odrv4 I__6478 (
            .O(N__43073),
            .I(\pid_front.N_75 ));
    Odrv4 I__6477 (
            .O(N__43070),
            .I(\pid_front.N_75 ));
    CascadeMux I__6476 (
            .O(N__43065),
            .I(N__43060));
    InMux I__6475 (
            .O(N__43064),
            .I(N__43057));
    InMux I__6474 (
            .O(N__43063),
            .I(N__43052));
    InMux I__6473 (
            .O(N__43060),
            .I(N__43052));
    LocalMux I__6472 (
            .O(N__43057),
            .I(\dron_frame_decoder_1.WDTZ0Z_14 ));
    LocalMux I__6471 (
            .O(N__43052),
            .I(\dron_frame_decoder_1.WDTZ0Z_14 ));
    InMux I__6470 (
            .O(N__43047),
            .I(N__43042));
    InMux I__6469 (
            .O(N__43046),
            .I(N__43039));
    InMux I__6468 (
            .O(N__43045),
            .I(N__43036));
    LocalMux I__6467 (
            .O(N__43042),
            .I(\dron_frame_decoder_1.WDTZ0Z_15 ));
    LocalMux I__6466 (
            .O(N__43039),
            .I(\dron_frame_decoder_1.WDTZ0Z_15 ));
    LocalMux I__6465 (
            .O(N__43036),
            .I(\dron_frame_decoder_1.WDTZ0Z_15 ));
    CascadeMux I__6464 (
            .O(N__43029),
            .I(\dron_frame_decoder_1.WDT10lt14_0_cascade_ ));
    CascadeMux I__6463 (
            .O(N__43026),
            .I(\dron_frame_decoder_1.N_218_cascade_ ));
    InMux I__6462 (
            .O(N__43023),
            .I(N__43020));
    LocalMux I__6461 (
            .O(N__43020),
            .I(N__43017));
    Span4Mux_v I__6460 (
            .O(N__43017),
            .I(N__43013));
    InMux I__6459 (
            .O(N__43016),
            .I(N__43010));
    Odrv4 I__6458 (
            .O(N__43013),
            .I(\pid_front.un11lto30_i_a2_6_and ));
    LocalMux I__6457 (
            .O(N__43010),
            .I(\pid_front.un11lto30_i_a2_6_and ));
    InMux I__6456 (
            .O(N__43005),
            .I(N__43002));
    LocalMux I__6455 (
            .O(N__43002),
            .I(\pid_front.source_pid_1_sqmuxa_1_0_o2_sx ));
    InMux I__6454 (
            .O(N__42999),
            .I(N__42996));
    LocalMux I__6453 (
            .O(N__42996),
            .I(N__42993));
    Odrv4 I__6452 (
            .O(N__42993),
            .I(\pid_front.N_389 ));
    CascadeMux I__6451 (
            .O(N__42990),
            .I(\pid_front.N_102_cascade_ ));
    CascadeMux I__6450 (
            .O(N__42987),
            .I(\pid_front.un1_reset_0_i_cascade_ ));
    CascadeMux I__6449 (
            .O(N__42984),
            .I(N__42981));
    InMux I__6448 (
            .O(N__42981),
            .I(N__42975));
    InMux I__6447 (
            .O(N__42980),
            .I(N__42975));
    LocalMux I__6446 (
            .O(N__42975),
            .I(N__42972));
    Odrv12 I__6445 (
            .O(N__42972),
            .I(\scaler_4.un3_source_data_0_cry_6_c_RNIOUNN ));
    InMux I__6444 (
            .O(N__42969),
            .I(\scaler_4.un3_source_data_0_cry_6 ));
    InMux I__6443 (
            .O(N__42966),
            .I(N__42962));
    InMux I__6442 (
            .O(N__42965),
            .I(N__42959));
    LocalMux I__6441 (
            .O(N__42962),
            .I(N__42956));
    LocalMux I__6440 (
            .O(N__42959),
            .I(N__42953));
    Odrv4 I__6439 (
            .O(N__42956),
            .I(\scaler_4.un3_source_data_0_cry_7_c_RNIP0PN ));
    Odrv12 I__6438 (
            .O(N__42953),
            .I(\scaler_4.un3_source_data_0_cry_7_c_RNIP0PN ));
    InMux I__6437 (
            .O(N__42948),
            .I(bfn_9_12_0_));
    InMux I__6436 (
            .O(N__42945),
            .I(\scaler_4.un3_source_data_0_cry_8 ));
    CascadeMux I__6435 (
            .O(N__42942),
            .I(N__42939));
    InMux I__6434 (
            .O(N__42939),
            .I(N__42936));
    LocalMux I__6433 (
            .O(N__42936),
            .I(N__42933));
    Odrv4 I__6432 (
            .O(N__42933),
            .I(\scaler_4.un3_source_data_0_cry_8_c_RNIS918 ));
    InMux I__6431 (
            .O(N__42930),
            .I(N__42926));
    InMux I__6430 (
            .O(N__42929),
            .I(N__42923));
    LocalMux I__6429 (
            .O(N__42926),
            .I(N__42920));
    LocalMux I__6428 (
            .O(N__42923),
            .I(\dron_frame_decoder_1.WDTZ0Z_8 ));
    Odrv4 I__6427 (
            .O(N__42920),
            .I(\dron_frame_decoder_1.WDTZ0Z_8 ));
    InMux I__6426 (
            .O(N__42915),
            .I(N__42911));
    InMux I__6425 (
            .O(N__42914),
            .I(N__42908));
    LocalMux I__6424 (
            .O(N__42911),
            .I(\dron_frame_decoder_1.WDTZ0Z_5 ));
    LocalMux I__6423 (
            .O(N__42908),
            .I(\dron_frame_decoder_1.WDTZ0Z_5 ));
    CascadeMux I__6422 (
            .O(N__42903),
            .I(N__42899));
    InMux I__6421 (
            .O(N__42902),
            .I(N__42896));
    InMux I__6420 (
            .O(N__42899),
            .I(N__42893));
    LocalMux I__6419 (
            .O(N__42896),
            .I(\dron_frame_decoder_1.WDTZ0Z_9 ));
    LocalMux I__6418 (
            .O(N__42893),
            .I(\dron_frame_decoder_1.WDTZ0Z_9 ));
    InMux I__6417 (
            .O(N__42888),
            .I(N__42884));
    InMux I__6416 (
            .O(N__42887),
            .I(N__42881));
    LocalMux I__6415 (
            .O(N__42884),
            .I(\dron_frame_decoder_1.WDTZ0Z_4 ));
    LocalMux I__6414 (
            .O(N__42881),
            .I(\dron_frame_decoder_1.WDTZ0Z_4 ));
    CascadeMux I__6413 (
            .O(N__42876),
            .I(\dron_frame_decoder_1.WDT10_0_i_1_cascade_ ));
    CascadeMux I__6412 (
            .O(N__42873),
            .I(N__42869));
    InMux I__6411 (
            .O(N__42872),
            .I(N__42866));
    InMux I__6410 (
            .O(N__42869),
            .I(N__42863));
    LocalMux I__6409 (
            .O(N__42866),
            .I(\dron_frame_decoder_1.WDT10_0_i ));
    LocalMux I__6408 (
            .O(N__42863),
            .I(\dron_frame_decoder_1.WDT10_0_i ));
    InMux I__6407 (
            .O(N__42858),
            .I(N__42854));
    InMux I__6406 (
            .O(N__42857),
            .I(N__42851));
    LocalMux I__6405 (
            .O(N__42854),
            .I(\dron_frame_decoder_1.WDTZ0Z_6 ));
    LocalMux I__6404 (
            .O(N__42851),
            .I(\dron_frame_decoder_1.WDTZ0Z_6 ));
    InMux I__6403 (
            .O(N__42846),
            .I(N__42842));
    InMux I__6402 (
            .O(N__42845),
            .I(N__42839));
    LocalMux I__6401 (
            .O(N__42842),
            .I(\dron_frame_decoder_1.WDTZ0Z_7 ));
    LocalMux I__6400 (
            .O(N__42839),
            .I(\dron_frame_decoder_1.WDTZ0Z_7 ));
    CascadeMux I__6399 (
            .O(N__42834),
            .I(N__42830));
    InMux I__6398 (
            .O(N__42833),
            .I(N__42827));
    InMux I__6397 (
            .O(N__42830),
            .I(N__42824));
    LocalMux I__6396 (
            .O(N__42827),
            .I(\dron_frame_decoder_1.WDTZ0Z_10 ));
    LocalMux I__6395 (
            .O(N__42824),
            .I(\dron_frame_decoder_1.WDTZ0Z_10 ));
    InMux I__6394 (
            .O(N__42819),
            .I(N__42816));
    LocalMux I__6393 (
            .O(N__42816),
            .I(\dron_frame_decoder_1.WDT10lto9_3 ));
    InMux I__6392 (
            .O(N__42813),
            .I(N__42810));
    LocalMux I__6391 (
            .O(N__42810),
            .I(\dron_frame_decoder_1.WDT10lt12_0 ));
    InMux I__6390 (
            .O(N__42807),
            .I(N__42802));
    InMux I__6389 (
            .O(N__42806),
            .I(N__42797));
    InMux I__6388 (
            .O(N__42805),
            .I(N__42797));
    LocalMux I__6387 (
            .O(N__42802),
            .I(\dron_frame_decoder_1.WDTZ0Z_11 ));
    LocalMux I__6386 (
            .O(N__42797),
            .I(\dron_frame_decoder_1.WDTZ0Z_11 ));
    InMux I__6385 (
            .O(N__42792),
            .I(N__42786));
    InMux I__6384 (
            .O(N__42791),
            .I(N__42783));
    InMux I__6383 (
            .O(N__42790),
            .I(N__42778));
    InMux I__6382 (
            .O(N__42789),
            .I(N__42778));
    LocalMux I__6381 (
            .O(N__42786),
            .I(\dron_frame_decoder_1.WDTZ0Z_13 ));
    LocalMux I__6380 (
            .O(N__42783),
            .I(\dron_frame_decoder_1.WDTZ0Z_13 ));
    LocalMux I__6379 (
            .O(N__42778),
            .I(\dron_frame_decoder_1.WDTZ0Z_13 ));
    CascadeMux I__6378 (
            .O(N__42771),
            .I(\dron_frame_decoder_1.WDT10lt12_0_cascade_ ));
    InMux I__6377 (
            .O(N__42768),
            .I(N__42763));
    InMux I__6376 (
            .O(N__42767),
            .I(N__42758));
    InMux I__6375 (
            .O(N__42766),
            .I(N__42758));
    LocalMux I__6374 (
            .O(N__42763),
            .I(\dron_frame_decoder_1.WDTZ0Z_12 ));
    LocalMux I__6373 (
            .O(N__42758),
            .I(\dron_frame_decoder_1.WDTZ0Z_12 ));
    InMux I__6372 (
            .O(N__42753),
            .I(N__42750));
    LocalMux I__6371 (
            .O(N__42750),
            .I(N__42744));
    InMux I__6370 (
            .O(N__42749),
            .I(N__42741));
    InMux I__6369 (
            .O(N__42748),
            .I(N__42738));
    InMux I__6368 (
            .O(N__42747),
            .I(N__42735));
    Odrv12 I__6367 (
            .O(N__42744),
            .I(frame_decoder_CH4data_0));
    LocalMux I__6366 (
            .O(N__42741),
            .I(frame_decoder_CH4data_0));
    LocalMux I__6365 (
            .O(N__42738),
            .I(frame_decoder_CH4data_0));
    LocalMux I__6364 (
            .O(N__42735),
            .I(frame_decoder_CH4data_0));
    InMux I__6363 (
            .O(N__42726),
            .I(N__42723));
    LocalMux I__6362 (
            .O(N__42723),
            .I(N__42718));
    InMux I__6361 (
            .O(N__42722),
            .I(N__42715));
    CascadeMux I__6360 (
            .O(N__42721),
            .I(N__42711));
    Span4Mux_v I__6359 (
            .O(N__42718),
            .I(N__42708));
    LocalMux I__6358 (
            .O(N__42715),
            .I(N__42705));
    InMux I__6357 (
            .O(N__42714),
            .I(N__42702));
    InMux I__6356 (
            .O(N__42711),
            .I(N__42699));
    Odrv4 I__6355 (
            .O(N__42708),
            .I(frame_decoder_OFF4data_0));
    Odrv4 I__6354 (
            .O(N__42705),
            .I(frame_decoder_OFF4data_0));
    LocalMux I__6353 (
            .O(N__42702),
            .I(frame_decoder_OFF4data_0));
    LocalMux I__6352 (
            .O(N__42699),
            .I(frame_decoder_OFF4data_0));
    InMux I__6351 (
            .O(N__42690),
            .I(N__42687));
    LocalMux I__6350 (
            .O(N__42687),
            .I(frame_decoder_CH4data_1));
    CascadeMux I__6349 (
            .O(N__42684),
            .I(N__42681));
    InMux I__6348 (
            .O(N__42681),
            .I(N__42678));
    LocalMux I__6347 (
            .O(N__42678),
            .I(frame_decoder_OFF4data_1));
    InMux I__6346 (
            .O(N__42675),
            .I(N__42670));
    InMux I__6345 (
            .O(N__42674),
            .I(N__42667));
    CascadeMux I__6344 (
            .O(N__42673),
            .I(N__42664));
    LocalMux I__6343 (
            .O(N__42670),
            .I(N__42658));
    LocalMux I__6342 (
            .O(N__42667),
            .I(N__42658));
    InMux I__6341 (
            .O(N__42664),
            .I(N__42653));
    InMux I__6340 (
            .O(N__42663),
            .I(N__42653));
    Span4Mux_h I__6339 (
            .O(N__42658),
            .I(N__42650));
    LocalMux I__6338 (
            .O(N__42653),
            .I(N__42647));
    Odrv4 I__6337 (
            .O(N__42650),
            .I(\scaler_4.un2_source_data_0 ));
    Odrv12 I__6336 (
            .O(N__42647),
            .I(\scaler_4.un2_source_data_0 ));
    InMux I__6335 (
            .O(N__42642),
            .I(\scaler_4.un3_source_data_0_cry_0 ));
    InMux I__6334 (
            .O(N__42639),
            .I(N__42636));
    LocalMux I__6333 (
            .O(N__42636),
            .I(frame_decoder_CH4data_2));
    CascadeMux I__6332 (
            .O(N__42633),
            .I(N__42630));
    InMux I__6331 (
            .O(N__42630),
            .I(N__42627));
    LocalMux I__6330 (
            .O(N__42627),
            .I(frame_decoder_OFF4data_2));
    CascadeMux I__6329 (
            .O(N__42624),
            .I(N__42621));
    InMux I__6328 (
            .O(N__42621),
            .I(N__42615));
    InMux I__6327 (
            .O(N__42620),
            .I(N__42615));
    LocalMux I__6326 (
            .O(N__42615),
            .I(N__42612));
    Odrv4 I__6325 (
            .O(N__42612),
            .I(\scaler_4.un3_source_data_0_cry_1_c_RNI74CL ));
    InMux I__6324 (
            .O(N__42609),
            .I(\scaler_4.un3_source_data_0_cry_1 ));
    InMux I__6323 (
            .O(N__42606),
            .I(N__42603));
    LocalMux I__6322 (
            .O(N__42603),
            .I(frame_decoder_CH4data_3));
    CascadeMux I__6321 (
            .O(N__42600),
            .I(N__42597));
    InMux I__6320 (
            .O(N__42597),
            .I(N__42594));
    LocalMux I__6319 (
            .O(N__42594),
            .I(frame_decoder_OFF4data_3));
    CascadeMux I__6318 (
            .O(N__42591),
            .I(N__42588));
    InMux I__6317 (
            .O(N__42588),
            .I(N__42582));
    InMux I__6316 (
            .O(N__42587),
            .I(N__42582));
    LocalMux I__6315 (
            .O(N__42582),
            .I(N__42579));
    Odrv4 I__6314 (
            .O(N__42579),
            .I(\scaler_4.un3_source_data_0_cry_2_c_RNIA8DL ));
    InMux I__6313 (
            .O(N__42576),
            .I(\scaler_4.un3_source_data_0_cry_2 ));
    InMux I__6312 (
            .O(N__42573),
            .I(N__42570));
    LocalMux I__6311 (
            .O(N__42570),
            .I(frame_decoder_CH4data_4));
    CascadeMux I__6310 (
            .O(N__42567),
            .I(N__42564));
    InMux I__6309 (
            .O(N__42564),
            .I(N__42561));
    LocalMux I__6308 (
            .O(N__42561),
            .I(frame_decoder_OFF4data_4));
    CascadeMux I__6307 (
            .O(N__42558),
            .I(N__42555));
    InMux I__6306 (
            .O(N__42555),
            .I(N__42549));
    InMux I__6305 (
            .O(N__42554),
            .I(N__42549));
    LocalMux I__6304 (
            .O(N__42549),
            .I(N__42546));
    Odrv4 I__6303 (
            .O(N__42546),
            .I(\scaler_4.un3_source_data_0_cry_3_c_RNIDCEL ));
    InMux I__6302 (
            .O(N__42543),
            .I(\scaler_4.un3_source_data_0_cry_3 ));
    InMux I__6301 (
            .O(N__42540),
            .I(N__42537));
    LocalMux I__6300 (
            .O(N__42537),
            .I(frame_decoder_CH4data_5));
    CascadeMux I__6299 (
            .O(N__42534),
            .I(N__42531));
    InMux I__6298 (
            .O(N__42531),
            .I(N__42528));
    LocalMux I__6297 (
            .O(N__42528),
            .I(frame_decoder_OFF4data_5));
    CascadeMux I__6296 (
            .O(N__42525),
            .I(N__42522));
    InMux I__6295 (
            .O(N__42522),
            .I(N__42516));
    InMux I__6294 (
            .O(N__42521),
            .I(N__42516));
    LocalMux I__6293 (
            .O(N__42516),
            .I(N__42513));
    Odrv4 I__6292 (
            .O(N__42513),
            .I(\scaler_4.un3_source_data_0_cry_4_c_RNIGGFL ));
    InMux I__6291 (
            .O(N__42510),
            .I(\scaler_4.un3_source_data_0_cry_4 ));
    InMux I__6290 (
            .O(N__42507),
            .I(N__42504));
    LocalMux I__6289 (
            .O(N__42504),
            .I(frame_decoder_CH4data_6));
    CascadeMux I__6288 (
            .O(N__42501),
            .I(N__42498));
    InMux I__6287 (
            .O(N__42498),
            .I(N__42495));
    LocalMux I__6286 (
            .O(N__42495),
            .I(frame_decoder_OFF4data_6));
    CascadeMux I__6285 (
            .O(N__42492),
            .I(N__42489));
    InMux I__6284 (
            .O(N__42489),
            .I(N__42483));
    InMux I__6283 (
            .O(N__42488),
            .I(N__42483));
    LocalMux I__6282 (
            .O(N__42483),
            .I(N__42480));
    Odrv12 I__6281 (
            .O(N__42480),
            .I(\scaler_4.un3_source_data_0_cry_5_c_RNIJKGL ));
    InMux I__6280 (
            .O(N__42477),
            .I(\scaler_4.un3_source_data_0_cry_5 ));
    InMux I__6279 (
            .O(N__42474),
            .I(N__42471));
    LocalMux I__6278 (
            .O(N__42471),
            .I(N__42468));
    Span4Mux_h I__6277 (
            .O(N__42468),
            .I(N__42465));
    Span4Mux_v I__6276 (
            .O(N__42465),
            .I(N__42462));
    Odrv4 I__6275 (
            .O(N__42462),
            .I(\scaler_4.un3_source_data_0_axb_7 ));
    InMux I__6274 (
            .O(N__42459),
            .I(\scaler_4.un2_source_data_0_cry_2 ));
    InMux I__6273 (
            .O(N__42456),
            .I(\scaler_4.un2_source_data_0_cry_3 ));
    InMux I__6272 (
            .O(N__42453),
            .I(\scaler_4.un2_source_data_0_cry_4 ));
    InMux I__6271 (
            .O(N__42450),
            .I(\scaler_4.un2_source_data_0_cry_5 ));
    InMux I__6270 (
            .O(N__42447),
            .I(\scaler_4.un2_source_data_0_cry_6 ));
    InMux I__6269 (
            .O(N__42444),
            .I(\scaler_4.un2_source_data_0_cry_7 ));
    InMux I__6268 (
            .O(N__42441),
            .I(bfn_9_9_0_));
    InMux I__6267 (
            .O(N__42438),
            .I(\scaler_4.un2_source_data_0_cry_9 ));
    InMux I__6266 (
            .O(N__42435),
            .I(N__42432));
    LocalMux I__6265 (
            .O(N__42432),
            .I(N__42429));
    Odrv4 I__6264 (
            .O(N__42429),
            .I(scaler_4_data_14));
    CEMux I__6263 (
            .O(N__42426),
            .I(N__42422));
    CEMux I__6262 (
            .O(N__42425),
            .I(N__42418));
    LocalMux I__6261 (
            .O(N__42422),
            .I(N__42415));
    CEMux I__6260 (
            .O(N__42421),
            .I(N__42412));
    LocalMux I__6259 (
            .O(N__42418),
            .I(N__42409));
    Span4Mux_v I__6258 (
            .O(N__42415),
            .I(N__42406));
    LocalMux I__6257 (
            .O(N__42412),
            .I(N__42403));
    Span4Mux_v I__6256 (
            .O(N__42409),
            .I(N__42396));
    Span4Mux_h I__6255 (
            .O(N__42406),
            .I(N__42396));
    Span4Mux_v I__6254 (
            .O(N__42403),
            .I(N__42396));
    Odrv4 I__6253 (
            .O(N__42396),
            .I(\scaler_4.debug_CH3_20A_c_0 ));
    InMux I__6252 (
            .O(N__42393),
            .I(\ppm_encoder_1.un1_rudder_cry_7 ));
    InMux I__6251 (
            .O(N__42390),
            .I(\ppm_encoder_1.un1_rudder_cry_8 ));
    InMux I__6250 (
            .O(N__42387),
            .I(\ppm_encoder_1.un1_rudder_cry_9 ));
    InMux I__6249 (
            .O(N__42384),
            .I(\ppm_encoder_1.un1_rudder_cry_10 ));
    InMux I__6248 (
            .O(N__42381),
            .I(\ppm_encoder_1.un1_rudder_cry_11 ));
    InMux I__6247 (
            .O(N__42378),
            .I(\ppm_encoder_1.un1_rudder_cry_12 ));
    InMux I__6246 (
            .O(N__42375),
            .I(bfn_9_7_0_));
    CascadeMux I__6245 (
            .O(N__42372),
            .I(N__42369));
    InMux I__6244 (
            .O(N__42369),
            .I(N__42366));
    LocalMux I__6243 (
            .O(N__42366),
            .I(N__42363));
    Span4Mux_h I__6242 (
            .O(N__42363),
            .I(N__42360));
    Odrv4 I__6241 (
            .O(N__42360),
            .I(\scaler_4.un2_source_data_0_cry_1_c_RNOZ0 ));
    InMux I__6240 (
            .O(N__42357),
            .I(N__42353));
    InMux I__6239 (
            .O(N__42356),
            .I(N__42350));
    LocalMux I__6238 (
            .O(N__42353),
            .I(N__42347));
    LocalMux I__6237 (
            .O(N__42350),
            .I(N__42344));
    Odrv4 I__6236 (
            .O(N__42347),
            .I(scaler_4_data_6));
    Odrv4 I__6235 (
            .O(N__42344),
            .I(scaler_4_data_6));
    InMux I__6234 (
            .O(N__42339),
            .I(\scaler_4.un2_source_data_0_cry_1 ));
    CascadeMux I__6233 (
            .O(N__42336),
            .I(N__42333));
    InMux I__6232 (
            .O(N__42333),
            .I(N__42330));
    LocalMux I__6231 (
            .O(N__42330),
            .I(\ppm_encoder_1.un2_throttle_iv_0_1_4 ));
    InMux I__6230 (
            .O(N__42327),
            .I(N__42324));
    LocalMux I__6229 (
            .O(N__42324),
            .I(N__42321));
    Span4Mux_v I__6228 (
            .O(N__42321),
            .I(N__42318));
    Odrv4 I__6227 (
            .O(N__42318),
            .I(\ppm_encoder_1.un1_throttle_cry_3_THRU_CO ));
    InMux I__6226 (
            .O(N__42315),
            .I(N__42311));
    InMux I__6225 (
            .O(N__42314),
            .I(N__42308));
    LocalMux I__6224 (
            .O(N__42311),
            .I(N__42305));
    LocalMux I__6223 (
            .O(N__42308),
            .I(N__42302));
    Span4Mux_v I__6222 (
            .O(N__42305),
            .I(N__42299));
    Span12Mux_h I__6221 (
            .O(N__42302),
            .I(N__42296));
    Span4Mux_h I__6220 (
            .O(N__42299),
            .I(N__42293));
    Odrv12 I__6219 (
            .O(N__42296),
            .I(throttle_order_4));
    Odrv4 I__6218 (
            .O(N__42293),
            .I(throttle_order_4));
    CascadeMux I__6217 (
            .O(N__42288),
            .I(N__42283));
    InMux I__6216 (
            .O(N__42287),
            .I(N__42276));
    InMux I__6215 (
            .O(N__42286),
            .I(N__42276));
    InMux I__6214 (
            .O(N__42283),
            .I(N__42276));
    LocalMux I__6213 (
            .O(N__42276),
            .I(\ppm_encoder_1.throttleZ0Z_4 ));
    InMux I__6212 (
            .O(N__42273),
            .I(\ppm_encoder_1.un1_rudder_cry_6 ));
    CascadeMux I__6211 (
            .O(N__42270),
            .I(\ppm_encoder_1.un2_throttle_iv_0_2_8_cascade_ ));
    CascadeMux I__6210 (
            .O(N__42267),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_8_cascade_ ));
    InMux I__6209 (
            .O(N__42264),
            .I(N__42261));
    LocalMux I__6208 (
            .O(N__42261),
            .I(\ppm_encoder_1.un2_throttle_iv_0_1_8 ));
    CascadeMux I__6207 (
            .O(N__42258),
            .I(\ppm_encoder_1.un2_throttle_iv_0_2_3_cascade_ ));
    CascadeMux I__6206 (
            .O(N__42255),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_3_cascade_ ));
    CascadeMux I__6205 (
            .O(N__42252),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_4_cascade_ ));
    CascadeMux I__6204 (
            .O(N__42249),
            .I(\ppm_encoder_1.elevator_RNIC96OZ0Z_5_cascade_ ));
    InMux I__6203 (
            .O(N__42246),
            .I(N__42243));
    LocalMux I__6202 (
            .O(N__42243),
            .I(\ppm_encoder_1.un2_throttle_iv_0_0_5 ));
    CascadeMux I__6201 (
            .O(N__42240),
            .I(\ppm_encoder_1.un2_throttle_iv_0_1_5_cascade_ ));
    CascadeMux I__6200 (
            .O(N__42237),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_5_cascade_ ));
    InMux I__6199 (
            .O(N__42234),
            .I(N__42228));
    InMux I__6198 (
            .O(N__42233),
            .I(N__42228));
    LocalMux I__6197 (
            .O(N__42228),
            .I(\ppm_encoder_1.elevatorZ0Z_5 ));
    CascadeMux I__6196 (
            .O(N__42225),
            .I(\ppm_encoder_1.elevator_RNIFC6OZ0Z_8_cascade_ ));
    CascadeMux I__6195 (
            .O(N__42222),
            .I(\pid_front.un1_pid_prereg_0_25_cascade_ ));
    InMux I__6194 (
            .O(N__42219),
            .I(N__42210));
    InMux I__6193 (
            .O(N__42218),
            .I(N__42210));
    InMux I__6192 (
            .O(N__42217),
            .I(N__42210));
    LocalMux I__6191 (
            .O(N__42210),
            .I(\pid_front.un1_pid_prereg_0_24 ));
    CascadeMux I__6190 (
            .O(N__42207),
            .I(N__42203));
    CascadeMux I__6189 (
            .O(N__42206),
            .I(N__42199));
    InMux I__6188 (
            .O(N__42203),
            .I(N__42192));
    InMux I__6187 (
            .O(N__42202),
            .I(N__42192));
    InMux I__6186 (
            .O(N__42199),
            .I(N__42192));
    LocalMux I__6185 (
            .O(N__42192),
            .I(\pid_front.un1_pid_prereg_0_26 ));
    InMux I__6184 (
            .O(N__42189),
            .I(N__42174));
    InMux I__6183 (
            .O(N__42188),
            .I(N__42174));
    InMux I__6182 (
            .O(N__42187),
            .I(N__42174));
    InMux I__6181 (
            .O(N__42186),
            .I(N__42174));
    InMux I__6180 (
            .O(N__42185),
            .I(N__42174));
    LocalMux I__6179 (
            .O(N__42174),
            .I(\pid_front.un1_pid_prereg_0_25 ));
    CascadeMux I__6178 (
            .O(N__42171),
            .I(N__42168));
    InMux I__6177 (
            .O(N__42168),
            .I(N__42163));
    InMux I__6176 (
            .O(N__42167),
            .I(N__42158));
    InMux I__6175 (
            .O(N__42166),
            .I(N__42158));
    LocalMux I__6174 (
            .O(N__42163),
            .I(\pid_front.un1_pid_prereg_0_23 ));
    LocalMux I__6173 (
            .O(N__42158),
            .I(\pid_front.un1_pid_prereg_0_23 ));
    CascadeMux I__6172 (
            .O(N__42153),
            .I(N__42150));
    InMux I__6171 (
            .O(N__42150),
            .I(N__42147));
    LocalMux I__6170 (
            .O(N__42147),
            .I(N__42142));
    InMux I__6169 (
            .O(N__42146),
            .I(N__42137));
    InMux I__6168 (
            .O(N__42145),
            .I(N__42137));
    Span4Mux_s1_v I__6167 (
            .O(N__42142),
            .I(N__42134));
    LocalMux I__6166 (
            .O(N__42137),
            .I(\ppm_encoder_1.throttleZ0Z_5 ));
    Odrv4 I__6165 (
            .O(N__42134),
            .I(\ppm_encoder_1.throttleZ0Z_5 ));
    CascadeMux I__6164 (
            .O(N__42129),
            .I(\pid_front.un1_pid_prereg_0_22_cascade_ ));
    InMux I__6163 (
            .O(N__42126),
            .I(N__42122));
    InMux I__6162 (
            .O(N__42125),
            .I(N__42119));
    LocalMux I__6161 (
            .O(N__42122),
            .I(\pid_front.un1_pid_prereg_0_20 ));
    LocalMux I__6160 (
            .O(N__42119),
            .I(\pid_front.un1_pid_prereg_0_20 ));
    InMux I__6159 (
            .O(N__42114),
            .I(N__42105));
    InMux I__6158 (
            .O(N__42113),
            .I(N__42105));
    InMux I__6157 (
            .O(N__42112),
            .I(N__42105));
    LocalMux I__6156 (
            .O(N__42105),
            .I(\pid_front.un1_pid_prereg_0_21 ));
    CascadeMux I__6155 (
            .O(N__42102),
            .I(\pid_front.un1_pid_prereg_0_20_cascade_ ));
    InMux I__6154 (
            .O(N__42099),
            .I(N__42096));
    LocalMux I__6153 (
            .O(N__42096),
            .I(N__42092));
    InMux I__6152 (
            .O(N__42095),
            .I(N__42089));
    Odrv4 I__6151 (
            .O(N__42092),
            .I(\pid_front.un1_pid_prereg_0_22 ));
    LocalMux I__6150 (
            .O(N__42089),
            .I(\pid_front.un1_pid_prereg_0_22 ));
    InMux I__6149 (
            .O(N__42084),
            .I(N__42081));
    LocalMux I__6148 (
            .O(N__42081),
            .I(\pid_front.source_pid_1_sqmuxa_1_0_a4_3 ));
    CascadeMux I__6147 (
            .O(N__42078),
            .I(\pid_front.N_98_cascade_ ));
    CascadeMux I__6146 (
            .O(N__42075),
            .I(\pid_front.un1_pid_prereg_0_9_cascade_ ));
    CascadeMux I__6145 (
            .O(N__42072),
            .I(\pid_front.un1_pid_prereg_0_10_cascade_ ));
    InMux I__6144 (
            .O(N__42069),
            .I(N__42063));
    InMux I__6143 (
            .O(N__42068),
            .I(N__42063));
    LocalMux I__6142 (
            .O(N__42063),
            .I(\pid_front.un1_pid_prereg_0_8 ));
    CascadeMux I__6141 (
            .O(N__42060),
            .I(\pid_front.un1_pid_prereg_0_8_cascade_ ));
    InMux I__6140 (
            .O(N__42057),
            .I(N__42053));
    InMux I__6139 (
            .O(N__42056),
            .I(N__42050));
    LocalMux I__6138 (
            .O(N__42053),
            .I(\pid_front.un1_pid_prereg_0_9 ));
    LocalMux I__6137 (
            .O(N__42050),
            .I(\pid_front.un1_pid_prereg_0_9 ));
    InMux I__6136 (
            .O(N__42045),
            .I(N__42042));
    LocalMux I__6135 (
            .O(N__42042),
            .I(N__42039));
    Odrv4 I__6134 (
            .O(N__42039),
            .I(\pid_front.N_11_i ));
    InMux I__6133 (
            .O(N__42036),
            .I(N__42033));
    LocalMux I__6132 (
            .O(N__42033),
            .I(N__42030));
    Odrv4 I__6131 (
            .O(N__42030),
            .I(\pid_front.un11lto30_i_a2_0_and ));
    InMux I__6130 (
            .O(N__42027),
            .I(N__42024));
    LocalMux I__6129 (
            .O(N__42024),
            .I(N__42021));
    Odrv4 I__6128 (
            .O(N__42021),
            .I(\pid_front.un11lto30_i_a2_2_and ));
    InMux I__6127 (
            .O(N__42018),
            .I(N__42013));
    InMux I__6126 (
            .O(N__42017),
            .I(N__42008));
    InMux I__6125 (
            .O(N__42016),
            .I(N__42008));
    LocalMux I__6124 (
            .O(N__42013),
            .I(\pid_front.pid_preregZ0Z_14 ));
    LocalMux I__6123 (
            .O(N__42008),
            .I(\pid_front.pid_preregZ0Z_14 ));
    InMux I__6122 (
            .O(N__42003),
            .I(N__42000));
    LocalMux I__6121 (
            .O(N__42000),
            .I(N__41997));
    Odrv4 I__6120 (
            .O(N__41997),
            .I(\pid_front.un11lto30_i_a2_4_and ));
    InMux I__6119 (
            .O(N__41994),
            .I(N__41990));
    InMux I__6118 (
            .O(N__41993),
            .I(N__41987));
    LocalMux I__6117 (
            .O(N__41990),
            .I(N__41984));
    LocalMux I__6116 (
            .O(N__41987),
            .I(N__41979));
    Span4Mux_v I__6115 (
            .O(N__41984),
            .I(N__41979));
    Odrv4 I__6114 (
            .O(N__41979),
            .I(\pid_front.un11lto30_i_a2_5_and ));
    CascadeMux I__6113 (
            .O(N__41976),
            .I(\pid_front.un11lto30_i_a2_4_and_cascade_ ));
    InMux I__6112 (
            .O(N__41973),
            .I(N__41970));
    LocalMux I__6111 (
            .O(N__41970),
            .I(N__41967));
    Odrv4 I__6110 (
            .O(N__41967),
            .I(\pid_front.source_pid_1_sqmuxa_1_0_a2_0_0 ));
    InMux I__6109 (
            .O(N__41964),
            .I(bfn_8_16_0_));
    CascadeMux I__6108 (
            .O(N__41961),
            .I(N__41957));
    InMux I__6107 (
            .O(N__41960),
            .I(N__41952));
    InMux I__6106 (
            .O(N__41957),
            .I(N__41944));
    InMux I__6105 (
            .O(N__41956),
            .I(N__41944));
    InMux I__6104 (
            .O(N__41955),
            .I(N__41944));
    LocalMux I__6103 (
            .O(N__41952),
            .I(N__41941));
    InMux I__6102 (
            .O(N__41951),
            .I(N__41938));
    LocalMux I__6101 (
            .O(N__41944),
            .I(N__41935));
    Span4Mux_v I__6100 (
            .O(N__41941),
            .I(N__41930));
    LocalMux I__6099 (
            .O(N__41938),
            .I(N__41930));
    Span4Mux_v I__6098 (
            .O(N__41935),
            .I(N__41927));
    Span4Mux_h I__6097 (
            .O(N__41930),
            .I(N__41924));
    Odrv4 I__6096 (
            .O(N__41927),
            .I(\uart_pc.N_143 ));
    Odrv4 I__6095 (
            .O(N__41924),
            .I(\uart_pc.N_143 ));
    InMux I__6094 (
            .O(N__41919),
            .I(N__41916));
    LocalMux I__6093 (
            .O(N__41916),
            .I(N__41910));
    CascadeMux I__6092 (
            .O(N__41915),
            .I(N__41907));
    CascadeMux I__6091 (
            .O(N__41914),
            .I(N__41903));
    CascadeMux I__6090 (
            .O(N__41913),
            .I(N__41900));
    Span4Mux_v I__6089 (
            .O(N__41910),
            .I(N__41897));
    InMux I__6088 (
            .O(N__41907),
            .I(N__41894));
    InMux I__6087 (
            .O(N__41906),
            .I(N__41887));
    InMux I__6086 (
            .O(N__41903),
            .I(N__41887));
    InMux I__6085 (
            .O(N__41900),
            .I(N__41887));
    Span4Mux_h I__6084 (
            .O(N__41897),
            .I(N__41880));
    LocalMux I__6083 (
            .O(N__41894),
            .I(N__41880));
    LocalMux I__6082 (
            .O(N__41887),
            .I(N__41880));
    Odrv4 I__6081 (
            .O(N__41880),
            .I(\uart_pc.timer_Count_0_sqmuxa ));
    InMux I__6080 (
            .O(N__41877),
            .I(N__41874));
    LocalMux I__6079 (
            .O(N__41874),
            .I(N__41869));
    CascadeMux I__6078 (
            .O(N__41873),
            .I(N__41865));
    InMux I__6077 (
            .O(N__41872),
            .I(N__41862));
    Span4Mux_h I__6076 (
            .O(N__41869),
            .I(N__41859));
    InMux I__6075 (
            .O(N__41868),
            .I(N__41854));
    InMux I__6074 (
            .O(N__41865),
            .I(N__41854));
    LocalMux I__6073 (
            .O(N__41862),
            .I(\uart_pc.timer_CountZ0Z_0 ));
    Odrv4 I__6072 (
            .O(N__41859),
            .I(\uart_pc.timer_CountZ0Z_0 ));
    LocalMux I__6071 (
            .O(N__41854),
            .I(\uart_pc.timer_CountZ0Z_0 ));
    InMux I__6070 (
            .O(N__41847),
            .I(N__41843));
    InMux I__6069 (
            .O(N__41846),
            .I(N__41840));
    LocalMux I__6068 (
            .O(N__41843),
            .I(\pid_front.un11lto30_i_a2_3_and ));
    LocalMux I__6067 (
            .O(N__41840),
            .I(\pid_front.un11lto30_i_a2_3_and ));
    CascadeMux I__6066 (
            .O(N__41835),
            .I(N__41832));
    InMux I__6065 (
            .O(N__41832),
            .I(N__41829));
    LocalMux I__6064 (
            .O(N__41829),
            .I(\pid_front.source_pid_1_sqmuxa_1_0_a2_1_4 ));
    InMux I__6063 (
            .O(N__41826),
            .I(\dron_frame_decoder_1.un1_WDT_cry_10 ));
    InMux I__6062 (
            .O(N__41823),
            .I(\dron_frame_decoder_1.un1_WDT_cry_11 ));
    InMux I__6061 (
            .O(N__41820),
            .I(\dron_frame_decoder_1.un1_WDT_cry_12 ));
    InMux I__6060 (
            .O(N__41817),
            .I(\dron_frame_decoder_1.un1_WDT_cry_13 ));
    InMux I__6059 (
            .O(N__41814),
            .I(\dron_frame_decoder_1.un1_WDT_cry_14 ));
    SRMux I__6058 (
            .O(N__41811),
            .I(N__41807));
    SRMux I__6057 (
            .O(N__41810),
            .I(N__41804));
    LocalMux I__6056 (
            .O(N__41807),
            .I(N__41801));
    LocalMux I__6055 (
            .O(N__41804),
            .I(N__41798));
    Span4Mux_v I__6054 (
            .O(N__41801),
            .I(N__41795));
    Span4Mux_v I__6053 (
            .O(N__41798),
            .I(N__41790));
    Span4Mux_h I__6052 (
            .O(N__41795),
            .I(N__41790));
    Odrv4 I__6051 (
            .O(N__41790),
            .I(\dron_frame_decoder_1.source_data_valid_2_sqmuxa_iZ0 ));
    InMux I__6050 (
            .O(N__41787),
            .I(N__41784));
    LocalMux I__6049 (
            .O(N__41784),
            .I(\dron_frame_decoder_1.WDTZ0Z_2 ));
    InMux I__6048 (
            .O(N__41781),
            .I(\dron_frame_decoder_1.un1_WDT_cry_1 ));
    InMux I__6047 (
            .O(N__41778),
            .I(N__41775));
    LocalMux I__6046 (
            .O(N__41775),
            .I(\dron_frame_decoder_1.WDTZ0Z_3 ));
    InMux I__6045 (
            .O(N__41772),
            .I(\dron_frame_decoder_1.un1_WDT_cry_2 ));
    InMux I__6044 (
            .O(N__41769),
            .I(\dron_frame_decoder_1.un1_WDT_cry_3 ));
    InMux I__6043 (
            .O(N__41766),
            .I(\dron_frame_decoder_1.un1_WDT_cry_4 ));
    InMux I__6042 (
            .O(N__41763),
            .I(\dron_frame_decoder_1.un1_WDT_cry_5 ));
    InMux I__6041 (
            .O(N__41760),
            .I(\dron_frame_decoder_1.un1_WDT_cry_6 ));
    InMux I__6040 (
            .O(N__41757),
            .I(bfn_8_14_0_));
    InMux I__6039 (
            .O(N__41754),
            .I(\dron_frame_decoder_1.un1_WDT_cry_8 ));
    InMux I__6038 (
            .O(N__41751),
            .I(\dron_frame_decoder_1.un1_WDT_cry_9 ));
    CEMux I__6037 (
            .O(N__41748),
            .I(N__41745));
    LocalMux I__6036 (
            .O(N__41745),
            .I(N__41742));
    Span4Mux_v I__6035 (
            .O(N__41742),
            .I(N__41739));
    Span4Mux_h I__6034 (
            .O(N__41739),
            .I(N__41736));
    Odrv4 I__6033 (
            .O(N__41736),
            .I(\Commands_frame_decoder.source_offset4data_1_sqmuxa_0 ));
    InMux I__6032 (
            .O(N__41733),
            .I(N__41730));
    LocalMux I__6031 (
            .O(N__41730),
            .I(\dron_frame_decoder_1.WDTZ0Z_0 ));
    InMux I__6030 (
            .O(N__41727),
            .I(N__41724));
    LocalMux I__6029 (
            .O(N__41724),
            .I(\dron_frame_decoder_1.WDTZ0Z_1 ));
    InMux I__6028 (
            .O(N__41721),
            .I(\dron_frame_decoder_1.un1_WDT_cry_0 ));
    CascadeMux I__6027 (
            .O(N__41718),
            .I(\uart_drone.timer_Count_RNIES9Q1Z0Z_2_cascade_ ));
    InMux I__6026 (
            .O(N__41715),
            .I(N__41711));
    InMux I__6025 (
            .O(N__41714),
            .I(N__41708));
    LocalMux I__6024 (
            .O(N__41711),
            .I(N__41704));
    LocalMux I__6023 (
            .O(N__41708),
            .I(N__41701));
    InMux I__6022 (
            .O(N__41707),
            .I(N__41697));
    Span4Mux_v I__6021 (
            .O(N__41704),
            .I(N__41694));
    Span4Mux_h I__6020 (
            .O(N__41701),
            .I(N__41691));
    InMux I__6019 (
            .O(N__41700),
            .I(N__41688));
    LocalMux I__6018 (
            .O(N__41697),
            .I(\uart_pc.N_152 ));
    Odrv4 I__6017 (
            .O(N__41694),
            .I(\uart_pc.N_152 ));
    Odrv4 I__6016 (
            .O(N__41691),
            .I(\uart_pc.N_152 ));
    LocalMux I__6015 (
            .O(N__41688),
            .I(\uart_pc.N_152 ));
    CascadeMux I__6014 (
            .O(N__41679),
            .I(N__41674));
    InMux I__6013 (
            .O(N__41678),
            .I(N__41671));
    InMux I__6012 (
            .O(N__41677),
            .I(N__41668));
    InMux I__6011 (
            .O(N__41674),
            .I(N__41665));
    LocalMux I__6010 (
            .O(N__41671),
            .I(N__41662));
    LocalMux I__6009 (
            .O(N__41668),
            .I(N__41659));
    LocalMux I__6008 (
            .O(N__41665),
            .I(\uart_pc.un1_state_4_0 ));
    Odrv4 I__6007 (
            .O(N__41662),
            .I(\uart_pc.un1_state_4_0 ));
    Odrv4 I__6006 (
            .O(N__41659),
            .I(\uart_pc.un1_state_4_0 ));
    CascadeMux I__6005 (
            .O(N__41652),
            .I(N__41646));
    InMux I__6004 (
            .O(N__41651),
            .I(N__41642));
    InMux I__6003 (
            .O(N__41650),
            .I(N__41639));
    InMux I__6002 (
            .O(N__41649),
            .I(N__41636));
    InMux I__6001 (
            .O(N__41646),
            .I(N__41633));
    CascadeMux I__6000 (
            .O(N__41645),
            .I(N__41630));
    LocalMux I__5999 (
            .O(N__41642),
            .I(N__41624));
    LocalMux I__5998 (
            .O(N__41639),
            .I(N__41619));
    LocalMux I__5997 (
            .O(N__41636),
            .I(N__41619));
    LocalMux I__5996 (
            .O(N__41633),
            .I(N__41616));
    InMux I__5995 (
            .O(N__41630),
            .I(N__41611));
    InMux I__5994 (
            .O(N__41629),
            .I(N__41611));
    InMux I__5993 (
            .O(N__41628),
            .I(N__41606));
    InMux I__5992 (
            .O(N__41627),
            .I(N__41606));
    Span4Mux_v I__5991 (
            .O(N__41624),
            .I(N__41601));
    Span4Mux_v I__5990 (
            .O(N__41619),
            .I(N__41601));
    Span4Mux_v I__5989 (
            .O(N__41616),
            .I(N__41596));
    LocalMux I__5988 (
            .O(N__41611),
            .I(N__41596));
    LocalMux I__5987 (
            .O(N__41606),
            .I(\uart_pc.stateZ0Z_3 ));
    Odrv4 I__5986 (
            .O(N__41601),
            .I(\uart_pc.stateZ0Z_3 ));
    Odrv4 I__5985 (
            .O(N__41596),
            .I(\uart_pc.stateZ0Z_3 ));
    InMux I__5984 (
            .O(N__41589),
            .I(N__41568));
    InMux I__5983 (
            .O(N__41588),
            .I(N__41568));
    InMux I__5982 (
            .O(N__41587),
            .I(N__41568));
    InMux I__5981 (
            .O(N__41586),
            .I(N__41568));
    InMux I__5980 (
            .O(N__41585),
            .I(N__41568));
    InMux I__5979 (
            .O(N__41584),
            .I(N__41568));
    InMux I__5978 (
            .O(N__41583),
            .I(N__41568));
    LocalMux I__5977 (
            .O(N__41568),
            .I(N__41562));
    InMux I__5976 (
            .O(N__41567),
            .I(N__41559));
    InMux I__5975 (
            .O(N__41566),
            .I(N__41556));
    InMux I__5974 (
            .O(N__41565),
            .I(N__41552));
    Span4Mux_h I__5973 (
            .O(N__41562),
            .I(N__41549));
    LocalMux I__5972 (
            .O(N__41559),
            .I(N__41544));
    LocalMux I__5971 (
            .O(N__41556),
            .I(N__41544));
    InMux I__5970 (
            .O(N__41555),
            .I(N__41541));
    LocalMux I__5969 (
            .O(N__41552),
            .I(\uart_pc.bit_CountZ0Z_0 ));
    Odrv4 I__5968 (
            .O(N__41549),
            .I(\uart_pc.bit_CountZ0Z_0 ));
    Odrv4 I__5967 (
            .O(N__41544),
            .I(\uart_pc.bit_CountZ0Z_0 ));
    LocalMux I__5966 (
            .O(N__41541),
            .I(\uart_pc.bit_CountZ0Z_0 ));
    CEMux I__5965 (
            .O(N__41532),
            .I(N__41528));
    CEMux I__5964 (
            .O(N__41531),
            .I(N__41525));
    LocalMux I__5963 (
            .O(N__41528),
            .I(N__41522));
    LocalMux I__5962 (
            .O(N__41525),
            .I(N__41519));
    Span4Mux_h I__5961 (
            .O(N__41522),
            .I(N__41516));
    Span4Mux_h I__5960 (
            .O(N__41519),
            .I(N__41513));
    Span4Mux_h I__5959 (
            .O(N__41516),
            .I(N__41510));
    Span4Mux_v I__5958 (
            .O(N__41513),
            .I(N__41507));
    Odrv4 I__5957 (
            .O(N__41510),
            .I(\Commands_frame_decoder.source_CH4data_1_sqmuxa_0 ));
    Odrv4 I__5956 (
            .O(N__41507),
            .I(\Commands_frame_decoder.source_CH4data_1_sqmuxa_0 ));
    InMux I__5955 (
            .O(N__41502),
            .I(N__41497));
    InMux I__5954 (
            .O(N__41501),
            .I(N__41494));
    CascadeMux I__5953 (
            .O(N__41500),
            .I(N__41491));
    LocalMux I__5952 (
            .O(N__41497),
            .I(N__41488));
    LocalMux I__5951 (
            .O(N__41494),
            .I(N__41485));
    InMux I__5950 (
            .O(N__41491),
            .I(N__41482));
    Span4Mux_h I__5949 (
            .O(N__41488),
            .I(N__41479));
    Span4Mux_h I__5948 (
            .O(N__41485),
            .I(N__41476));
    LocalMux I__5947 (
            .O(N__41482),
            .I(throttle_order_11));
    Odrv4 I__5946 (
            .O(N__41479),
            .I(throttle_order_11));
    Odrv4 I__5945 (
            .O(N__41476),
            .I(throttle_order_11));
    InMux I__5944 (
            .O(N__41469),
            .I(N__41466));
    LocalMux I__5943 (
            .O(N__41466),
            .I(N__41463));
    Odrv4 I__5942 (
            .O(N__41463),
            .I(\ppm_encoder_1.un1_throttle_cry_10_THRU_CO ));
    InMux I__5941 (
            .O(N__41460),
            .I(\ppm_encoder_1.un1_throttle_cry_10 ));
    InMux I__5940 (
            .O(N__41457),
            .I(\ppm_encoder_1.un1_throttle_cry_11 ));
    InMux I__5939 (
            .O(N__41454),
            .I(\ppm_encoder_1.un1_throttle_cry_12 ));
    InMux I__5938 (
            .O(N__41451),
            .I(\ppm_encoder_1.un1_throttle_cry_13 ));
    InMux I__5937 (
            .O(N__41448),
            .I(N__41445));
    LocalMux I__5936 (
            .O(N__41445),
            .I(N__41442));
    Odrv4 I__5935 (
            .O(N__41442),
            .I(\ppm_encoder_1.un1_throttle_cry_5_THRU_CO ));
    CascadeMux I__5934 (
            .O(N__41439),
            .I(N__41436));
    InMux I__5933 (
            .O(N__41436),
            .I(N__41432));
    InMux I__5932 (
            .O(N__41435),
            .I(N__41428));
    LocalMux I__5931 (
            .O(N__41432),
            .I(N__41425));
    InMux I__5930 (
            .O(N__41431),
            .I(N__41422));
    LocalMux I__5929 (
            .O(N__41428),
            .I(N__41419));
    Span4Mux_h I__5928 (
            .O(N__41425),
            .I(N__41416));
    LocalMux I__5927 (
            .O(N__41422),
            .I(throttle_order_6));
    Odrv4 I__5926 (
            .O(N__41419),
            .I(throttle_order_6));
    Odrv4 I__5925 (
            .O(N__41416),
            .I(throttle_order_6));
    InMux I__5924 (
            .O(N__41409),
            .I(N__41404));
    CascadeMux I__5923 (
            .O(N__41408),
            .I(N__41401));
    InMux I__5922 (
            .O(N__41407),
            .I(N__41398));
    LocalMux I__5921 (
            .O(N__41404),
            .I(N__41395));
    InMux I__5920 (
            .O(N__41401),
            .I(N__41392));
    LocalMux I__5919 (
            .O(N__41398),
            .I(N__41389));
    Span4Mux_h I__5918 (
            .O(N__41395),
            .I(N__41386));
    LocalMux I__5917 (
            .O(N__41392),
            .I(throttle_order_8));
    Odrv12 I__5916 (
            .O(N__41389),
            .I(throttle_order_8));
    Odrv4 I__5915 (
            .O(N__41386),
            .I(throttle_order_8));
    InMux I__5914 (
            .O(N__41379),
            .I(N__41376));
    LocalMux I__5913 (
            .O(N__41376),
            .I(\ppm_encoder_1.un1_throttle_cry_7_THRU_CO ));
    IoInMux I__5912 (
            .O(N__41373),
            .I(N__41370));
    LocalMux I__5911 (
            .O(N__41370),
            .I(N__41367));
    IoSpan4Mux I__5910 (
            .O(N__41367),
            .I(N__41364));
    Span4Mux_s3_v I__5909 (
            .O(N__41364),
            .I(N__41359));
    InMux I__5908 (
            .O(N__41363),
            .I(N__41354));
    InMux I__5907 (
            .O(N__41362),
            .I(N__41354));
    Sp12to4 I__5906 (
            .O(N__41359),
            .I(N__41351));
    LocalMux I__5905 (
            .O(N__41354),
            .I(N__41348));
    Span12Mux_s8_v I__5904 (
            .O(N__41351),
            .I(N__41345));
    Span4Mux_h I__5903 (
            .O(N__41348),
            .I(N__41341));
    Span12Mux_h I__5902 (
            .O(N__41345),
            .I(N__41338));
    InMux I__5901 (
            .O(N__41344),
            .I(N__41335));
    Span4Mux_h I__5900 (
            .O(N__41341),
            .I(N__41332));
    Odrv12 I__5899 (
            .O(N__41338),
            .I(debug_CH3_20A_c));
    LocalMux I__5898 (
            .O(N__41335),
            .I(debug_CH3_20A_c));
    Odrv4 I__5897 (
            .O(N__41332),
            .I(debug_CH3_20A_c));
    InMux I__5896 (
            .O(N__41325),
            .I(N__41322));
    LocalMux I__5895 (
            .O(N__41322),
            .I(N__41318));
    InMux I__5894 (
            .O(N__41321),
            .I(N__41315));
    Span4Mux_v I__5893 (
            .O(N__41318),
            .I(N__41310));
    LocalMux I__5892 (
            .O(N__41315),
            .I(N__41310));
    Span4Mux_h I__5891 (
            .O(N__41310),
            .I(N__41307));
    Odrv4 I__5890 (
            .O(N__41307),
            .I(throttle_order_3));
    InMux I__5889 (
            .O(N__41304),
            .I(N__41301));
    LocalMux I__5888 (
            .O(N__41301),
            .I(\ppm_encoder_1.un1_throttle_cry_2_THRU_CO ));
    InMux I__5887 (
            .O(N__41298),
            .I(\ppm_encoder_1.un1_throttle_cry_2 ));
    InMux I__5886 (
            .O(N__41295),
            .I(\ppm_encoder_1.un1_throttle_cry_3 ));
    InMux I__5885 (
            .O(N__41292),
            .I(N__41288));
    InMux I__5884 (
            .O(N__41291),
            .I(N__41285));
    LocalMux I__5883 (
            .O(N__41288),
            .I(N__41282));
    LocalMux I__5882 (
            .O(N__41285),
            .I(N__41279));
    Span4Mux_h I__5881 (
            .O(N__41282),
            .I(N__41276));
    Span4Mux_h I__5880 (
            .O(N__41279),
            .I(N__41273));
    Span4Mux_v I__5879 (
            .O(N__41276),
            .I(N__41270));
    Span4Mux_v I__5878 (
            .O(N__41273),
            .I(N__41267));
    Span4Mux_v I__5877 (
            .O(N__41270),
            .I(N__41264));
    Span4Mux_h I__5876 (
            .O(N__41267),
            .I(N__41261));
    Odrv4 I__5875 (
            .O(N__41264),
            .I(throttle_order_5));
    Odrv4 I__5874 (
            .O(N__41261),
            .I(throttle_order_5));
    InMux I__5873 (
            .O(N__41256),
            .I(N__41253));
    LocalMux I__5872 (
            .O(N__41253),
            .I(N__41250));
    Odrv4 I__5871 (
            .O(N__41250),
            .I(\ppm_encoder_1.un1_throttle_cry_4_THRU_CO ));
    InMux I__5870 (
            .O(N__41247),
            .I(\ppm_encoder_1.un1_throttle_cry_4 ));
    InMux I__5869 (
            .O(N__41244),
            .I(\ppm_encoder_1.un1_throttle_cry_5 ));
    InMux I__5868 (
            .O(N__41241),
            .I(\ppm_encoder_1.un1_throttle_cry_6 ));
    InMux I__5867 (
            .O(N__41238),
            .I(bfn_8_9_0_));
    InMux I__5866 (
            .O(N__41235),
            .I(N__41232));
    LocalMux I__5865 (
            .O(N__41232),
            .I(N__41228));
    InMux I__5864 (
            .O(N__41231),
            .I(N__41225));
    Span4Mux_v I__5863 (
            .O(N__41228),
            .I(N__41219));
    LocalMux I__5862 (
            .O(N__41225),
            .I(N__41219));
    InMux I__5861 (
            .O(N__41224),
            .I(N__41216));
    Span4Mux_h I__5860 (
            .O(N__41219),
            .I(N__41213));
    LocalMux I__5859 (
            .O(N__41216),
            .I(throttle_order_9));
    Odrv4 I__5858 (
            .O(N__41213),
            .I(throttle_order_9));
    InMux I__5857 (
            .O(N__41208),
            .I(N__41205));
    LocalMux I__5856 (
            .O(N__41205),
            .I(N__41202));
    Odrv4 I__5855 (
            .O(N__41202),
            .I(\ppm_encoder_1.un1_throttle_cry_8_THRU_CO ));
    InMux I__5854 (
            .O(N__41199),
            .I(\ppm_encoder_1.un1_throttle_cry_8 ));
    InMux I__5853 (
            .O(N__41196),
            .I(\ppm_encoder_1.un1_throttle_cry_9 ));
    InMux I__5852 (
            .O(N__41193),
            .I(\ppm_encoder_1.un1_throttle_cry_0 ));
    InMux I__5851 (
            .O(N__41190),
            .I(\ppm_encoder_1.un1_throttle_cry_1 ));
    InMux I__5850 (
            .O(N__41187),
            .I(\reset_module_System.count_1_cry_18 ));
    InMux I__5849 (
            .O(N__41184),
            .I(N__41180));
    InMux I__5848 (
            .O(N__41183),
            .I(N__41177));
    LocalMux I__5847 (
            .O(N__41180),
            .I(N__41174));
    LocalMux I__5846 (
            .O(N__41177),
            .I(\reset_module_System.countZ0Z_20 ));
    Odrv4 I__5845 (
            .O(N__41174),
            .I(\reset_module_System.countZ0Z_20 ));
    InMux I__5844 (
            .O(N__41169),
            .I(\reset_module_System.count_1_cry_19 ));
    InMux I__5843 (
            .O(N__41166),
            .I(\reset_module_System.count_1_cry_20 ));
    InMux I__5842 (
            .O(N__41163),
            .I(N__41159));
    InMux I__5841 (
            .O(N__41162),
            .I(N__41156));
    LocalMux I__5840 (
            .O(N__41159),
            .I(\reset_module_System.countZ0Z_10 ));
    LocalMux I__5839 (
            .O(N__41156),
            .I(\reset_module_System.countZ0Z_10 ));
    InMux I__5838 (
            .O(N__41151),
            .I(N__41147));
    InMux I__5837 (
            .O(N__41150),
            .I(N__41144));
    LocalMux I__5836 (
            .O(N__41147),
            .I(\reset_module_System.countZ0Z_11 ));
    LocalMux I__5835 (
            .O(N__41144),
            .I(\reset_module_System.countZ0Z_11 ));
    InMux I__5834 (
            .O(N__41139),
            .I(N__41136));
    LocalMux I__5833 (
            .O(N__41136),
            .I(\reset_module_System.reset6_3 ));
    InMux I__5832 (
            .O(N__41133),
            .I(N__41129));
    InMux I__5831 (
            .O(N__41132),
            .I(N__41126));
    LocalMux I__5830 (
            .O(N__41129),
            .I(\reset_module_System.countZ0Z_19 ));
    LocalMux I__5829 (
            .O(N__41126),
            .I(\reset_module_System.countZ0Z_19 ));
    InMux I__5828 (
            .O(N__41121),
            .I(N__41118));
    LocalMux I__5827 (
            .O(N__41118),
            .I(N__41114));
    InMux I__5826 (
            .O(N__41117),
            .I(N__41111));
    Odrv4 I__5825 (
            .O(N__41114),
            .I(\reset_module_System.countZ0Z_15 ));
    LocalMux I__5824 (
            .O(N__41111),
            .I(\reset_module_System.countZ0Z_15 ));
    CascadeMux I__5823 (
            .O(N__41106),
            .I(N__41102));
    InMux I__5822 (
            .O(N__41105),
            .I(N__41099));
    InMux I__5821 (
            .O(N__41102),
            .I(N__41096));
    LocalMux I__5820 (
            .O(N__41099),
            .I(\reset_module_System.countZ0Z_21 ));
    LocalMux I__5819 (
            .O(N__41096),
            .I(\reset_module_System.countZ0Z_21 ));
    InMux I__5818 (
            .O(N__41091),
            .I(N__41088));
    LocalMux I__5817 (
            .O(N__41088),
            .I(N__41084));
    InMux I__5816 (
            .O(N__41087),
            .I(N__41081));
    Odrv4 I__5815 (
            .O(N__41084),
            .I(\reset_module_System.countZ0Z_13 ));
    LocalMux I__5814 (
            .O(N__41081),
            .I(\reset_module_System.countZ0Z_13 ));
    InMux I__5813 (
            .O(N__41076),
            .I(N__41073));
    LocalMux I__5812 (
            .O(N__41073),
            .I(N__41070));
    Odrv4 I__5811 (
            .O(N__41070),
            .I(uart_input_drone_c));
    InMux I__5810 (
            .O(N__41067),
            .I(N__41064));
    LocalMux I__5809 (
            .O(N__41064),
            .I(N__41061));
    Span4Mux_h I__5808 (
            .O(N__41061),
            .I(N__41058));
    Odrv4 I__5807 (
            .O(N__41058),
            .I(\uart_drone_sync.aux_0__0__0_0 ));
    InMux I__5806 (
            .O(N__41055),
            .I(N__41052));
    LocalMux I__5805 (
            .O(N__41052),
            .I(N__41046));
    InMux I__5804 (
            .O(N__41051),
            .I(N__41041));
    InMux I__5803 (
            .O(N__41050),
            .I(N__41041));
    InMux I__5802 (
            .O(N__41049),
            .I(N__41038));
    Odrv4 I__5801 (
            .O(N__41046),
            .I(\reset_module_System.countZ0Z_0 ));
    LocalMux I__5800 (
            .O(N__41041),
            .I(\reset_module_System.countZ0Z_0 ));
    LocalMux I__5799 (
            .O(N__41038),
            .I(\reset_module_System.countZ0Z_0 ));
    CascadeMux I__5798 (
            .O(N__41031),
            .I(N__41027));
    InMux I__5797 (
            .O(N__41030),
            .I(N__41023));
    InMux I__5796 (
            .O(N__41027),
            .I(N__41018));
    InMux I__5795 (
            .O(N__41026),
            .I(N__41018));
    LocalMux I__5794 (
            .O(N__41023),
            .I(N__41012));
    LocalMux I__5793 (
            .O(N__41018),
            .I(N__41012));
    InMux I__5792 (
            .O(N__41017),
            .I(N__41009));
    Span4Mux_s3_v I__5791 (
            .O(N__41012),
            .I(N__41006));
    LocalMux I__5790 (
            .O(N__41009),
            .I(\reset_module_System.reset6_15 ));
    Odrv4 I__5789 (
            .O(N__41006),
            .I(\reset_module_System.reset6_15 ));
    InMux I__5788 (
            .O(N__41001),
            .I(N__40998));
    LocalMux I__5787 (
            .O(N__40998),
            .I(N__40993));
    InMux I__5786 (
            .O(N__40997),
            .I(N__40988));
    InMux I__5785 (
            .O(N__40996),
            .I(N__40988));
    Odrv4 I__5784 (
            .O(N__40993),
            .I(\reset_module_System.reset6_19 ));
    LocalMux I__5783 (
            .O(N__40988),
            .I(\reset_module_System.reset6_19 ));
    CascadeMux I__5782 (
            .O(N__40983),
            .I(\reset_module_System.count_1_1_cascade_ ));
    InMux I__5781 (
            .O(N__40980),
            .I(N__40977));
    LocalMux I__5780 (
            .O(N__40977),
            .I(N__40974));
    Span4Mux_v I__5779 (
            .O(N__40974),
            .I(N__40968));
    InMux I__5778 (
            .O(N__40973),
            .I(N__40965));
    InMux I__5777 (
            .O(N__40972),
            .I(N__40962));
    InMux I__5776 (
            .O(N__40971),
            .I(N__40959));
    Odrv4 I__5775 (
            .O(N__40968),
            .I(\reset_module_System.reset6_14 ));
    LocalMux I__5774 (
            .O(N__40965),
            .I(\reset_module_System.reset6_14 ));
    LocalMux I__5773 (
            .O(N__40962),
            .I(\reset_module_System.reset6_14 ));
    LocalMux I__5772 (
            .O(N__40959),
            .I(\reset_module_System.reset6_14 ));
    CascadeMux I__5771 (
            .O(N__40950),
            .I(N__40946));
    InMux I__5770 (
            .O(N__40949),
            .I(N__40942));
    InMux I__5769 (
            .O(N__40946),
            .I(N__40939));
    InMux I__5768 (
            .O(N__40945),
            .I(N__40936));
    LocalMux I__5767 (
            .O(N__40942),
            .I(N__40933));
    LocalMux I__5766 (
            .O(N__40939),
            .I(N__40930));
    LocalMux I__5765 (
            .O(N__40936),
            .I(\reset_module_System.countZ0Z_1 ));
    Odrv4 I__5764 (
            .O(N__40933),
            .I(\reset_module_System.countZ0Z_1 ));
    Odrv12 I__5763 (
            .O(N__40930),
            .I(\reset_module_System.countZ0Z_1 ));
    InMux I__5762 (
            .O(N__40923),
            .I(\reset_module_System.count_1_cry_9 ));
    InMux I__5761 (
            .O(N__40920),
            .I(\reset_module_System.count_1_cry_10 ));
    InMux I__5760 (
            .O(N__40917),
            .I(N__40914));
    LocalMux I__5759 (
            .O(N__40914),
            .I(N__40910));
    InMux I__5758 (
            .O(N__40913),
            .I(N__40907));
    Odrv12 I__5757 (
            .O(N__40910),
            .I(\reset_module_System.countZ0Z_12 ));
    LocalMux I__5756 (
            .O(N__40907),
            .I(\reset_module_System.countZ0Z_12 ));
    InMux I__5755 (
            .O(N__40902),
            .I(\reset_module_System.count_1_cry_11 ));
    InMux I__5754 (
            .O(N__40899),
            .I(\reset_module_System.count_1_cry_12 ));
    InMux I__5753 (
            .O(N__40896),
            .I(N__40892));
    InMux I__5752 (
            .O(N__40895),
            .I(N__40889));
    LocalMux I__5751 (
            .O(N__40892),
            .I(\reset_module_System.countZ0Z_14 ));
    LocalMux I__5750 (
            .O(N__40889),
            .I(\reset_module_System.countZ0Z_14 ));
    InMux I__5749 (
            .O(N__40884),
            .I(\reset_module_System.count_1_cry_13 ));
    InMux I__5748 (
            .O(N__40881),
            .I(\reset_module_System.count_1_cry_14 ));
    InMux I__5747 (
            .O(N__40878),
            .I(N__40875));
    LocalMux I__5746 (
            .O(N__40875),
            .I(N__40871));
    InMux I__5745 (
            .O(N__40874),
            .I(N__40868));
    Odrv4 I__5744 (
            .O(N__40871),
            .I(\reset_module_System.countZ0Z_16 ));
    LocalMux I__5743 (
            .O(N__40868),
            .I(\reset_module_System.countZ0Z_16 ));
    InMux I__5742 (
            .O(N__40863),
            .I(\reset_module_System.count_1_cry_15 ));
    CascadeMux I__5741 (
            .O(N__40860),
            .I(N__40856));
    InMux I__5740 (
            .O(N__40859),
            .I(N__40853));
    InMux I__5739 (
            .O(N__40856),
            .I(N__40850));
    LocalMux I__5738 (
            .O(N__40853),
            .I(\reset_module_System.countZ0Z_17 ));
    LocalMux I__5737 (
            .O(N__40850),
            .I(\reset_module_System.countZ0Z_17 ));
    InMux I__5736 (
            .O(N__40845),
            .I(bfn_8_3_0_));
    CascadeMux I__5735 (
            .O(N__40842),
            .I(N__40838));
    InMux I__5734 (
            .O(N__40841),
            .I(N__40835));
    InMux I__5733 (
            .O(N__40838),
            .I(N__40832));
    LocalMux I__5732 (
            .O(N__40835),
            .I(\reset_module_System.countZ0Z_18 ));
    LocalMux I__5731 (
            .O(N__40832),
            .I(\reset_module_System.countZ0Z_18 ));
    InMux I__5730 (
            .O(N__40827),
            .I(\reset_module_System.count_1_cry_17 ));
    CascadeMux I__5729 (
            .O(N__40824),
            .I(N__40821));
    InMux I__5728 (
            .O(N__40821),
            .I(N__40817));
    InMux I__5727 (
            .O(N__40820),
            .I(N__40814));
    LocalMux I__5726 (
            .O(N__40817),
            .I(\reset_module_System.countZ0Z_2 ));
    LocalMux I__5725 (
            .O(N__40814),
            .I(\reset_module_System.countZ0Z_2 ));
    InMux I__5724 (
            .O(N__40809),
            .I(N__40806));
    LocalMux I__5723 (
            .O(N__40806),
            .I(\reset_module_System.count_1_2 ));
    InMux I__5722 (
            .O(N__40803),
            .I(\reset_module_System.count_1_cry_1 ));
    InMux I__5721 (
            .O(N__40800),
            .I(N__40796));
    InMux I__5720 (
            .O(N__40799),
            .I(N__40793));
    LocalMux I__5719 (
            .O(N__40796),
            .I(\reset_module_System.countZ0Z_3 ));
    LocalMux I__5718 (
            .O(N__40793),
            .I(\reset_module_System.countZ0Z_3 ));
    InMux I__5717 (
            .O(N__40788),
            .I(\reset_module_System.count_1_cry_2 ));
    InMux I__5716 (
            .O(N__40785),
            .I(N__40781));
    InMux I__5715 (
            .O(N__40784),
            .I(N__40778));
    LocalMux I__5714 (
            .O(N__40781),
            .I(\reset_module_System.countZ0Z_4 ));
    LocalMux I__5713 (
            .O(N__40778),
            .I(\reset_module_System.countZ0Z_4 ));
    InMux I__5712 (
            .O(N__40773),
            .I(\reset_module_System.count_1_cry_3 ));
    InMux I__5711 (
            .O(N__40770),
            .I(N__40766));
    InMux I__5710 (
            .O(N__40769),
            .I(N__40763));
    LocalMux I__5709 (
            .O(N__40766),
            .I(\reset_module_System.countZ0Z_5 ));
    LocalMux I__5708 (
            .O(N__40763),
            .I(\reset_module_System.countZ0Z_5 ));
    InMux I__5707 (
            .O(N__40758),
            .I(\reset_module_System.count_1_cry_4 ));
    InMux I__5706 (
            .O(N__40755),
            .I(N__40751));
    InMux I__5705 (
            .O(N__40754),
            .I(N__40748));
    LocalMux I__5704 (
            .O(N__40751),
            .I(\reset_module_System.countZ0Z_6 ));
    LocalMux I__5703 (
            .O(N__40748),
            .I(\reset_module_System.countZ0Z_6 ));
    InMux I__5702 (
            .O(N__40743),
            .I(\reset_module_System.count_1_cry_5 ));
    InMux I__5701 (
            .O(N__40740),
            .I(N__40736));
    InMux I__5700 (
            .O(N__40739),
            .I(N__40733));
    LocalMux I__5699 (
            .O(N__40736),
            .I(\reset_module_System.countZ0Z_7 ));
    LocalMux I__5698 (
            .O(N__40733),
            .I(\reset_module_System.countZ0Z_7 ));
    InMux I__5697 (
            .O(N__40728),
            .I(\reset_module_System.count_1_cry_6 ));
    InMux I__5696 (
            .O(N__40725),
            .I(N__40721));
    InMux I__5695 (
            .O(N__40724),
            .I(N__40718));
    LocalMux I__5694 (
            .O(N__40721),
            .I(\reset_module_System.countZ0Z_8 ));
    LocalMux I__5693 (
            .O(N__40718),
            .I(\reset_module_System.countZ0Z_8 ));
    InMux I__5692 (
            .O(N__40713),
            .I(\reset_module_System.count_1_cry_7 ));
    CascadeMux I__5691 (
            .O(N__40710),
            .I(N__40706));
    InMux I__5690 (
            .O(N__40709),
            .I(N__40703));
    InMux I__5689 (
            .O(N__40706),
            .I(N__40700));
    LocalMux I__5688 (
            .O(N__40703),
            .I(\reset_module_System.countZ0Z_9 ));
    LocalMux I__5687 (
            .O(N__40700),
            .I(\reset_module_System.countZ0Z_9 ));
    InMux I__5686 (
            .O(N__40695),
            .I(bfn_8_2_0_));
    InMux I__5685 (
            .O(N__40692),
            .I(N__40689));
    LocalMux I__5684 (
            .O(N__40689),
            .I(N__40686));
    Odrv4 I__5683 (
            .O(N__40686),
            .I(\dron_frame_decoder_1.drone_altitude_10 ));
    InMux I__5682 (
            .O(N__40683),
            .I(N__40680));
    LocalMux I__5681 (
            .O(N__40680),
            .I(drone_altitude_12));
    InMux I__5680 (
            .O(N__40677),
            .I(N__40674));
    LocalMux I__5679 (
            .O(N__40674),
            .I(drone_altitude_13));
    InMux I__5678 (
            .O(N__40671),
            .I(N__40668));
    LocalMux I__5677 (
            .O(N__40668),
            .I(drone_altitude_14));
    InMux I__5676 (
            .O(N__40665),
            .I(N__40662));
    LocalMux I__5675 (
            .O(N__40662),
            .I(N__40659));
    Odrv4 I__5674 (
            .O(N__40659),
            .I(drone_altitude_15));
    InMux I__5673 (
            .O(N__40656),
            .I(N__40653));
    LocalMux I__5672 (
            .O(N__40653),
            .I(N__40650));
    Span4Mux_h I__5671 (
            .O(N__40650),
            .I(N__40647));
    Odrv4 I__5670 (
            .O(N__40647),
            .I(\dron_frame_decoder_1.drone_altitude_8 ));
    InMux I__5669 (
            .O(N__40644),
            .I(N__40641));
    LocalMux I__5668 (
            .O(N__40641),
            .I(N__40638));
    Span4Mux_h I__5667 (
            .O(N__40638),
            .I(N__40635));
    Odrv4 I__5666 (
            .O(N__40635),
            .I(\dron_frame_decoder_1.drone_altitude_9 ));
    CascadeMux I__5665 (
            .O(N__40632),
            .I(\pid_front.N_99_cascade_ ));
    CascadeMux I__5664 (
            .O(N__40629),
            .I(N__40626));
    InMux I__5663 (
            .O(N__40626),
            .I(N__40623));
    LocalMux I__5662 (
            .O(N__40623),
            .I(N__40620));
    Span4Mux_v I__5661 (
            .O(N__40620),
            .I(N__40617));
    Odrv4 I__5660 (
            .O(N__40617),
            .I(\pid_alt.error_axbZ0Z_12 ));
    InMux I__5659 (
            .O(N__40614),
            .I(N__40611));
    LocalMux I__5658 (
            .O(N__40611),
            .I(N__40608));
    Span4Mux_h I__5657 (
            .O(N__40608),
            .I(N__40605));
    Odrv4 I__5656 (
            .O(N__40605),
            .I(\pid_alt.error_axbZ0Z_13 ));
    InMux I__5655 (
            .O(N__40602),
            .I(N__40599));
    LocalMux I__5654 (
            .O(N__40599),
            .I(N__40596));
    Span4Mux_h I__5653 (
            .O(N__40596),
            .I(N__40593));
    Odrv4 I__5652 (
            .O(N__40593),
            .I(\pid_alt.error_axbZ0Z_14 ));
    InMux I__5651 (
            .O(N__40590),
            .I(\uart_pc.un4_timer_Count_1_cry_1 ));
    InMux I__5650 (
            .O(N__40587),
            .I(\uart_pc.un4_timer_Count_1_cry_2 ));
    InMux I__5649 (
            .O(N__40584),
            .I(\uart_pc.un4_timer_Count_1_cry_3 ));
    InMux I__5648 (
            .O(N__40581),
            .I(N__40578));
    LocalMux I__5647 (
            .O(N__40578),
            .I(N__40574));
    InMux I__5646 (
            .O(N__40577),
            .I(N__40571));
    Span4Mux_v I__5645 (
            .O(N__40574),
            .I(N__40566));
    LocalMux I__5644 (
            .O(N__40571),
            .I(N__40566));
    Span4Mux_v I__5643 (
            .O(N__40566),
            .I(N__40563));
    Odrv4 I__5642 (
            .O(N__40563),
            .I(\uart_pc.N_126_li ));
    InMux I__5641 (
            .O(N__40560),
            .I(N__40556));
    InMux I__5640 (
            .O(N__40559),
            .I(N__40553));
    LocalMux I__5639 (
            .O(N__40556),
            .I(N__40546));
    LocalMux I__5638 (
            .O(N__40553),
            .I(N__40546));
    InMux I__5637 (
            .O(N__40552),
            .I(N__40543));
    InMux I__5636 (
            .O(N__40551),
            .I(N__40540));
    Span4Mux_v I__5635 (
            .O(N__40546),
            .I(N__40535));
    LocalMux I__5634 (
            .O(N__40543),
            .I(N__40535));
    LocalMux I__5633 (
            .O(N__40540),
            .I(N__40532));
    Span4Mux_v I__5632 (
            .O(N__40535),
            .I(N__40528));
    Span4Mux_v I__5631 (
            .O(N__40532),
            .I(N__40525));
    InMux I__5630 (
            .O(N__40531),
            .I(N__40522));
    Span4Mux_h I__5629 (
            .O(N__40528),
            .I(N__40514));
    Span4Mux_h I__5628 (
            .O(N__40525),
            .I(N__40514));
    LocalMux I__5627 (
            .O(N__40522),
            .I(N__40514));
    InMux I__5626 (
            .O(N__40521),
            .I(N__40511));
    Odrv4 I__5625 (
            .O(N__40514),
            .I(\uart_pc.stateZ0Z_4 ));
    LocalMux I__5624 (
            .O(N__40511),
            .I(\uart_pc.stateZ0Z_4 ));
    CascadeMux I__5623 (
            .O(N__40506),
            .I(N__40503));
    InMux I__5622 (
            .O(N__40503),
            .I(N__40500));
    LocalMux I__5621 (
            .O(N__40500),
            .I(\uart_pc.un1_state_2_0_a3_0 ));
    CascadeMux I__5620 (
            .O(N__40497),
            .I(N__40494));
    InMux I__5619 (
            .O(N__40494),
            .I(N__40482));
    InMux I__5618 (
            .O(N__40493),
            .I(N__40482));
    InMux I__5617 (
            .O(N__40492),
            .I(N__40469));
    InMux I__5616 (
            .O(N__40491),
            .I(N__40469));
    InMux I__5615 (
            .O(N__40490),
            .I(N__40469));
    InMux I__5614 (
            .O(N__40489),
            .I(N__40469));
    InMux I__5613 (
            .O(N__40488),
            .I(N__40469));
    InMux I__5612 (
            .O(N__40487),
            .I(N__40469));
    LocalMux I__5611 (
            .O(N__40482),
            .I(N__40466));
    LocalMux I__5610 (
            .O(N__40469),
            .I(N__40463));
    Span4Mux_v I__5609 (
            .O(N__40466),
            .I(N__40460));
    Span4Mux_v I__5608 (
            .O(N__40463),
            .I(N__40455));
    Span4Mux_h I__5607 (
            .O(N__40460),
            .I(N__40455));
    Sp12to4 I__5606 (
            .O(N__40455),
            .I(N__40452));
    Odrv12 I__5605 (
            .O(N__40452),
            .I(\uart_pc.un1_state_2_0 ));
    InMux I__5604 (
            .O(N__40449),
            .I(N__40446));
    LocalMux I__5603 (
            .O(N__40446),
            .I(\uart_pc.timer_Count_RNO_0Z0Z_3 ));
    InMux I__5602 (
            .O(N__40443),
            .I(N__40436));
    InMux I__5601 (
            .O(N__40442),
            .I(N__40429));
    InMux I__5600 (
            .O(N__40441),
            .I(N__40429));
    InMux I__5599 (
            .O(N__40440),
            .I(N__40429));
    CascadeMux I__5598 (
            .O(N__40439),
            .I(N__40424));
    LocalMux I__5597 (
            .O(N__40436),
            .I(N__40420));
    LocalMux I__5596 (
            .O(N__40429),
            .I(N__40417));
    InMux I__5595 (
            .O(N__40428),
            .I(N__40410));
    InMux I__5594 (
            .O(N__40427),
            .I(N__40410));
    InMux I__5593 (
            .O(N__40424),
            .I(N__40410));
    InMux I__5592 (
            .O(N__40423),
            .I(N__40407));
    Span4Mux_h I__5591 (
            .O(N__40420),
            .I(N__40402));
    Span4Mux_h I__5590 (
            .O(N__40417),
            .I(N__40402));
    LocalMux I__5589 (
            .O(N__40410),
            .I(N__40399));
    LocalMux I__5588 (
            .O(N__40407),
            .I(\uart_pc.timer_CountZ1Z_3 ));
    Odrv4 I__5587 (
            .O(N__40402),
            .I(\uart_pc.timer_CountZ1Z_3 ));
    Odrv4 I__5586 (
            .O(N__40399),
            .I(\uart_pc.timer_CountZ1Z_3 ));
    InMux I__5585 (
            .O(N__40392),
            .I(N__40389));
    LocalMux I__5584 (
            .O(N__40389),
            .I(\uart_pc.timer_Count_RNO_0Z0Z_4 ));
    InMux I__5583 (
            .O(N__40386),
            .I(N__40379));
    InMux I__5582 (
            .O(N__40385),
            .I(N__40372));
    InMux I__5581 (
            .O(N__40384),
            .I(N__40372));
    InMux I__5580 (
            .O(N__40383),
            .I(N__40372));
    InMux I__5579 (
            .O(N__40382),
            .I(N__40366));
    LocalMux I__5578 (
            .O(N__40379),
            .I(N__40362));
    LocalMux I__5577 (
            .O(N__40372),
            .I(N__40359));
    InMux I__5576 (
            .O(N__40371),
            .I(N__40352));
    InMux I__5575 (
            .O(N__40370),
            .I(N__40352));
    InMux I__5574 (
            .O(N__40369),
            .I(N__40352));
    LocalMux I__5573 (
            .O(N__40366),
            .I(N__40349));
    InMux I__5572 (
            .O(N__40365),
            .I(N__40346));
    Span4Mux_h I__5571 (
            .O(N__40362),
            .I(N__40341));
    Span4Mux_h I__5570 (
            .O(N__40359),
            .I(N__40341));
    LocalMux I__5569 (
            .O(N__40352),
            .I(N__40338));
    Odrv12 I__5568 (
            .O(N__40349),
            .I(\uart_pc.timer_CountZ0Z_4 ));
    LocalMux I__5567 (
            .O(N__40346),
            .I(\uart_pc.timer_CountZ0Z_4 ));
    Odrv4 I__5566 (
            .O(N__40341),
            .I(\uart_pc.timer_CountZ0Z_4 ));
    Odrv4 I__5565 (
            .O(N__40338),
            .I(\uart_pc.timer_CountZ0Z_4 ));
    InMux I__5564 (
            .O(N__40329),
            .I(N__40326));
    LocalMux I__5563 (
            .O(N__40326),
            .I(\uart_pc.timer_Count_RNO_0Z0Z_2 ));
    CascadeMux I__5562 (
            .O(N__40323),
            .I(N__40319));
    InMux I__5561 (
            .O(N__40322),
            .I(N__40316));
    InMux I__5560 (
            .O(N__40319),
            .I(N__40313));
    LocalMux I__5559 (
            .O(N__40316),
            .I(N__40309));
    LocalMux I__5558 (
            .O(N__40313),
            .I(N__40306));
    InMux I__5557 (
            .O(N__40312),
            .I(N__40303));
    Span4Mux_h I__5556 (
            .O(N__40309),
            .I(N__40298));
    Span4Mux_h I__5555 (
            .O(N__40306),
            .I(N__40298));
    LocalMux I__5554 (
            .O(N__40303),
            .I(\uart_pc.timer_CountZ1Z_2 ));
    Odrv4 I__5553 (
            .O(N__40298),
            .I(\uart_pc.timer_CountZ1Z_2 ));
    InMux I__5552 (
            .O(N__40293),
            .I(N__40290));
    LocalMux I__5551 (
            .O(N__40290),
            .I(N__40287));
    Span4Mux_v I__5550 (
            .O(N__40287),
            .I(N__40284));
    Span4Mux_v I__5549 (
            .O(N__40284),
            .I(N__40280));
    InMux I__5548 (
            .O(N__40283),
            .I(N__40277));
    Span4Mux_h I__5547 (
            .O(N__40280),
            .I(N__40274));
    LocalMux I__5546 (
            .O(N__40277),
            .I(N__40271));
    Odrv4 I__5545 (
            .O(N__40274),
            .I(\Commands_frame_decoder.source_offset4data_1_sqmuxa ));
    Odrv12 I__5544 (
            .O(N__40271),
            .I(\Commands_frame_decoder.source_offset4data_1_sqmuxa ));
    CascadeMux I__5543 (
            .O(N__40266),
            .I(\uart_pc.un1_state_4_0_cascade_ ));
    CascadeMux I__5542 (
            .O(N__40263),
            .I(N__40260));
    InMux I__5541 (
            .O(N__40260),
            .I(N__40257));
    LocalMux I__5540 (
            .O(N__40257),
            .I(\uart_pc.CO0 ));
    IoInMux I__5539 (
            .O(N__40254),
            .I(N__40251));
    LocalMux I__5538 (
            .O(N__40251),
            .I(N__40247));
    InMux I__5537 (
            .O(N__40250),
            .I(N__40244));
    Span4Mux_s1_v I__5536 (
            .O(N__40247),
            .I(N__40234));
    LocalMux I__5535 (
            .O(N__40244),
            .I(N__40231));
    InMux I__5534 (
            .O(N__40243),
            .I(N__40228));
    CascadeMux I__5533 (
            .O(N__40242),
            .I(N__40225));
    CascadeMux I__5532 (
            .O(N__40241),
            .I(N__40222));
    CascadeMux I__5531 (
            .O(N__40240),
            .I(N__40219));
    CascadeMux I__5530 (
            .O(N__40239),
            .I(N__40216));
    InMux I__5529 (
            .O(N__40238),
            .I(N__40209));
    InMux I__5528 (
            .O(N__40237),
            .I(N__40206));
    Span4Mux_v I__5527 (
            .O(N__40234),
            .I(N__40202));
    Span4Mux_v I__5526 (
            .O(N__40231),
            .I(N__40197));
    LocalMux I__5525 (
            .O(N__40228),
            .I(N__40197));
    InMux I__5524 (
            .O(N__40225),
            .I(N__40180));
    InMux I__5523 (
            .O(N__40222),
            .I(N__40180));
    InMux I__5522 (
            .O(N__40219),
            .I(N__40180));
    InMux I__5521 (
            .O(N__40216),
            .I(N__40180));
    InMux I__5520 (
            .O(N__40215),
            .I(N__40180));
    InMux I__5519 (
            .O(N__40214),
            .I(N__40180));
    InMux I__5518 (
            .O(N__40213),
            .I(N__40180));
    InMux I__5517 (
            .O(N__40212),
            .I(N__40180));
    LocalMux I__5516 (
            .O(N__40209),
            .I(N__40177));
    LocalMux I__5515 (
            .O(N__40206),
            .I(N__40174));
    InMux I__5514 (
            .O(N__40205),
            .I(N__40171));
    Span4Mux_h I__5513 (
            .O(N__40202),
            .I(N__40168));
    Span4Mux_h I__5512 (
            .O(N__40197),
            .I(N__40165));
    LocalMux I__5511 (
            .O(N__40180),
            .I(N__40156));
    Span4Mux_v I__5510 (
            .O(N__40177),
            .I(N__40156));
    Span4Mux_h I__5509 (
            .O(N__40174),
            .I(N__40156));
    LocalMux I__5508 (
            .O(N__40171),
            .I(N__40156));
    Span4Mux_h I__5507 (
            .O(N__40168),
            .I(N__40151));
    Span4Mux_v I__5506 (
            .O(N__40165),
            .I(N__40151));
    Span4Mux_v I__5505 (
            .O(N__40156),
            .I(N__40148));
    Odrv4 I__5504 (
            .O(N__40151),
            .I(debug_CH2_18A_c));
    Odrv4 I__5503 (
            .O(N__40148),
            .I(debug_CH2_18A_c));
    CascadeMux I__5502 (
            .O(N__40143),
            .I(N__40139));
    InMux I__5501 (
            .O(N__40142),
            .I(N__40133));
    InMux I__5500 (
            .O(N__40139),
            .I(N__40133));
    InMux I__5499 (
            .O(N__40138),
            .I(N__40130));
    LocalMux I__5498 (
            .O(N__40133),
            .I(N__40127));
    LocalMux I__5497 (
            .O(N__40130),
            .I(\uart_pc.stateZ0Z_1 ));
    Odrv4 I__5496 (
            .O(N__40127),
            .I(\uart_pc.stateZ0Z_1 ));
    CascadeMux I__5495 (
            .O(N__40122),
            .I(\uart_pc.state_srsts_i_0_2_cascade_ ));
    CascadeMux I__5494 (
            .O(N__40119),
            .I(N__40115));
    InMux I__5493 (
            .O(N__40118),
            .I(N__40111));
    InMux I__5492 (
            .O(N__40115),
            .I(N__40108));
    InMux I__5491 (
            .O(N__40114),
            .I(N__40104));
    LocalMux I__5490 (
            .O(N__40111),
            .I(N__40099));
    LocalMux I__5489 (
            .O(N__40108),
            .I(N__40099));
    InMux I__5488 (
            .O(N__40107),
            .I(N__40096));
    LocalMux I__5487 (
            .O(N__40104),
            .I(\uart_pc.stateZ0Z_2 ));
    Odrv4 I__5486 (
            .O(N__40099),
            .I(\uart_pc.stateZ0Z_2 ));
    LocalMux I__5485 (
            .O(N__40096),
            .I(\uart_pc.stateZ0Z_2 ));
    InMux I__5484 (
            .O(N__40089),
            .I(N__40086));
    LocalMux I__5483 (
            .O(N__40086),
            .I(N__40082));
    InMux I__5482 (
            .O(N__40085),
            .I(N__40079));
    Span4Mux_v I__5481 (
            .O(N__40082),
            .I(N__40076));
    LocalMux I__5480 (
            .O(N__40079),
            .I(\uart_pc.timer_CountZ1Z_1 ));
    Odrv4 I__5479 (
            .O(N__40076),
            .I(\uart_pc.timer_CountZ1Z_1 ));
    CascadeMux I__5478 (
            .O(N__40071),
            .I(N__40066));
    InMux I__5477 (
            .O(N__40070),
            .I(N__40063));
    InMux I__5476 (
            .O(N__40069),
            .I(N__40058));
    InMux I__5475 (
            .O(N__40066),
            .I(N__40058));
    LocalMux I__5474 (
            .O(N__40063),
            .I(N__40053));
    LocalMux I__5473 (
            .O(N__40058),
            .I(N__40053));
    Odrv4 I__5472 (
            .O(N__40053),
            .I(\uart_drone.N_126_li ));
    CascadeMux I__5471 (
            .O(N__40050),
            .I(N__40047));
    InMux I__5470 (
            .O(N__40047),
            .I(N__40044));
    LocalMux I__5469 (
            .O(N__40044),
            .I(N__40041));
    Span4Mux_v I__5468 (
            .O(N__40041),
            .I(N__40038));
    Odrv4 I__5467 (
            .O(N__40038),
            .I(\uart_drone.un1_state_2_0_a3_0 ));
    CascadeMux I__5466 (
            .O(N__40035),
            .I(N__40032));
    InMux I__5465 (
            .O(N__40032),
            .I(N__40028));
    InMux I__5464 (
            .O(N__40031),
            .I(N__40025));
    LocalMux I__5463 (
            .O(N__40028),
            .I(\uart_pc.stateZ0Z_0 ));
    LocalMux I__5462 (
            .O(N__40025),
            .I(\uart_pc.stateZ0Z_0 ));
    InMux I__5461 (
            .O(N__40020),
            .I(N__40014));
    InMux I__5460 (
            .O(N__40019),
            .I(N__40014));
    LocalMux I__5459 (
            .O(N__40014),
            .I(N__40011));
    Odrv4 I__5458 (
            .O(N__40011),
            .I(\uart_pc.un1_state_7_0 ));
    CascadeMux I__5457 (
            .O(N__40008),
            .I(N__40002));
    CascadeMux I__5456 (
            .O(N__40007),
            .I(N__39998));
    CascadeMux I__5455 (
            .O(N__40006),
            .I(N__39994));
    InMux I__5454 (
            .O(N__40005),
            .I(N__39976));
    InMux I__5453 (
            .O(N__40002),
            .I(N__39976));
    InMux I__5452 (
            .O(N__40001),
            .I(N__39976));
    InMux I__5451 (
            .O(N__39998),
            .I(N__39976));
    InMux I__5450 (
            .O(N__39997),
            .I(N__39976));
    InMux I__5449 (
            .O(N__39994),
            .I(N__39976));
    InMux I__5448 (
            .O(N__39993),
            .I(N__39976));
    InMux I__5447 (
            .O(N__39992),
            .I(N__39971));
    InMux I__5446 (
            .O(N__39991),
            .I(N__39971));
    LocalMux I__5445 (
            .O(N__39976),
            .I(N__39968));
    LocalMux I__5444 (
            .O(N__39971),
            .I(N__39962));
    Span4Mux_v I__5443 (
            .O(N__39968),
            .I(N__39962));
    InMux I__5442 (
            .O(N__39967),
            .I(N__39959));
    Odrv4 I__5441 (
            .O(N__39962),
            .I(\uart_pc.bit_CountZ0Z_1 ));
    LocalMux I__5440 (
            .O(N__39959),
            .I(\uart_pc.bit_CountZ0Z_1 ));
    InMux I__5439 (
            .O(N__39954),
            .I(N__39933));
    InMux I__5438 (
            .O(N__39953),
            .I(N__39933));
    InMux I__5437 (
            .O(N__39952),
            .I(N__39933));
    InMux I__5436 (
            .O(N__39951),
            .I(N__39933));
    InMux I__5435 (
            .O(N__39950),
            .I(N__39933));
    InMux I__5434 (
            .O(N__39949),
            .I(N__39933));
    InMux I__5433 (
            .O(N__39948),
            .I(N__39933));
    LocalMux I__5432 (
            .O(N__39933),
            .I(N__39929));
    InMux I__5431 (
            .O(N__39932),
            .I(N__39925));
    Span4Mux_v I__5430 (
            .O(N__39929),
            .I(N__39922));
    InMux I__5429 (
            .O(N__39928),
            .I(N__39919));
    LocalMux I__5428 (
            .O(N__39925),
            .I(\uart_pc.bit_CountZ0Z_2 ));
    Odrv4 I__5427 (
            .O(N__39922),
            .I(\uart_pc.bit_CountZ0Z_2 ));
    LocalMux I__5426 (
            .O(N__39919),
            .I(\uart_pc.bit_CountZ0Z_2 ));
    SRMux I__5425 (
            .O(N__39912),
            .I(N__39909));
    LocalMux I__5424 (
            .O(N__39909),
            .I(N__39906));
    Span4Mux_h I__5423 (
            .O(N__39906),
            .I(N__39903));
    Span4Mux_v I__5422 (
            .O(N__39903),
            .I(N__39900));
    Odrv4 I__5421 (
            .O(N__39900),
            .I(\uart_pc.state_RNIEAGSZ0Z_4 ));
    InMux I__5420 (
            .O(N__39897),
            .I(N__39893));
    InMux I__5419 (
            .O(N__39896),
            .I(N__39890));
    LocalMux I__5418 (
            .O(N__39893),
            .I(N__39887));
    LocalMux I__5417 (
            .O(N__39890),
            .I(N__39884));
    Span4Mux_v I__5416 (
            .O(N__39887),
            .I(N__39881));
    Span4Mux_v I__5415 (
            .O(N__39884),
            .I(N__39876));
    Span4Mux_h I__5414 (
            .O(N__39881),
            .I(N__39876));
    Odrv4 I__5413 (
            .O(N__39876),
            .I(\Commands_frame_decoder.source_xy_ki_1_sqmuxa ));
    CascadeMux I__5412 (
            .O(N__39873),
            .I(N__39869));
    InMux I__5411 (
            .O(N__39872),
            .I(N__39860));
    InMux I__5410 (
            .O(N__39869),
            .I(N__39860));
    InMux I__5409 (
            .O(N__39868),
            .I(N__39860));
    InMux I__5408 (
            .O(N__39867),
            .I(N__39857));
    LocalMux I__5407 (
            .O(N__39860),
            .I(N__39854));
    LocalMux I__5406 (
            .O(N__39857),
            .I(\uart_drone.timer_CountZ0Z_0 ));
    Odrv4 I__5405 (
            .O(N__39854),
            .I(\uart_drone.timer_CountZ0Z_0 ));
    InMux I__5404 (
            .O(N__39849),
            .I(N__39846));
    LocalMux I__5403 (
            .O(N__39846),
            .I(N__39843));
    Odrv4 I__5402 (
            .O(N__39843),
            .I(\uart_drone.timer_Count_RNO_0_0_3 ));
    CascadeMux I__5401 (
            .O(N__39840),
            .I(N__39836));
    InMux I__5400 (
            .O(N__39839),
            .I(N__39830));
    InMux I__5399 (
            .O(N__39836),
            .I(N__39830));
    InMux I__5398 (
            .O(N__39835),
            .I(N__39827));
    LocalMux I__5397 (
            .O(N__39830),
            .I(N__39824));
    LocalMux I__5396 (
            .O(N__39827),
            .I(N__39819));
    Span4Mux_h I__5395 (
            .O(N__39824),
            .I(N__39819));
    Odrv4 I__5394 (
            .O(N__39819),
            .I(\uart_drone.timer_CountZ1Z_2 ));
    InMux I__5393 (
            .O(N__39816),
            .I(N__39813));
    LocalMux I__5392 (
            .O(N__39813),
            .I(N__39807));
    InMux I__5391 (
            .O(N__39812),
            .I(N__39802));
    InMux I__5390 (
            .O(N__39811),
            .I(N__39802));
    InMux I__5389 (
            .O(N__39810),
            .I(N__39799));
    Span4Mux_v I__5388 (
            .O(N__39807),
            .I(N__39792));
    LocalMux I__5387 (
            .O(N__39802),
            .I(N__39792));
    LocalMux I__5386 (
            .O(N__39799),
            .I(N__39789));
    InMux I__5385 (
            .O(N__39798),
            .I(N__39784));
    InMux I__5384 (
            .O(N__39797),
            .I(N__39784));
    Odrv4 I__5383 (
            .O(N__39792),
            .I(\uart_drone.N_143 ));
    Odrv4 I__5382 (
            .O(N__39789),
            .I(\uart_drone.N_143 ));
    LocalMux I__5381 (
            .O(N__39784),
            .I(\uart_drone.N_143 ));
    CascadeMux I__5380 (
            .O(N__39777),
            .I(N__39771));
    CascadeMux I__5379 (
            .O(N__39776),
            .I(N__39768));
    CascadeMux I__5378 (
            .O(N__39775),
            .I(N__39764));
    CascadeMux I__5377 (
            .O(N__39774),
            .I(N__39761));
    InMux I__5376 (
            .O(N__39771),
            .I(N__39756));
    InMux I__5375 (
            .O(N__39768),
            .I(N__39756));
    InMux I__5374 (
            .O(N__39767),
            .I(N__39753));
    InMux I__5373 (
            .O(N__39764),
            .I(N__39748));
    InMux I__5372 (
            .O(N__39761),
            .I(N__39748));
    LocalMux I__5371 (
            .O(N__39756),
            .I(N__39745));
    LocalMux I__5370 (
            .O(N__39753),
            .I(N__39742));
    LocalMux I__5369 (
            .O(N__39748),
            .I(N__39737));
    Span4Mux_h I__5368 (
            .O(N__39745),
            .I(N__39737));
    Span4Mux_h I__5367 (
            .O(N__39742),
            .I(N__39734));
    Odrv4 I__5366 (
            .O(N__39737),
            .I(\uart_drone.timer_Count_0_sqmuxa ));
    Odrv4 I__5365 (
            .O(N__39734),
            .I(\uart_drone.timer_Count_0_sqmuxa ));
    CascadeMux I__5364 (
            .O(N__39729),
            .I(\uart_pc.state_srsts_0_0_0_cascade_ ));
    InMux I__5363 (
            .O(N__39726),
            .I(N__39723));
    LocalMux I__5362 (
            .O(N__39723),
            .I(N__39720));
    Odrv4 I__5361 (
            .O(N__39720),
            .I(\uart_pc_sync.aux_3__0_Z0Z_0 ));
    InMux I__5360 (
            .O(N__39717),
            .I(N__39714));
    LocalMux I__5359 (
            .O(N__39714),
            .I(\uart_pc_sync.aux_1__0_Z0Z_0 ));
    InMux I__5358 (
            .O(N__39711),
            .I(N__39708));
    LocalMux I__5357 (
            .O(N__39708),
            .I(\uart_pc_sync.aux_2__0_Z0Z_0 ));
    CascadeMux I__5356 (
            .O(N__39705),
            .I(\uart_drone.state_srsts_0_0_0_cascade_ ));
    InMux I__5355 (
            .O(N__39702),
            .I(N__39696));
    InMux I__5354 (
            .O(N__39701),
            .I(N__39696));
    LocalMux I__5353 (
            .O(N__39696),
            .I(\uart_drone.stateZ0Z_0 ));
    InMux I__5352 (
            .O(N__39693),
            .I(N__39688));
    InMux I__5351 (
            .O(N__39692),
            .I(N__39683));
    InMux I__5350 (
            .O(N__39691),
            .I(N__39683));
    LocalMux I__5349 (
            .O(N__39688),
            .I(\uart_drone.stateZ0Z_1 ));
    LocalMux I__5348 (
            .O(N__39683),
            .I(\uart_drone.stateZ0Z_1 ));
    CascadeMux I__5347 (
            .O(N__39678),
            .I(\uart_drone.state_srsts_i_0_2_cascade_ ));
    InMux I__5346 (
            .O(N__39675),
            .I(N__39672));
    LocalMux I__5345 (
            .O(N__39672),
            .I(\reset_module_System.reset6_13 ));
    CascadeMux I__5344 (
            .O(N__39669),
            .I(\reset_module_System.reset6_17_cascade_ ));
    InMux I__5343 (
            .O(N__39666),
            .I(N__39663));
    LocalMux I__5342 (
            .O(N__39663),
            .I(\reset_module_System.reset6_11 ));
    CascadeMux I__5341 (
            .O(N__39660),
            .I(\reset_module_System.reset6_19_cascade_ ));
    InMux I__5340 (
            .O(N__39657),
            .I(N__39654));
    LocalMux I__5339 (
            .O(N__39654),
            .I(N__39651));
    Span4Mux_h I__5338 (
            .O(N__39651),
            .I(N__39648));
    Span4Mux_v I__5337 (
            .O(N__39648),
            .I(N__39645));
    Odrv4 I__5336 (
            .O(N__39645),
            .I(scaler_4_data_5));
    InMux I__5335 (
            .O(N__39642),
            .I(N__39639));
    LocalMux I__5334 (
            .O(N__39639),
            .I(N__39636));
    Span12Mux_s9_h I__5333 (
            .O(N__39636),
            .I(N__39633));
    Odrv12 I__5332 (
            .O(N__39633),
            .I(uart_input_pc_c));
    InMux I__5331 (
            .O(N__39630),
            .I(N__39627));
    LocalMux I__5330 (
            .O(N__39627),
            .I(\uart_pc_sync.aux_0__0_Z0Z_0 ));
    InMux I__5329 (
            .O(N__39624),
            .I(N__39621));
    LocalMux I__5328 (
            .O(N__39621),
            .I(N__39617));
    InMux I__5327 (
            .O(N__39620),
            .I(N__39614));
    Span4Mux_h I__5326 (
            .O(N__39617),
            .I(N__39611));
    LocalMux I__5325 (
            .O(N__39614),
            .I(\pid_alt.error_i_acummZ0Z_11 ));
    Odrv4 I__5324 (
            .O(N__39611),
            .I(\pid_alt.error_i_acummZ0Z_11 ));
    InMux I__5323 (
            .O(N__39606),
            .I(N__39601));
    InMux I__5322 (
            .O(N__39605),
            .I(N__39598));
    InMux I__5321 (
            .O(N__39604),
            .I(N__39595));
    LocalMux I__5320 (
            .O(N__39601),
            .I(N__39592));
    LocalMux I__5319 (
            .O(N__39598),
            .I(N__39589));
    LocalMux I__5318 (
            .O(N__39595),
            .I(N__39586));
    Span4Mux_v I__5317 (
            .O(N__39592),
            .I(N__39581));
    Span4Mux_v I__5316 (
            .O(N__39589),
            .I(N__39581));
    Odrv4 I__5315 (
            .O(N__39586),
            .I(\pid_alt.error_i_acumm_preregZ0Z_6 ));
    Odrv4 I__5314 (
            .O(N__39581),
            .I(\pid_alt.error_i_acumm_preregZ0Z_6 ));
    InMux I__5313 (
            .O(N__39576),
            .I(N__39573));
    LocalMux I__5312 (
            .O(N__39573),
            .I(N__39569));
    InMux I__5311 (
            .O(N__39572),
            .I(N__39566));
    Span4Mux_h I__5310 (
            .O(N__39569),
            .I(N__39563));
    LocalMux I__5309 (
            .O(N__39566),
            .I(\pid_alt.error_i_acummZ0Z_6 ));
    Odrv4 I__5308 (
            .O(N__39563),
            .I(\pid_alt.error_i_acummZ0Z_6 ));
    InMux I__5307 (
            .O(N__39558),
            .I(N__39553));
    InMux I__5306 (
            .O(N__39557),
            .I(N__39550));
    CascadeMux I__5305 (
            .O(N__39556),
            .I(N__39547));
    LocalMux I__5304 (
            .O(N__39553),
            .I(N__39544));
    LocalMux I__5303 (
            .O(N__39550),
            .I(N__39541));
    InMux I__5302 (
            .O(N__39547),
            .I(N__39538));
    Span4Mux_v I__5301 (
            .O(N__39544),
            .I(N__39535));
    Span4Mux_h I__5300 (
            .O(N__39541),
            .I(N__39532));
    LocalMux I__5299 (
            .O(N__39538),
            .I(N__39529));
    Odrv4 I__5298 (
            .O(N__39535),
            .I(\pid_alt.error_i_acumm_preregZ0Z_7 ));
    Odrv4 I__5297 (
            .O(N__39532),
            .I(\pid_alt.error_i_acumm_preregZ0Z_7 ));
    Odrv4 I__5296 (
            .O(N__39529),
            .I(\pid_alt.error_i_acumm_preregZ0Z_7 ));
    InMux I__5295 (
            .O(N__39522),
            .I(N__39519));
    LocalMux I__5294 (
            .O(N__39519),
            .I(N__39515));
    InMux I__5293 (
            .O(N__39518),
            .I(N__39512));
    Span4Mux_h I__5292 (
            .O(N__39515),
            .I(N__39509));
    LocalMux I__5291 (
            .O(N__39512),
            .I(\pid_alt.error_i_acummZ0Z_7 ));
    Odrv4 I__5290 (
            .O(N__39509),
            .I(\pid_alt.error_i_acummZ0Z_7 ));
    InMux I__5289 (
            .O(N__39504),
            .I(N__39501));
    LocalMux I__5288 (
            .O(N__39501),
            .I(N__39496));
    InMux I__5287 (
            .O(N__39500),
            .I(N__39493));
    InMux I__5286 (
            .O(N__39499),
            .I(N__39490));
    Span4Mux_v I__5285 (
            .O(N__39496),
            .I(N__39487));
    LocalMux I__5284 (
            .O(N__39493),
            .I(\pid_alt.error_i_acumm_preregZ0Z_8 ));
    LocalMux I__5283 (
            .O(N__39490),
            .I(\pid_alt.error_i_acumm_preregZ0Z_8 ));
    Odrv4 I__5282 (
            .O(N__39487),
            .I(\pid_alt.error_i_acumm_preregZ0Z_8 ));
    InMux I__5281 (
            .O(N__39480),
            .I(N__39476));
    CascadeMux I__5280 (
            .O(N__39479),
            .I(N__39473));
    LocalMux I__5279 (
            .O(N__39476),
            .I(N__39470));
    InMux I__5278 (
            .O(N__39473),
            .I(N__39467));
    Span4Mux_h I__5277 (
            .O(N__39470),
            .I(N__39464));
    LocalMux I__5276 (
            .O(N__39467),
            .I(\pid_alt.error_i_acummZ0Z_8 ));
    Odrv4 I__5275 (
            .O(N__39464),
            .I(\pid_alt.error_i_acummZ0Z_8 ));
    CascadeMux I__5274 (
            .O(N__39459),
            .I(N__39455));
    CascadeMux I__5273 (
            .O(N__39458),
            .I(N__39452));
    InMux I__5272 (
            .O(N__39455),
            .I(N__39443));
    InMux I__5271 (
            .O(N__39452),
            .I(N__39443));
    InMux I__5270 (
            .O(N__39451),
            .I(N__39434));
    InMux I__5269 (
            .O(N__39450),
            .I(N__39434));
    InMux I__5268 (
            .O(N__39449),
            .I(N__39434));
    InMux I__5267 (
            .O(N__39448),
            .I(N__39434));
    LocalMux I__5266 (
            .O(N__39443),
            .I(N__39426));
    LocalMux I__5265 (
            .O(N__39434),
            .I(N__39426));
    InMux I__5264 (
            .O(N__39433),
            .I(N__39419));
    InMux I__5263 (
            .O(N__39432),
            .I(N__39419));
    InMux I__5262 (
            .O(N__39431),
            .I(N__39419));
    Span4Mux_v I__5261 (
            .O(N__39426),
            .I(N__39414));
    LocalMux I__5260 (
            .O(N__39419),
            .I(N__39414));
    Odrv4 I__5259 (
            .O(N__39414),
            .I(\pid_alt.N_158 ));
    InMux I__5258 (
            .O(N__39411),
            .I(N__39407));
    InMux I__5257 (
            .O(N__39410),
            .I(N__39404));
    LocalMux I__5256 (
            .O(N__39407),
            .I(N__39399));
    LocalMux I__5255 (
            .O(N__39404),
            .I(N__39399));
    Span4Mux_h I__5254 (
            .O(N__39399),
            .I(N__39395));
    InMux I__5253 (
            .O(N__39398),
            .I(N__39392));
    Odrv4 I__5252 (
            .O(N__39395),
            .I(\pid_alt.error_i_acumm_preregZ0Z_9 ));
    LocalMux I__5251 (
            .O(N__39392),
            .I(\pid_alt.error_i_acumm_preregZ0Z_9 ));
    InMux I__5250 (
            .O(N__39387),
            .I(N__39383));
    InMux I__5249 (
            .O(N__39386),
            .I(N__39380));
    LocalMux I__5248 (
            .O(N__39383),
            .I(N__39377));
    LocalMux I__5247 (
            .O(N__39380),
            .I(N__39372));
    Span4Mux_h I__5246 (
            .O(N__39377),
            .I(N__39372));
    Odrv4 I__5245 (
            .O(N__39372),
            .I(\pid_alt.error_i_acummZ0Z_9 ));
    InMux I__5244 (
            .O(N__39369),
            .I(N__39365));
    InMux I__5243 (
            .O(N__39368),
            .I(N__39362));
    LocalMux I__5242 (
            .O(N__39365),
            .I(N__39358));
    LocalMux I__5241 (
            .O(N__39362),
            .I(N__39355));
    InMux I__5240 (
            .O(N__39361),
            .I(N__39352));
    Span4Mux_h I__5239 (
            .O(N__39358),
            .I(N__39349));
    Odrv4 I__5238 (
            .O(N__39355),
            .I(\pid_alt.error_i_acumm7lto12 ));
    LocalMux I__5237 (
            .O(N__39352),
            .I(\pid_alt.error_i_acumm7lto12 ));
    Odrv4 I__5236 (
            .O(N__39349),
            .I(\pid_alt.error_i_acumm7lto12 ));
    InMux I__5235 (
            .O(N__39342),
            .I(N__39338));
    InMux I__5234 (
            .O(N__39341),
            .I(N__39335));
    LocalMux I__5233 (
            .O(N__39338),
            .I(\pid_alt.N_9_0 ));
    LocalMux I__5232 (
            .O(N__39335),
            .I(\pid_alt.N_9_0 ));
    InMux I__5231 (
            .O(N__39330),
            .I(N__39326));
    CascadeMux I__5230 (
            .O(N__39329),
            .I(N__39323));
    LocalMux I__5229 (
            .O(N__39326),
            .I(N__39320));
    InMux I__5228 (
            .O(N__39323),
            .I(N__39317));
    Span4Mux_h I__5227 (
            .O(N__39320),
            .I(N__39314));
    LocalMux I__5226 (
            .O(N__39317),
            .I(\pid_alt.error_i_acummZ0Z_12 ));
    Odrv4 I__5225 (
            .O(N__39314),
            .I(\pid_alt.error_i_acummZ0Z_12 ));
    InMux I__5224 (
            .O(N__39309),
            .I(N__39304));
    InMux I__5223 (
            .O(N__39308),
            .I(N__39299));
    InMux I__5222 (
            .O(N__39307),
            .I(N__39299));
    LocalMux I__5221 (
            .O(N__39304),
            .I(N__39295));
    LocalMux I__5220 (
            .O(N__39299),
            .I(N__39292));
    InMux I__5219 (
            .O(N__39298),
            .I(N__39280));
    Span12Mux_h I__5218 (
            .O(N__39295),
            .I(N__39277));
    Span4Mux_h I__5217 (
            .O(N__39292),
            .I(N__39274));
    InMux I__5216 (
            .O(N__39291),
            .I(N__39271));
    InMux I__5215 (
            .O(N__39290),
            .I(N__39264));
    InMux I__5214 (
            .O(N__39289),
            .I(N__39264));
    InMux I__5213 (
            .O(N__39288),
            .I(N__39264));
    InMux I__5212 (
            .O(N__39287),
            .I(N__39253));
    InMux I__5211 (
            .O(N__39286),
            .I(N__39253));
    InMux I__5210 (
            .O(N__39285),
            .I(N__39253));
    InMux I__5209 (
            .O(N__39284),
            .I(N__39253));
    InMux I__5208 (
            .O(N__39283),
            .I(N__39253));
    LocalMux I__5207 (
            .O(N__39280),
            .I(\Commands_frame_decoder.N_403 ));
    Odrv12 I__5206 (
            .O(N__39277),
            .I(\Commands_frame_decoder.N_403 ));
    Odrv4 I__5205 (
            .O(N__39274),
            .I(\Commands_frame_decoder.N_403 ));
    LocalMux I__5204 (
            .O(N__39271),
            .I(\Commands_frame_decoder.N_403 ));
    LocalMux I__5203 (
            .O(N__39264),
            .I(\Commands_frame_decoder.N_403 ));
    LocalMux I__5202 (
            .O(N__39253),
            .I(\Commands_frame_decoder.N_403 ));
    InMux I__5201 (
            .O(N__39240),
            .I(N__39236));
    InMux I__5200 (
            .O(N__39239),
            .I(N__39233));
    LocalMux I__5199 (
            .O(N__39236),
            .I(N__39230));
    LocalMux I__5198 (
            .O(N__39233),
            .I(N__39227));
    Span4Mux_h I__5197 (
            .O(N__39230),
            .I(N__39224));
    Span4Mux_h I__5196 (
            .O(N__39227),
            .I(N__39221));
    Sp12to4 I__5195 (
            .O(N__39224),
            .I(N__39217));
    Span4Mux_v I__5194 (
            .O(N__39221),
            .I(N__39214));
    InMux I__5193 (
            .O(N__39220),
            .I(N__39211));
    Span12Mux_v I__5192 (
            .O(N__39217),
            .I(N__39208));
    Span4Mux_v I__5191 (
            .O(N__39214),
            .I(N__39205));
    LocalMux I__5190 (
            .O(N__39211),
            .I(\Commands_frame_decoder.stateZ0Z_10 ));
    Odrv12 I__5189 (
            .O(N__39208),
            .I(\Commands_frame_decoder.stateZ0Z_10 ));
    Odrv4 I__5188 (
            .O(N__39205),
            .I(\Commands_frame_decoder.stateZ0Z_10 ));
    InMux I__5187 (
            .O(N__39198),
            .I(N__39195));
    LocalMux I__5186 (
            .O(N__39195),
            .I(N__39192));
    Span4Mux_v I__5185 (
            .O(N__39192),
            .I(N__39189));
    Span4Mux_s1_h I__5184 (
            .O(N__39189),
            .I(N__39186));
    Span4Mux_h I__5183 (
            .O(N__39186),
            .I(N__39183));
    Odrv4 I__5182 (
            .O(N__39183),
            .I(alt_kp_6));
    InMux I__5181 (
            .O(N__39180),
            .I(N__39177));
    LocalMux I__5180 (
            .O(N__39177),
            .I(N__39174));
    Span4Mux_v I__5179 (
            .O(N__39174),
            .I(N__39171));
    Span4Mux_h I__5178 (
            .O(N__39171),
            .I(N__39168));
    Odrv4 I__5177 (
            .O(N__39168),
            .I(alt_kp_7));
    CEMux I__5176 (
            .O(N__39165),
            .I(N__39162));
    LocalMux I__5175 (
            .O(N__39162),
            .I(N__39159));
    Span4Mux_v I__5174 (
            .O(N__39159),
            .I(N__39156));
    Span4Mux_v I__5173 (
            .O(N__39156),
            .I(N__39153));
    Span4Mux_v I__5172 (
            .O(N__39153),
            .I(N__39150));
    Odrv4 I__5171 (
            .O(N__39150),
            .I(\Commands_frame_decoder.state_RNIF38SZ0Z_6 ));
    InMux I__5170 (
            .O(N__39147),
            .I(N__39144));
    LocalMux I__5169 (
            .O(N__39144),
            .I(drone_altitude_i_10));
    CascadeMux I__5168 (
            .O(N__39141),
            .I(N__39138));
    InMux I__5167 (
            .O(N__39138),
            .I(N__39135));
    LocalMux I__5166 (
            .O(N__39135),
            .I(alt_command_4));
    CascadeMux I__5165 (
            .O(N__39132),
            .I(N__39129));
    InMux I__5164 (
            .O(N__39129),
            .I(N__39126));
    LocalMux I__5163 (
            .O(N__39126),
            .I(alt_command_5));
    CascadeMux I__5162 (
            .O(N__39123),
            .I(N__39120));
    InMux I__5161 (
            .O(N__39120),
            .I(N__39117));
    LocalMux I__5160 (
            .O(N__39117),
            .I(alt_command_6));
    CascadeMux I__5159 (
            .O(N__39114),
            .I(N__39111));
    InMux I__5158 (
            .O(N__39111),
            .I(N__39108));
    LocalMux I__5157 (
            .O(N__39108),
            .I(alt_command_7));
    CEMux I__5156 (
            .O(N__39105),
            .I(N__39102));
    LocalMux I__5155 (
            .O(N__39102),
            .I(N__39099));
    Odrv12 I__5154 (
            .O(N__39099),
            .I(\Commands_frame_decoder.un1_sink_data_valid_2_0_0 ));
    InMux I__5153 (
            .O(N__39096),
            .I(N__39091));
    InMux I__5152 (
            .O(N__39095),
            .I(N__39088));
    InMux I__5151 (
            .O(N__39094),
            .I(N__39085));
    LocalMux I__5150 (
            .O(N__39091),
            .I(\pid_alt.error_i_acumm_preregZ0Z_10 ));
    LocalMux I__5149 (
            .O(N__39088),
            .I(\pid_alt.error_i_acumm_preregZ0Z_10 ));
    LocalMux I__5148 (
            .O(N__39085),
            .I(\pid_alt.error_i_acumm_preregZ0Z_10 ));
    InMux I__5147 (
            .O(N__39078),
            .I(N__39075));
    LocalMux I__5146 (
            .O(N__39075),
            .I(N__39071));
    InMux I__5145 (
            .O(N__39074),
            .I(N__39068));
    Span4Mux_h I__5144 (
            .O(N__39071),
            .I(N__39065));
    LocalMux I__5143 (
            .O(N__39068),
            .I(\pid_alt.error_i_acummZ0Z_10 ));
    Odrv4 I__5142 (
            .O(N__39065),
            .I(\pid_alt.error_i_acummZ0Z_10 ));
    InMux I__5141 (
            .O(N__39060),
            .I(N__39056));
    CascadeMux I__5140 (
            .O(N__39059),
            .I(N__39053));
    LocalMux I__5139 (
            .O(N__39056),
            .I(N__39049));
    InMux I__5138 (
            .O(N__39053),
            .I(N__39046));
    CascadeMux I__5137 (
            .O(N__39052),
            .I(N__39043));
    Span4Mux_h I__5136 (
            .O(N__39049),
            .I(N__39038));
    LocalMux I__5135 (
            .O(N__39046),
            .I(N__39038));
    InMux I__5134 (
            .O(N__39043),
            .I(N__39035));
    Odrv4 I__5133 (
            .O(N__39038),
            .I(\pid_alt.error_i_acumm_preregZ0Z_11 ));
    LocalMux I__5132 (
            .O(N__39035),
            .I(\pid_alt.error_i_acumm_preregZ0Z_11 ));
    InMux I__5131 (
            .O(N__39030),
            .I(N__39027));
    LocalMux I__5130 (
            .O(N__39027),
            .I(\dron_frame_decoder_1.drone_altitude_6 ));
    InMux I__5129 (
            .O(N__39024),
            .I(N__39021));
    LocalMux I__5128 (
            .O(N__39021),
            .I(drone_altitude_i_6));
    InMux I__5127 (
            .O(N__39018),
            .I(N__39015));
    LocalMux I__5126 (
            .O(N__39015),
            .I(\dron_frame_decoder_1.drone_altitude_7 ));
    InMux I__5125 (
            .O(N__39012),
            .I(N__39009));
    LocalMux I__5124 (
            .O(N__39009),
            .I(drone_altitude_i_7));
    InMux I__5123 (
            .O(N__39006),
            .I(N__39003));
    LocalMux I__5122 (
            .O(N__39003),
            .I(drone_altitude_i_8));
    InMux I__5121 (
            .O(N__39000),
            .I(N__38997));
    LocalMux I__5120 (
            .O(N__38997),
            .I(drone_altitude_i_9));
    InMux I__5119 (
            .O(N__38994),
            .I(N__38991));
    LocalMux I__5118 (
            .O(N__38991),
            .I(N__38988));
    Span4Mux_v I__5117 (
            .O(N__38988),
            .I(N__38985));
    Span4Mux_s1_h I__5116 (
            .O(N__38985),
            .I(N__38982));
    Span4Mux_h I__5115 (
            .O(N__38982),
            .I(N__38979));
    Odrv4 I__5114 (
            .O(N__38979),
            .I(alt_kp_0));
    InMux I__5113 (
            .O(N__38976),
            .I(N__38973));
    LocalMux I__5112 (
            .O(N__38973),
            .I(N__38970));
    Span12Mux_s11_v I__5111 (
            .O(N__38970),
            .I(N__38967));
    Odrv12 I__5110 (
            .O(N__38967),
            .I(alt_kp_1));
    InMux I__5109 (
            .O(N__38964),
            .I(N__38961));
    LocalMux I__5108 (
            .O(N__38961),
            .I(N__38958));
    Span4Mux_v I__5107 (
            .O(N__38958),
            .I(N__38955));
    Span4Mux_h I__5106 (
            .O(N__38955),
            .I(N__38952));
    Odrv4 I__5105 (
            .O(N__38952),
            .I(alt_kp_2));
    InMux I__5104 (
            .O(N__38949),
            .I(N__38946));
    LocalMux I__5103 (
            .O(N__38946),
            .I(N__38943));
    Span4Mux_v I__5102 (
            .O(N__38943),
            .I(N__38940));
    Span4Mux_v I__5101 (
            .O(N__38940),
            .I(N__38937));
    Span4Mux_h I__5100 (
            .O(N__38937),
            .I(N__38934));
    Odrv4 I__5099 (
            .O(N__38934),
            .I(alt_kp_3));
    InMux I__5098 (
            .O(N__38931),
            .I(N__38928));
    LocalMux I__5097 (
            .O(N__38928),
            .I(N__38925));
    Span4Mux_v I__5096 (
            .O(N__38925),
            .I(N__38922));
    Span4Mux_h I__5095 (
            .O(N__38922),
            .I(N__38919));
    Odrv4 I__5094 (
            .O(N__38919),
            .I(alt_kp_5));
    InMux I__5093 (
            .O(N__38916),
            .I(N__38912));
    InMux I__5092 (
            .O(N__38915),
            .I(N__38908));
    LocalMux I__5091 (
            .O(N__38912),
            .I(N__38905));
    InMux I__5090 (
            .O(N__38911),
            .I(N__38902));
    LocalMux I__5089 (
            .O(N__38908),
            .I(N__38897));
    Span4Mux_v I__5088 (
            .O(N__38905),
            .I(N__38897));
    LocalMux I__5087 (
            .O(N__38902),
            .I(N__38894));
    Span4Mux_v I__5086 (
            .O(N__38897),
            .I(N__38891));
    Span12Mux_s5_h I__5085 (
            .O(N__38894),
            .I(N__38887));
    Span4Mux_h I__5084 (
            .O(N__38891),
            .I(N__38884));
    InMux I__5083 (
            .O(N__38890),
            .I(N__38881));
    Odrv12 I__5082 (
            .O(N__38887),
            .I(drone_altitude_0));
    Odrv4 I__5081 (
            .O(N__38884),
            .I(drone_altitude_0));
    LocalMux I__5080 (
            .O(N__38881),
            .I(drone_altitude_0));
    InMux I__5079 (
            .O(N__38874),
            .I(N__38871));
    LocalMux I__5078 (
            .O(N__38871),
            .I(drone_altitude_1));
    InMux I__5077 (
            .O(N__38868),
            .I(N__38865));
    LocalMux I__5076 (
            .O(N__38865),
            .I(\dron_frame_decoder_1.drone_altitude_4 ));
    InMux I__5075 (
            .O(N__38862),
            .I(N__38859));
    LocalMux I__5074 (
            .O(N__38859),
            .I(drone_altitude_i_4));
    InMux I__5073 (
            .O(N__38856),
            .I(N__38853));
    LocalMux I__5072 (
            .O(N__38853),
            .I(\dron_frame_decoder_1.drone_altitude_5 ));
    InMux I__5071 (
            .O(N__38850),
            .I(N__38847));
    LocalMux I__5070 (
            .O(N__38847),
            .I(drone_altitude_i_5));
    InMux I__5069 (
            .O(N__38844),
            .I(N__38841));
    LocalMux I__5068 (
            .O(N__38841),
            .I(N__38838));
    Odrv4 I__5067 (
            .O(N__38838),
            .I(\pid_alt.error_d_reg_prev_esr_RNI64JA4Z0Z_12 ));
    InMux I__5066 (
            .O(N__38835),
            .I(N__38832));
    LocalMux I__5065 (
            .O(N__38832),
            .I(\pid_alt.error_d_reg_prev_esr_RNIJGHMZ0Z_12 ));
    InMux I__5064 (
            .O(N__38829),
            .I(N__38822));
    InMux I__5063 (
            .O(N__38828),
            .I(N__38822));
    InMux I__5062 (
            .O(N__38827),
            .I(N__38819));
    LocalMux I__5061 (
            .O(N__38822),
            .I(N__38816));
    LocalMux I__5060 (
            .O(N__38819),
            .I(N__38813));
    Span4Mux_v I__5059 (
            .O(N__38816),
            .I(N__38810));
    Odrv4 I__5058 (
            .O(N__38813),
            .I(\pid_alt.error_i_acumm_esr_RNIJ6LMZ0Z_13 ));
    Odrv4 I__5057 (
            .O(N__38810),
            .I(\pid_alt.error_i_acumm_esr_RNIJ6LMZ0Z_13 ));
    CascadeMux I__5056 (
            .O(N__38805),
            .I(\pid_alt.error_d_reg_prev_esr_RNIJGHMZ0Z_12_cascade_ ));
    CascadeMux I__5055 (
            .O(N__38802),
            .I(N__38799));
    InMux I__5054 (
            .O(N__38799),
            .I(N__38795));
    InMux I__5053 (
            .O(N__38798),
            .I(N__38792));
    LocalMux I__5052 (
            .O(N__38795),
            .I(N__38789));
    LocalMux I__5051 (
            .O(N__38792),
            .I(\pid_alt.error_d_reg_prev_esr_RNISAO32Z0Z_12 ));
    Odrv4 I__5050 (
            .O(N__38789),
            .I(\pid_alt.error_d_reg_prev_esr_RNISAO32Z0Z_12 ));
    InMux I__5049 (
            .O(N__38784),
            .I(N__38780));
    InMux I__5048 (
            .O(N__38783),
            .I(N__38777));
    LocalMux I__5047 (
            .O(N__38780),
            .I(N__38774));
    LocalMux I__5046 (
            .O(N__38777),
            .I(N__38771));
    Span4Mux_v I__5045 (
            .O(N__38774),
            .I(N__38766));
    Span4Mux_h I__5044 (
            .O(N__38771),
            .I(N__38766));
    Span4Mux_v I__5043 (
            .O(N__38766),
            .I(N__38763));
    Odrv4 I__5042 (
            .O(N__38763),
            .I(\pid_alt.error_p_regZ0Z_13 ));
    InMux I__5041 (
            .O(N__38760),
            .I(N__38756));
    InMux I__5040 (
            .O(N__38759),
            .I(N__38753));
    LocalMux I__5039 (
            .O(N__38756),
            .I(N__38750));
    LocalMux I__5038 (
            .O(N__38753),
            .I(N__38747));
    Span4Mux_v I__5037 (
            .O(N__38750),
            .I(N__38742));
    Span4Mux_h I__5036 (
            .O(N__38747),
            .I(N__38742));
    Span4Mux_v I__5035 (
            .O(N__38742),
            .I(N__38739));
    Odrv4 I__5034 (
            .O(N__38739),
            .I(\pid_alt.error_d_reg_prevZ0Z_13 ));
    InMux I__5033 (
            .O(N__38736),
            .I(N__38733));
    LocalMux I__5032 (
            .O(N__38733),
            .I(N__38730));
    Span4Mux_v I__5031 (
            .O(N__38730),
            .I(N__38726));
    InMux I__5030 (
            .O(N__38729),
            .I(N__38723));
    Span4Mux_v I__5029 (
            .O(N__38726),
            .I(N__38720));
    LocalMux I__5028 (
            .O(N__38723),
            .I(N__38716));
    Sp12to4 I__5027 (
            .O(N__38720),
            .I(N__38713));
    InMux I__5026 (
            .O(N__38719),
            .I(N__38710));
    Span4Mux_v I__5025 (
            .O(N__38716),
            .I(N__38707));
    Span12Mux_s5_h I__5024 (
            .O(N__38713),
            .I(N__38702));
    LocalMux I__5023 (
            .O(N__38710),
            .I(N__38702));
    Span4Mux_v I__5022 (
            .O(N__38707),
            .I(N__38699));
    Span12Mux_v I__5021 (
            .O(N__38702),
            .I(N__38696));
    Odrv4 I__5020 (
            .O(N__38699),
            .I(\pid_alt.error_d_regZ0Z_13 ));
    Odrv12 I__5019 (
            .O(N__38696),
            .I(\pid_alt.error_d_regZ0Z_13 ));
    InMux I__5018 (
            .O(N__38691),
            .I(N__38685));
    InMux I__5017 (
            .O(N__38690),
            .I(N__38685));
    LocalMux I__5016 (
            .O(N__38685),
            .I(\pid_alt.error_d_reg_prev_esr_RNIMJHM_0Z0Z_13 ));
    CascadeMux I__5015 (
            .O(N__38682),
            .I(N__38678));
    CascadeMux I__5014 (
            .O(N__38681),
            .I(N__38675));
    InMux I__5013 (
            .O(N__38678),
            .I(N__38672));
    InMux I__5012 (
            .O(N__38675),
            .I(N__38669));
    LocalMux I__5011 (
            .O(N__38672),
            .I(N__38666));
    LocalMux I__5010 (
            .O(N__38669),
            .I(\pid_alt.error_d_reg_prev_esr_RNIAPQ62Z0Z_11 ));
    Odrv4 I__5009 (
            .O(N__38666),
            .I(\pid_alt.error_d_reg_prev_esr_RNIAPQ62Z0Z_11 ));
    InMux I__5008 (
            .O(N__38661),
            .I(N__38655));
    InMux I__5007 (
            .O(N__38660),
            .I(N__38655));
    LocalMux I__5006 (
            .O(N__38655),
            .I(\pid_alt.error_d_reg_prevZ0Z_12 ));
    InMux I__5005 (
            .O(N__38652),
            .I(N__38646));
    InMux I__5004 (
            .O(N__38651),
            .I(N__38646));
    LocalMux I__5003 (
            .O(N__38646),
            .I(N__38643));
    Span4Mux_v I__5002 (
            .O(N__38643),
            .I(N__38640));
    Span4Mux_h I__5001 (
            .O(N__38640),
            .I(N__38637));
    Odrv4 I__5000 (
            .O(N__38637),
            .I(\pid_alt.error_p_regZ0Z_12 ));
    InMux I__4999 (
            .O(N__38634),
            .I(N__38627));
    InMux I__4998 (
            .O(N__38633),
            .I(N__38627));
    InMux I__4997 (
            .O(N__38632),
            .I(N__38624));
    LocalMux I__4996 (
            .O(N__38627),
            .I(N__38619));
    LocalMux I__4995 (
            .O(N__38624),
            .I(N__38619));
    Span12Mux_v I__4994 (
            .O(N__38619),
            .I(N__38616));
    Odrv12 I__4993 (
            .O(N__38616),
            .I(\pid_alt.error_d_regZ0Z_12 ));
    InMux I__4992 (
            .O(N__38613),
            .I(N__38610));
    LocalMux I__4991 (
            .O(N__38610),
            .I(\pid_alt.error_d_reg_prev_esr_RNIJGHM_0Z0Z_12 ));
    InMux I__4990 (
            .O(N__38607),
            .I(N__38603));
    CascadeMux I__4989 (
            .O(N__38606),
            .I(N__38600));
    LocalMux I__4988 (
            .O(N__38603),
            .I(N__38597));
    InMux I__4987 (
            .O(N__38600),
            .I(N__38594));
    Span4Mux_h I__4986 (
            .O(N__38597),
            .I(N__38589));
    LocalMux I__4985 (
            .O(N__38594),
            .I(N__38589));
    Odrv4 I__4984 (
            .O(N__38589),
            .I(\pid_alt.error_d_reg_prev_esr_RNI1FP62Z0Z_10 ));
    InMux I__4983 (
            .O(N__38586),
            .I(N__38580));
    InMux I__4982 (
            .O(N__38585),
            .I(N__38580));
    LocalMux I__4981 (
            .O(N__38580),
            .I(N__38577));
    Odrv12 I__4980 (
            .O(N__38577),
            .I(\pid_alt.error_d_reg_prev_esr_RNIGDHMZ0Z_11 ));
    CascadeMux I__4979 (
            .O(N__38574),
            .I(\pid_alt.error_d_reg_prev_esr_RNIJGHM_0Z0Z_12_cascade_ ));
    InMux I__4978 (
            .O(N__38571),
            .I(N__38566));
    InMux I__4977 (
            .O(N__38570),
            .I(N__38561));
    InMux I__4976 (
            .O(N__38569),
            .I(N__38561));
    LocalMux I__4975 (
            .O(N__38566),
            .I(N__38558));
    LocalMux I__4974 (
            .O(N__38561),
            .I(N__38555));
    Span4Mux_v I__4973 (
            .O(N__38558),
            .I(N__38552));
    Span4Mux_v I__4972 (
            .O(N__38555),
            .I(N__38549));
    Odrv4 I__4971 (
            .O(N__38552),
            .I(\pid_alt.error_i_reg_esr_RNI7RNPZ0Z_12 ));
    Odrv4 I__4970 (
            .O(N__38549),
            .I(\pid_alt.error_i_reg_esr_RNI7RNPZ0Z_12 ));
    InMux I__4969 (
            .O(N__38544),
            .I(N__38541));
    LocalMux I__4968 (
            .O(N__38541),
            .I(N__38538));
    Odrv4 I__4967 (
            .O(N__38538),
            .I(\pid_alt.error_d_reg_prev_esr_RNIB8KD4Z0Z_11 ));
    InMux I__4966 (
            .O(N__38535),
            .I(N__38531));
    InMux I__4965 (
            .O(N__38534),
            .I(N__38528));
    LocalMux I__4964 (
            .O(N__38531),
            .I(N__38525));
    LocalMux I__4963 (
            .O(N__38528),
            .I(N__38522));
    Span4Mux_h I__4962 (
            .O(N__38525),
            .I(N__38519));
    Odrv4 I__4961 (
            .O(N__38522),
            .I(\Commands_frame_decoder.stateZ0Z_2 ));
    Odrv4 I__4960 (
            .O(N__38519),
            .I(\Commands_frame_decoder.stateZ0Z_2 ));
    CascadeMux I__4959 (
            .O(N__38514),
            .I(\Commands_frame_decoder.un1_sink_data_valid_2_0_cascade_ ));
    CascadeMux I__4958 (
            .O(N__38511),
            .I(N__38507));
    CascadeMux I__4957 (
            .O(N__38510),
            .I(N__38503));
    InMux I__4956 (
            .O(N__38507),
            .I(N__38497));
    InMux I__4955 (
            .O(N__38506),
            .I(N__38497));
    InMux I__4954 (
            .O(N__38503),
            .I(N__38492));
    InMux I__4953 (
            .O(N__38502),
            .I(N__38492));
    LocalMux I__4952 (
            .O(N__38497),
            .I(N__38486));
    LocalMux I__4951 (
            .O(N__38492),
            .I(N__38486));
    InMux I__4950 (
            .O(N__38491),
            .I(N__38483));
    Odrv4 I__4949 (
            .O(N__38486),
            .I(\Commands_frame_decoder.un1_sink_data_valid_2_0 ));
    LocalMux I__4948 (
            .O(N__38483),
            .I(\Commands_frame_decoder.un1_sink_data_valid_2_0 ));
    InMux I__4947 (
            .O(N__38478),
            .I(N__38472));
    InMux I__4946 (
            .O(N__38477),
            .I(N__38472));
    LocalMux I__4945 (
            .O(N__38472),
            .I(\Commands_frame_decoder.stateZ0Z_3 ));
    CascadeMux I__4944 (
            .O(N__38469),
            .I(N__38466));
    InMux I__4943 (
            .O(N__38466),
            .I(N__38454));
    InMux I__4942 (
            .O(N__38465),
            .I(N__38454));
    CascadeMux I__4941 (
            .O(N__38464),
            .I(N__38451));
    CascadeMux I__4940 (
            .O(N__38463),
            .I(N__38444));
    InMux I__4939 (
            .O(N__38462),
            .I(N__38430));
    InMux I__4938 (
            .O(N__38461),
            .I(N__38430));
    InMux I__4937 (
            .O(N__38460),
            .I(N__38430));
    InMux I__4936 (
            .O(N__38459),
            .I(N__38430));
    LocalMux I__4935 (
            .O(N__38454),
            .I(N__38427));
    InMux I__4934 (
            .O(N__38451),
            .I(N__38414));
    InMux I__4933 (
            .O(N__38450),
            .I(N__38414));
    InMux I__4932 (
            .O(N__38449),
            .I(N__38414));
    InMux I__4931 (
            .O(N__38448),
            .I(N__38414));
    InMux I__4930 (
            .O(N__38447),
            .I(N__38414));
    InMux I__4929 (
            .O(N__38444),
            .I(N__38414));
    InMux I__4928 (
            .O(N__38443),
            .I(N__38403));
    InMux I__4927 (
            .O(N__38442),
            .I(N__38403));
    InMux I__4926 (
            .O(N__38441),
            .I(N__38403));
    InMux I__4925 (
            .O(N__38440),
            .I(N__38403));
    InMux I__4924 (
            .O(N__38439),
            .I(N__38403));
    LocalMux I__4923 (
            .O(N__38430),
            .I(N__38395));
    Span4Mux_v I__4922 (
            .O(N__38427),
            .I(N__38388));
    LocalMux I__4921 (
            .O(N__38414),
            .I(N__38388));
    LocalMux I__4920 (
            .O(N__38403),
            .I(N__38388));
    InMux I__4919 (
            .O(N__38402),
            .I(N__38383));
    InMux I__4918 (
            .O(N__38401),
            .I(N__38383));
    InMux I__4917 (
            .O(N__38400),
            .I(N__38378));
    InMux I__4916 (
            .O(N__38399),
            .I(N__38378));
    InMux I__4915 (
            .O(N__38398),
            .I(N__38375));
    Span4Mux_v I__4914 (
            .O(N__38395),
            .I(N__38369));
    Span4Mux_v I__4913 (
            .O(N__38388),
            .I(N__38369));
    LocalMux I__4912 (
            .O(N__38383),
            .I(N__38362));
    LocalMux I__4911 (
            .O(N__38378),
            .I(N__38357));
    LocalMux I__4910 (
            .O(N__38375),
            .I(N__38357));
    InMux I__4909 (
            .O(N__38374),
            .I(N__38354));
    Span4Mux_s3_h I__4908 (
            .O(N__38369),
            .I(N__38351));
    InMux I__4907 (
            .O(N__38368),
            .I(N__38348));
    InMux I__4906 (
            .O(N__38367),
            .I(N__38341));
    InMux I__4905 (
            .O(N__38366),
            .I(N__38341));
    InMux I__4904 (
            .O(N__38365),
            .I(N__38341));
    Span4Mux_h I__4903 (
            .O(N__38362),
            .I(N__38338));
    Span4Mux_h I__4902 (
            .O(N__38357),
            .I(N__38335));
    LocalMux I__4901 (
            .O(N__38354),
            .I(uart_pc_data_rdy));
    Odrv4 I__4900 (
            .O(N__38351),
            .I(uart_pc_data_rdy));
    LocalMux I__4899 (
            .O(N__38348),
            .I(uart_pc_data_rdy));
    LocalMux I__4898 (
            .O(N__38341),
            .I(uart_pc_data_rdy));
    Odrv4 I__4897 (
            .O(N__38338),
            .I(uart_pc_data_rdy));
    Odrv4 I__4896 (
            .O(N__38335),
            .I(uart_pc_data_rdy));
    InMux I__4895 (
            .O(N__38322),
            .I(N__38319));
    LocalMux I__4894 (
            .O(N__38319),
            .I(\Commands_frame_decoder.source_CH2data_1_sqmuxa ));
    CascadeMux I__4893 (
            .O(N__38316),
            .I(\Commands_frame_decoder.source_CH2data_1_sqmuxa_cascade_ ));
    InMux I__4892 (
            .O(N__38313),
            .I(N__38310));
    LocalMux I__4891 (
            .O(N__38310),
            .I(N__38306));
    InMux I__4890 (
            .O(N__38309),
            .I(N__38303));
    Span4Mux_h I__4889 (
            .O(N__38306),
            .I(N__38300));
    LocalMux I__4888 (
            .O(N__38303),
            .I(\Commands_frame_decoder.stateZ0Z_4 ));
    Odrv4 I__4887 (
            .O(N__38300),
            .I(\Commands_frame_decoder.stateZ0Z_4 ));
    InMux I__4886 (
            .O(N__38295),
            .I(N__38292));
    LocalMux I__4885 (
            .O(N__38292),
            .I(N__38289));
    Span4Mux_h I__4884 (
            .O(N__38289),
            .I(N__38286));
    Span4Mux_h I__4883 (
            .O(N__38286),
            .I(N__38283));
    Odrv4 I__4882 (
            .O(N__38283),
            .I(\pid_front.O_0_20 ));
    InMux I__4881 (
            .O(N__38280),
            .I(N__38277));
    LocalMux I__4880 (
            .O(N__38277),
            .I(N__38274));
    Odrv12 I__4879 (
            .O(N__38274),
            .I(\pid_front.O_0_6 ));
    InMux I__4878 (
            .O(N__38271),
            .I(N__38268));
    LocalMux I__4877 (
            .O(N__38268),
            .I(N__38265));
    Span4Mux_h I__4876 (
            .O(N__38265),
            .I(N__38262));
    Span4Mux_h I__4875 (
            .O(N__38262),
            .I(N__38259));
    Odrv4 I__4874 (
            .O(N__38259),
            .I(\pid_front.O_0_12 ));
    InMux I__4873 (
            .O(N__38256),
            .I(N__38252));
    InMux I__4872 (
            .O(N__38255),
            .I(N__38249));
    LocalMux I__4871 (
            .O(N__38252),
            .I(\uart_pc.data_AuxZ0Z_7 ));
    LocalMux I__4870 (
            .O(N__38249),
            .I(\uart_pc.data_AuxZ0Z_7 ));
    CascadeMux I__4869 (
            .O(N__38244),
            .I(\uart_pc.N_145_cascade_ ));
    InMux I__4868 (
            .O(N__38241),
            .I(N__38238));
    LocalMux I__4867 (
            .O(N__38238),
            .I(\uart_pc.N_144_1 ));
    CascadeMux I__4866 (
            .O(N__38235),
            .I(\uart_pc.N_144_1_cascade_ ));
    InMux I__4865 (
            .O(N__38232),
            .I(N__38228));
    InMux I__4864 (
            .O(N__38231),
            .I(N__38225));
    LocalMux I__4863 (
            .O(N__38228),
            .I(N__38222));
    LocalMux I__4862 (
            .O(N__38225),
            .I(\Commands_frame_decoder.stateZ0Z_12 ));
    Odrv4 I__4861 (
            .O(N__38222),
            .I(\Commands_frame_decoder.stateZ0Z_12 ));
    CascadeMux I__4860 (
            .O(N__38217),
            .I(N__38214));
    InMux I__4859 (
            .O(N__38214),
            .I(N__38210));
    CascadeMux I__4858 (
            .O(N__38213),
            .I(N__38206));
    LocalMux I__4857 (
            .O(N__38210),
            .I(N__38203));
    InMux I__4856 (
            .O(N__38209),
            .I(N__38197));
    InMux I__4855 (
            .O(N__38206),
            .I(N__38197));
    Span4Mux_h I__4854 (
            .O(N__38203),
            .I(N__38194));
    InMux I__4853 (
            .O(N__38202),
            .I(N__38191));
    LocalMux I__4852 (
            .O(N__38197),
            .I(\Commands_frame_decoder.stateZ0Z_6 ));
    Odrv4 I__4851 (
            .O(N__38194),
            .I(\Commands_frame_decoder.stateZ0Z_6 ));
    LocalMux I__4850 (
            .O(N__38191),
            .I(\Commands_frame_decoder.stateZ0Z_6 ));
    InMux I__4849 (
            .O(N__38184),
            .I(N__38181));
    LocalMux I__4848 (
            .O(N__38181),
            .I(N__38178));
    Span4Mux_v I__4847 (
            .O(N__38178),
            .I(N__38175));
    Span4Mux_h I__4846 (
            .O(N__38175),
            .I(N__38171));
    InMux I__4845 (
            .O(N__38174),
            .I(N__38168));
    Span4Mux_v I__4844 (
            .O(N__38171),
            .I(N__38165));
    LocalMux I__4843 (
            .O(N__38168),
            .I(alt_kp_4));
    Odrv4 I__4842 (
            .O(N__38165),
            .I(alt_kp_4));
    InMux I__4841 (
            .O(N__38160),
            .I(N__38157));
    LocalMux I__4840 (
            .O(N__38157),
            .I(N__38154));
    Span4Mux_h I__4839 (
            .O(N__38154),
            .I(N__38148));
    InMux I__4838 (
            .O(N__38153),
            .I(N__38145));
    InMux I__4837 (
            .O(N__38152),
            .I(N__38140));
    InMux I__4836 (
            .O(N__38151),
            .I(N__38140));
    Odrv4 I__4835 (
            .O(N__38148),
            .I(\uart_pc.data_rdyc_1 ));
    LocalMux I__4834 (
            .O(N__38145),
            .I(\uart_pc.data_rdyc_1 ));
    LocalMux I__4833 (
            .O(N__38140),
            .I(\uart_pc.data_rdyc_1 ));
    InMux I__4832 (
            .O(N__38133),
            .I(N__38130));
    LocalMux I__4831 (
            .O(N__38130),
            .I(\uart_pc.data_Auxce_0_0_0 ));
    CascadeMux I__4830 (
            .O(N__38127),
            .I(N__38123));
    CascadeMux I__4829 (
            .O(N__38126),
            .I(N__38120));
    InMux I__4828 (
            .O(N__38123),
            .I(N__38117));
    InMux I__4827 (
            .O(N__38120),
            .I(N__38114));
    LocalMux I__4826 (
            .O(N__38117),
            .I(\uart_pc.data_AuxZ1Z_0 ));
    LocalMux I__4825 (
            .O(N__38114),
            .I(\uart_pc.data_AuxZ1Z_0 ));
    InMux I__4824 (
            .O(N__38109),
            .I(N__38106));
    LocalMux I__4823 (
            .O(N__38106),
            .I(\uart_pc.data_Auxce_0_1 ));
    CascadeMux I__4822 (
            .O(N__38103),
            .I(N__38099));
    InMux I__4821 (
            .O(N__38102),
            .I(N__38096));
    InMux I__4820 (
            .O(N__38099),
            .I(N__38093));
    LocalMux I__4819 (
            .O(N__38096),
            .I(N__38090));
    LocalMux I__4818 (
            .O(N__38093),
            .I(\uart_pc.data_AuxZ1Z_1 ));
    Odrv4 I__4817 (
            .O(N__38090),
            .I(\uart_pc.data_AuxZ1Z_1 ));
    InMux I__4816 (
            .O(N__38085),
            .I(N__38082));
    LocalMux I__4815 (
            .O(N__38082),
            .I(\uart_pc.data_Auxce_0_0_2 ));
    CascadeMux I__4814 (
            .O(N__38079),
            .I(N__38075));
    InMux I__4813 (
            .O(N__38078),
            .I(N__38072));
    InMux I__4812 (
            .O(N__38075),
            .I(N__38069));
    LocalMux I__4811 (
            .O(N__38072),
            .I(\uart_pc.data_AuxZ1Z_2 ));
    LocalMux I__4810 (
            .O(N__38069),
            .I(\uart_pc.data_AuxZ1Z_2 ));
    InMux I__4809 (
            .O(N__38064),
            .I(N__38061));
    LocalMux I__4808 (
            .O(N__38061),
            .I(\uart_pc.data_Auxce_0_3 ));
    CascadeMux I__4807 (
            .O(N__38058),
            .I(N__38055));
    InMux I__4806 (
            .O(N__38055),
            .I(N__38051));
    InMux I__4805 (
            .O(N__38054),
            .I(N__38048));
    LocalMux I__4804 (
            .O(N__38051),
            .I(\uart_pc.data_AuxZ0Z_3 ));
    LocalMux I__4803 (
            .O(N__38048),
            .I(\uart_pc.data_AuxZ0Z_3 ));
    InMux I__4802 (
            .O(N__38043),
            .I(N__38040));
    LocalMux I__4801 (
            .O(N__38040),
            .I(\uart_pc.data_Auxce_0_0_4 ));
    CascadeMux I__4800 (
            .O(N__38037),
            .I(N__38034));
    InMux I__4799 (
            .O(N__38034),
            .I(N__38031));
    LocalMux I__4798 (
            .O(N__38031),
            .I(N__38027));
    InMux I__4797 (
            .O(N__38030),
            .I(N__38024));
    Span4Mux_v I__4796 (
            .O(N__38027),
            .I(N__38021));
    LocalMux I__4795 (
            .O(N__38024),
            .I(\uart_pc.data_AuxZ0Z_4 ));
    Odrv4 I__4794 (
            .O(N__38021),
            .I(\uart_pc.data_AuxZ0Z_4 ));
    InMux I__4793 (
            .O(N__38016),
            .I(N__38013));
    LocalMux I__4792 (
            .O(N__38013),
            .I(N__38010));
    Odrv4 I__4791 (
            .O(N__38010),
            .I(\uart_pc.data_Auxce_0_5 ));
    InMux I__4790 (
            .O(N__38007),
            .I(N__38003));
    InMux I__4789 (
            .O(N__38006),
            .I(N__38000));
    LocalMux I__4788 (
            .O(N__38003),
            .I(\uart_pc.data_AuxZ0Z_5 ));
    LocalMux I__4787 (
            .O(N__38000),
            .I(\uart_pc.data_AuxZ0Z_5 ));
    CascadeMux I__4786 (
            .O(N__37995),
            .I(N__37992));
    InMux I__4785 (
            .O(N__37992),
            .I(N__37989));
    LocalMux I__4784 (
            .O(N__37989),
            .I(N__37986));
    Sp12to4 I__4783 (
            .O(N__37986),
            .I(N__37983));
    Odrv12 I__4782 (
            .O(N__37983),
            .I(\uart_pc.data_Auxce_0_6 ));
    InMux I__4781 (
            .O(N__37980),
            .I(N__37976));
    InMux I__4780 (
            .O(N__37979),
            .I(N__37973));
    LocalMux I__4779 (
            .O(N__37976),
            .I(\uart_pc.data_AuxZ0Z_6 ));
    LocalMux I__4778 (
            .O(N__37973),
            .I(\uart_pc.data_AuxZ0Z_6 ));
    InMux I__4777 (
            .O(N__37968),
            .I(N__37962));
    InMux I__4776 (
            .O(N__37967),
            .I(N__37962));
    LocalMux I__4775 (
            .O(N__37962),
            .I(N__37958));
    InMux I__4774 (
            .O(N__37961),
            .I(N__37955));
    Span4Mux_h I__4773 (
            .O(N__37958),
            .I(N__37952));
    LocalMux I__4772 (
            .O(N__37955),
            .I(N__37949));
    Span4Mux_v I__4771 (
            .O(N__37952),
            .I(N__37946));
    Span4Mux_v I__4770 (
            .O(N__37949),
            .I(N__37943));
    Odrv4 I__4769 (
            .O(N__37946),
            .I(\pid_alt.pid_preregZ0Z_6 ));
    Odrv4 I__4768 (
            .O(N__37943),
            .I(\pid_alt.pid_preregZ0Z_6 ));
    InMux I__4767 (
            .O(N__37938),
            .I(N__37932));
    InMux I__4766 (
            .O(N__37937),
            .I(N__37932));
    LocalMux I__4765 (
            .O(N__37932),
            .I(N__37928));
    InMux I__4764 (
            .O(N__37931),
            .I(N__37925));
    Span4Mux_h I__4763 (
            .O(N__37928),
            .I(N__37922));
    LocalMux I__4762 (
            .O(N__37925),
            .I(N__37919));
    Span4Mux_v I__4761 (
            .O(N__37922),
            .I(N__37916));
    Span4Mux_v I__4760 (
            .O(N__37919),
            .I(N__37913));
    Odrv4 I__4759 (
            .O(N__37916),
            .I(\pid_alt.pid_preregZ0Z_7 ));
    Odrv4 I__4758 (
            .O(N__37913),
            .I(\pid_alt.pid_preregZ0Z_7 ));
    InMux I__4757 (
            .O(N__37908),
            .I(N__37902));
    InMux I__4756 (
            .O(N__37907),
            .I(N__37902));
    LocalMux I__4755 (
            .O(N__37902),
            .I(N__37898));
    InMux I__4754 (
            .O(N__37901),
            .I(N__37895));
    Span4Mux_h I__4753 (
            .O(N__37898),
            .I(N__37892));
    LocalMux I__4752 (
            .O(N__37895),
            .I(N__37889));
    Span4Mux_v I__4751 (
            .O(N__37892),
            .I(N__37886));
    Span4Mux_v I__4750 (
            .O(N__37889),
            .I(N__37883));
    Odrv4 I__4749 (
            .O(N__37886),
            .I(\pid_alt.pid_preregZ0Z_8 ));
    Odrv4 I__4748 (
            .O(N__37883),
            .I(\pid_alt.pid_preregZ0Z_8 ));
    CascadeMux I__4747 (
            .O(N__37878),
            .I(N__37874));
    InMux I__4746 (
            .O(N__37877),
            .I(N__37868));
    InMux I__4745 (
            .O(N__37874),
            .I(N__37868));
    CascadeMux I__4744 (
            .O(N__37873),
            .I(N__37865));
    LocalMux I__4743 (
            .O(N__37868),
            .I(N__37862));
    InMux I__4742 (
            .O(N__37865),
            .I(N__37859));
    Span4Mux_v I__4741 (
            .O(N__37862),
            .I(N__37856));
    LocalMux I__4740 (
            .O(N__37859),
            .I(N__37853));
    Span4Mux_v I__4739 (
            .O(N__37856),
            .I(N__37850));
    Span4Mux_v I__4738 (
            .O(N__37853),
            .I(N__37847));
    Odrv4 I__4737 (
            .O(N__37850),
            .I(\pid_alt.pid_preregZ0Z_9 ));
    Odrv4 I__4736 (
            .O(N__37847),
            .I(\pid_alt.pid_preregZ0Z_9 ));
    CascadeMux I__4735 (
            .O(N__37842),
            .I(N__37836));
    InMux I__4734 (
            .O(N__37841),
            .I(N__37821));
    InMux I__4733 (
            .O(N__37840),
            .I(N__37821));
    InMux I__4732 (
            .O(N__37839),
            .I(N__37821));
    InMux I__4731 (
            .O(N__37836),
            .I(N__37821));
    InMux I__4730 (
            .O(N__37835),
            .I(N__37821));
    InMux I__4729 (
            .O(N__37834),
            .I(N__37821));
    LocalMux I__4728 (
            .O(N__37821),
            .I(\pid_alt.source_pid_9_0_tz_6 ));
    SRMux I__4727 (
            .O(N__37818),
            .I(N__37815));
    LocalMux I__4726 (
            .O(N__37815),
            .I(N__37809));
    SRMux I__4725 (
            .O(N__37814),
            .I(N__37806));
    SRMux I__4724 (
            .O(N__37813),
            .I(N__37803));
    SRMux I__4723 (
            .O(N__37812),
            .I(N__37800));
    Span4Mux_v I__4722 (
            .O(N__37809),
            .I(N__37795));
    LocalMux I__4721 (
            .O(N__37806),
            .I(N__37795));
    LocalMux I__4720 (
            .O(N__37803),
            .I(N__37790));
    LocalMux I__4719 (
            .O(N__37800),
            .I(N__37790));
    Odrv4 I__4718 (
            .O(N__37795),
            .I(\pid_alt.un1_reset_0_i ));
    Odrv4 I__4717 (
            .O(N__37790),
            .I(\pid_alt.un1_reset_0_i ));
    InMux I__4716 (
            .O(N__37785),
            .I(\uart_drone.un4_timer_Count_1_cry_3 ));
    InMux I__4715 (
            .O(N__37782),
            .I(N__37779));
    LocalMux I__4714 (
            .O(N__37779),
            .I(\uart_drone.timer_Count_RNO_0_0_4 ));
    InMux I__4713 (
            .O(N__37776),
            .I(N__37771));
    InMux I__4712 (
            .O(N__37775),
            .I(N__37767));
    InMux I__4711 (
            .O(N__37774),
            .I(N__37764));
    LocalMux I__4710 (
            .O(N__37771),
            .I(N__37761));
    CascadeMux I__4709 (
            .O(N__37770),
            .I(N__37756));
    LocalMux I__4708 (
            .O(N__37767),
            .I(N__37753));
    LocalMux I__4707 (
            .O(N__37764),
            .I(N__37750));
    Span4Mux_h I__4706 (
            .O(N__37761),
            .I(N__37747));
    InMux I__4705 (
            .O(N__37760),
            .I(N__37744));
    InMux I__4704 (
            .O(N__37759),
            .I(N__37741));
    InMux I__4703 (
            .O(N__37756),
            .I(N__37738));
    Span4Mux_v I__4702 (
            .O(N__37753),
            .I(N__37725));
    Span4Mux_h I__4701 (
            .O(N__37750),
            .I(N__37725));
    Span4Mux_h I__4700 (
            .O(N__37747),
            .I(N__37725));
    LocalMux I__4699 (
            .O(N__37744),
            .I(N__37725));
    LocalMux I__4698 (
            .O(N__37741),
            .I(N__37725));
    LocalMux I__4697 (
            .O(N__37738),
            .I(N__37725));
    Span4Mux_v I__4696 (
            .O(N__37725),
            .I(N__37722));
    Odrv4 I__4695 (
            .O(N__37722),
            .I(\pid_alt.pid_preregZ0Z_13 ));
    InMux I__4694 (
            .O(N__37719),
            .I(N__37714));
    InMux I__4693 (
            .O(N__37718),
            .I(N__37703));
    InMux I__4692 (
            .O(N__37717),
            .I(N__37703));
    LocalMux I__4691 (
            .O(N__37714),
            .I(N__37700));
    InMux I__4690 (
            .O(N__37713),
            .I(N__37695));
    InMux I__4689 (
            .O(N__37712),
            .I(N__37695));
    InMux I__4688 (
            .O(N__37711),
            .I(N__37684));
    InMux I__4687 (
            .O(N__37710),
            .I(N__37684));
    InMux I__4686 (
            .O(N__37709),
            .I(N__37684));
    InMux I__4685 (
            .O(N__37708),
            .I(N__37684));
    LocalMux I__4684 (
            .O(N__37703),
            .I(N__37681));
    Span4Mux_v I__4683 (
            .O(N__37700),
            .I(N__37678));
    LocalMux I__4682 (
            .O(N__37695),
            .I(N__37675));
    InMux I__4681 (
            .O(N__37694),
            .I(N__37670));
    InMux I__4680 (
            .O(N__37693),
            .I(N__37670));
    LocalMux I__4679 (
            .O(N__37684),
            .I(N__37667));
    Span4Mux_v I__4678 (
            .O(N__37681),
            .I(N__37664));
    Span4Mux_v I__4677 (
            .O(N__37678),
            .I(N__37661));
    Span4Mux_h I__4676 (
            .O(N__37675),
            .I(N__37658));
    LocalMux I__4675 (
            .O(N__37670),
            .I(\pid_alt.N_539 ));
    Odrv4 I__4674 (
            .O(N__37667),
            .I(\pid_alt.N_539 ));
    Odrv4 I__4673 (
            .O(N__37664),
            .I(\pid_alt.N_539 ));
    Odrv4 I__4672 (
            .O(N__37661),
            .I(\pid_alt.N_539 ));
    Odrv4 I__4671 (
            .O(N__37658),
            .I(\pid_alt.N_539 ));
    CascadeMux I__4670 (
            .O(N__37647),
            .I(N__37643));
    CascadeMux I__4669 (
            .O(N__37646),
            .I(N__37639));
    InMux I__4668 (
            .O(N__37643),
            .I(N__37635));
    CascadeMux I__4667 (
            .O(N__37642),
            .I(N__37632));
    InMux I__4666 (
            .O(N__37639),
            .I(N__37625));
    InMux I__4665 (
            .O(N__37638),
            .I(N__37625));
    LocalMux I__4664 (
            .O(N__37635),
            .I(N__37620));
    InMux I__4663 (
            .O(N__37632),
            .I(N__37613));
    InMux I__4662 (
            .O(N__37631),
            .I(N__37613));
    InMux I__4661 (
            .O(N__37630),
            .I(N__37610));
    LocalMux I__4660 (
            .O(N__37625),
            .I(N__37607));
    InMux I__4659 (
            .O(N__37624),
            .I(N__37604));
    InMux I__4658 (
            .O(N__37623),
            .I(N__37601));
    Span4Mux_v I__4657 (
            .O(N__37620),
            .I(N__37598));
    InMux I__4656 (
            .O(N__37619),
            .I(N__37593));
    InMux I__4655 (
            .O(N__37618),
            .I(N__37593));
    LocalMux I__4654 (
            .O(N__37613),
            .I(N__37590));
    LocalMux I__4653 (
            .O(N__37610),
            .I(N__37587));
    Span4Mux_v I__4652 (
            .O(N__37607),
            .I(N__37584));
    LocalMux I__4651 (
            .O(N__37604),
            .I(N__37579));
    LocalMux I__4650 (
            .O(N__37601),
            .I(N__37579));
    Span4Mux_v I__4649 (
            .O(N__37598),
            .I(N__37576));
    LocalMux I__4648 (
            .O(N__37593),
            .I(N__37569));
    Span4Mux_v I__4647 (
            .O(N__37590),
            .I(N__37569));
    Span4Mux_h I__4646 (
            .O(N__37587),
            .I(N__37569));
    Span4Mux_v I__4645 (
            .O(N__37584),
            .I(N__37566));
    Span4Mux_h I__4644 (
            .O(N__37579),
            .I(N__37563));
    Span4Mux_v I__4643 (
            .O(N__37576),
            .I(N__37560));
    Span4Mux_v I__4642 (
            .O(N__37569),
            .I(N__37557));
    Odrv4 I__4641 (
            .O(N__37566),
            .I(\pid_alt.pid_preregZ0Z_24 ));
    Odrv4 I__4640 (
            .O(N__37563),
            .I(\pid_alt.pid_preregZ0Z_24 ));
    Odrv4 I__4639 (
            .O(N__37560),
            .I(\pid_alt.pid_preregZ0Z_24 ));
    Odrv4 I__4638 (
            .O(N__37557),
            .I(\pid_alt.pid_preregZ0Z_24 ));
    InMux I__4637 (
            .O(N__37548),
            .I(N__37543));
    InMux I__4636 (
            .O(N__37547),
            .I(N__37540));
    InMux I__4635 (
            .O(N__37546),
            .I(N__37537));
    LocalMux I__4634 (
            .O(N__37543),
            .I(N__37531));
    LocalMux I__4633 (
            .O(N__37540),
            .I(N__37531));
    LocalMux I__4632 (
            .O(N__37537),
            .I(N__37528));
    InMux I__4631 (
            .O(N__37536),
            .I(N__37525));
    Span12Mux_h I__4630 (
            .O(N__37531),
            .I(N__37522));
    Span4Mux_v I__4629 (
            .O(N__37528),
            .I(N__37517));
    LocalMux I__4628 (
            .O(N__37525),
            .I(N__37517));
    Odrv12 I__4627 (
            .O(N__37522),
            .I(\pid_alt.pid_preregZ0Z_12 ));
    Odrv4 I__4626 (
            .O(N__37517),
            .I(\pid_alt.pid_preregZ0Z_12 ));
    CascadeMux I__4625 (
            .O(N__37512),
            .I(\uart_drone.timer_Count_RNO_0_0_1_cascade_ ));
    InMux I__4624 (
            .O(N__37509),
            .I(N__37503));
    InMux I__4623 (
            .O(N__37508),
            .I(N__37503));
    LocalMux I__4622 (
            .O(N__37503),
            .I(\uart_drone.timer_CountZ1Z_1 ));
    InMux I__4621 (
            .O(N__37500),
            .I(N__37494));
    InMux I__4620 (
            .O(N__37499),
            .I(N__37494));
    LocalMux I__4619 (
            .O(N__37494),
            .I(N__37490));
    InMux I__4618 (
            .O(N__37493),
            .I(N__37487));
    Span4Mux_v I__4617 (
            .O(N__37490),
            .I(N__37484));
    LocalMux I__4616 (
            .O(N__37487),
            .I(N__37481));
    Span4Mux_v I__4615 (
            .O(N__37484),
            .I(N__37478));
    Span4Mux_v I__4614 (
            .O(N__37481),
            .I(N__37475));
    Odrv4 I__4613 (
            .O(N__37478),
            .I(\pid_alt.pid_preregZ0Z_10 ));
    Odrv4 I__4612 (
            .O(N__37475),
            .I(\pid_alt.pid_preregZ0Z_10 ));
    CascadeMux I__4611 (
            .O(N__37470),
            .I(\pid_alt.source_pid_1_sqmuxa_0_a2_1_4_cascade_ ));
    InMux I__4610 (
            .O(N__37467),
            .I(N__37464));
    LocalMux I__4609 (
            .O(N__37464),
            .I(N__37461));
    Odrv4 I__4608 (
            .O(N__37461),
            .I(\pid_alt.source_pid_1_sqmuxa_0_a2_1_5 ));
    InMux I__4607 (
            .O(N__37458),
            .I(N__37453));
    InMux I__4606 (
            .O(N__37457),
            .I(N__37448));
    InMux I__4605 (
            .O(N__37456),
            .I(N__37448));
    LocalMux I__4604 (
            .O(N__37453),
            .I(N__37443));
    LocalMux I__4603 (
            .O(N__37448),
            .I(N__37443));
    Span4Mux_h I__4602 (
            .O(N__37443),
            .I(N__37440));
    Span4Mux_v I__4601 (
            .O(N__37440),
            .I(N__37437));
    Odrv4 I__4600 (
            .O(N__37437),
            .I(\pid_alt.pid_preregZ0Z_11 ));
    InMux I__4599 (
            .O(N__37434),
            .I(N__37431));
    LocalMux I__4598 (
            .O(N__37431),
            .I(\uart_drone_sync.aux_1__0__0_0 ));
    InMux I__4597 (
            .O(N__37428),
            .I(N__37425));
    LocalMux I__4596 (
            .O(N__37425),
            .I(\uart_drone_sync.aux_2__0__0_0 ));
    InMux I__4595 (
            .O(N__37422),
            .I(N__37419));
    LocalMux I__4594 (
            .O(N__37419),
            .I(\uart_drone_sync.aux_3__0__0_0 ));
    InMux I__4593 (
            .O(N__37416),
            .I(N__37413));
    LocalMux I__4592 (
            .O(N__37413),
            .I(\uart_drone.timer_Count_RNO_0_0_2 ));
    InMux I__4591 (
            .O(N__37410),
            .I(\uart_drone.un4_timer_Count_1_cry_1 ));
    InMux I__4590 (
            .O(N__37407),
            .I(\uart_drone.un4_timer_Count_1_cry_2 ));
    InMux I__4589 (
            .O(N__37404),
            .I(N__37401));
    LocalMux I__4588 (
            .O(N__37401),
            .I(\pid_alt.m35_e_3 ));
    InMux I__4587 (
            .O(N__37398),
            .I(N__37395));
    LocalMux I__4586 (
            .O(N__37395),
            .I(N__37392));
    Odrv4 I__4585 (
            .O(N__37392),
            .I(\pid_alt.m35_e_2 ));
    CascadeMux I__4584 (
            .O(N__37389),
            .I(\pid_alt.N_9_0_cascade_ ));
    InMux I__4583 (
            .O(N__37386),
            .I(N__37383));
    LocalMux I__4582 (
            .O(N__37383),
            .I(N__37379));
    InMux I__4581 (
            .O(N__37382),
            .I(N__37376));
    Odrv4 I__4580 (
            .O(N__37379),
            .I(\pid_alt.error_i_acumm_preregZ0Z_1 ));
    LocalMux I__4579 (
            .O(N__37376),
            .I(\pid_alt.error_i_acumm_preregZ0Z_1 ));
    CascadeMux I__4578 (
            .O(N__37371),
            .I(\pid_alt.N_62_mux_cascade_ ));
    InMux I__4577 (
            .O(N__37368),
            .I(N__37365));
    LocalMux I__4576 (
            .O(N__37365),
            .I(N__37362));
    Span4Mux_h I__4575 (
            .O(N__37362),
            .I(N__37359));
    Odrv4 I__4574 (
            .O(N__37359),
            .I(\pid_alt.error_i_acummZ0Z_1 ));
    InMux I__4573 (
            .O(N__37356),
            .I(N__37353));
    LocalMux I__4572 (
            .O(N__37353),
            .I(N__37349));
    InMux I__4571 (
            .O(N__37352),
            .I(N__37346));
    Odrv4 I__4570 (
            .O(N__37349),
            .I(\pid_alt.error_i_acumm_preregZ0Z_2 ));
    LocalMux I__4569 (
            .O(N__37346),
            .I(\pid_alt.error_i_acumm_preregZ0Z_2 ));
    InMux I__4568 (
            .O(N__37341),
            .I(N__37338));
    LocalMux I__4567 (
            .O(N__37338),
            .I(N__37335));
    Span4Mux_h I__4566 (
            .O(N__37335),
            .I(N__37332));
    Odrv4 I__4565 (
            .O(N__37332),
            .I(\pid_alt.error_i_acummZ0Z_2 ));
    CascadeMux I__4564 (
            .O(N__37329),
            .I(\pid_alt.N_159_cascade_ ));
    InMux I__4563 (
            .O(N__37326),
            .I(N__37323));
    LocalMux I__4562 (
            .O(N__37323),
            .I(N__37319));
    InMux I__4561 (
            .O(N__37322),
            .I(N__37316));
    Odrv4 I__4560 (
            .O(N__37319),
            .I(\pid_alt.error_i_acumm_preregZ0Z_0 ));
    LocalMux I__4559 (
            .O(N__37316),
            .I(\pid_alt.error_i_acumm_preregZ0Z_0 ));
    InMux I__4558 (
            .O(N__37311),
            .I(N__37307));
    InMux I__4557 (
            .O(N__37310),
            .I(N__37304));
    LocalMux I__4556 (
            .O(N__37307),
            .I(N__37301));
    LocalMux I__4555 (
            .O(N__37304),
            .I(N__37296));
    Span4Mux_h I__4554 (
            .O(N__37301),
            .I(N__37296));
    Odrv4 I__4553 (
            .O(N__37296),
            .I(\pid_alt.error_i_acummZ0Z_0 ));
    InMux I__4552 (
            .O(N__37293),
            .I(N__37290));
    LocalMux I__4551 (
            .O(N__37290),
            .I(N__37287));
    Span12Mux_v I__4550 (
            .O(N__37287),
            .I(N__37284));
    Odrv12 I__4549 (
            .O(N__37284),
            .I(\pid_alt.error_i_acummZ0Z_4 ));
    InMux I__4548 (
            .O(N__37281),
            .I(N__37277));
    InMux I__4547 (
            .O(N__37280),
            .I(N__37274));
    LocalMux I__4546 (
            .O(N__37277),
            .I(N__37269));
    LocalMux I__4545 (
            .O(N__37274),
            .I(N__37269));
    Odrv4 I__4544 (
            .O(N__37269),
            .I(\pid_alt.error_i_acumm_preregZ0Z_3 ));
    CascadeMux I__4543 (
            .O(N__37266),
            .I(N__37262));
    CascadeMux I__4542 (
            .O(N__37265),
            .I(N__37259));
    InMux I__4541 (
            .O(N__37262),
            .I(N__37251));
    InMux I__4540 (
            .O(N__37259),
            .I(N__37251));
    InMux I__4539 (
            .O(N__37258),
            .I(N__37251));
    LocalMux I__4538 (
            .O(N__37251),
            .I(\pid_alt.N_159 ));
    CascadeMux I__4537 (
            .O(N__37248),
            .I(N__37244));
    InMux I__4536 (
            .O(N__37247),
            .I(N__37237));
    InMux I__4535 (
            .O(N__37244),
            .I(N__37226));
    InMux I__4534 (
            .O(N__37243),
            .I(N__37226));
    InMux I__4533 (
            .O(N__37242),
            .I(N__37226));
    InMux I__4532 (
            .O(N__37241),
            .I(N__37226));
    InMux I__4531 (
            .O(N__37240),
            .I(N__37226));
    LocalMux I__4530 (
            .O(N__37237),
            .I(N__37223));
    LocalMux I__4529 (
            .O(N__37226),
            .I(\pid_alt.error_i_acumm7lto4 ));
    Odrv12 I__4528 (
            .O(N__37223),
            .I(\pid_alt.error_i_acumm7lto4 ));
    InMux I__4527 (
            .O(N__37218),
            .I(N__37215));
    LocalMux I__4526 (
            .O(N__37215),
            .I(N__37212));
    Span4Mux_s3_h I__4525 (
            .O(N__37212),
            .I(N__37209));
    Span4Mux_v I__4524 (
            .O(N__37209),
            .I(N__37206));
    Odrv4 I__4523 (
            .O(N__37206),
            .I(\pid_alt.error_i_acummZ0Z_3 ));
    InMux I__4522 (
            .O(N__37203),
            .I(N__37198));
    InMux I__4521 (
            .O(N__37202),
            .I(N__37193));
    InMux I__4520 (
            .O(N__37201),
            .I(N__37193));
    LocalMux I__4519 (
            .O(N__37198),
            .I(N__37190));
    LocalMux I__4518 (
            .O(N__37193),
            .I(N__37187));
    Span4Mux_h I__4517 (
            .O(N__37190),
            .I(N__37184));
    Span4Mux_v I__4516 (
            .O(N__37187),
            .I(N__37181));
    Odrv4 I__4515 (
            .O(N__37184),
            .I(\pid_alt.error_i_reg_esr_RNIT8KA1Z0Z_5 ));
    Odrv4 I__4514 (
            .O(N__37181),
            .I(\pid_alt.error_i_reg_esr_RNIT8KA1Z0Z_5 ));
    InMux I__4513 (
            .O(N__37176),
            .I(N__37173));
    LocalMux I__4512 (
            .O(N__37173),
            .I(N__37168));
    InMux I__4511 (
            .O(N__37172),
            .I(N__37163));
    InMux I__4510 (
            .O(N__37171),
            .I(N__37163));
    Span4Mux_h I__4509 (
            .O(N__37168),
            .I(N__37160));
    LocalMux I__4508 (
            .O(N__37163),
            .I(N__37157));
    Odrv4 I__4507 (
            .O(N__37160),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_7_c_RNI6LNQ ));
    Odrv4 I__4506 (
            .O(N__37157),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_7_c_RNI6LNQ ));
    InMux I__4505 (
            .O(N__37152),
            .I(N__37149));
    LocalMux I__4504 (
            .O(N__37149),
            .I(N__37146));
    Span4Mux_v I__4503 (
            .O(N__37146),
            .I(N__37141));
    InMux I__4502 (
            .O(N__37145),
            .I(N__37136));
    InMux I__4501 (
            .O(N__37144),
            .I(N__37136));
    Odrv4 I__4500 (
            .O(N__37141),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_9_c_RNIQN3F ));
    LocalMux I__4499 (
            .O(N__37136),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_9_c_RNIQN3F ));
    CascadeMux I__4498 (
            .O(N__37131),
            .I(\pid_alt.m21_e_2_cascade_ ));
    InMux I__4497 (
            .O(N__37128),
            .I(N__37125));
    LocalMux I__4496 (
            .O(N__37125),
            .I(N__37122));
    Span4Mux_h I__4495 (
            .O(N__37122),
            .I(N__37119));
    Odrv4 I__4494 (
            .O(N__37119),
            .I(\pid_alt.m21_e_8 ));
    InMux I__4493 (
            .O(N__37116),
            .I(N__37113));
    LocalMux I__4492 (
            .O(N__37113),
            .I(\pid_alt.m21_e_9 ));
    CascadeMux I__4491 (
            .O(N__37110),
            .I(\pid_alt.m21_e_10_cascade_ ));
    CascadeMux I__4490 (
            .O(N__37107),
            .I(\pid_alt.N_111_cascade_ ));
    InMux I__4489 (
            .O(N__37104),
            .I(N__37101));
    LocalMux I__4488 (
            .O(N__37101),
            .I(N__37098));
    Span4Mux_s1_h I__4487 (
            .O(N__37098),
            .I(N__37093));
    InMux I__4486 (
            .O(N__37097),
            .I(N__37090));
    InMux I__4485 (
            .O(N__37096),
            .I(N__37087));
    Span4Mux_v I__4484 (
            .O(N__37093),
            .I(N__37082));
    LocalMux I__4483 (
            .O(N__37090),
            .I(N__37082));
    LocalMux I__4482 (
            .O(N__37087),
            .I(N__37079));
    Span4Mux_v I__4481 (
            .O(N__37082),
            .I(N__37076));
    Span4Mux_v I__4480 (
            .O(N__37079),
            .I(N__37073));
    Span4Mux_v I__4479 (
            .O(N__37076),
            .I(N__37068));
    Span4Mux_v I__4478 (
            .O(N__37073),
            .I(N__37068));
    Odrv4 I__4477 (
            .O(N__37068),
            .I(\pid_alt.error_11 ));
    InMux I__4476 (
            .O(N__37065),
            .I(\pid_alt.error_cry_10 ));
    InMux I__4475 (
            .O(N__37062),
            .I(N__37059));
    LocalMux I__4474 (
            .O(N__37059),
            .I(N__37054));
    InMux I__4473 (
            .O(N__37058),
            .I(N__37051));
    InMux I__4472 (
            .O(N__37057),
            .I(N__37048));
    Span4Mux_h I__4471 (
            .O(N__37054),
            .I(N__37045));
    LocalMux I__4470 (
            .O(N__37051),
            .I(N__37042));
    LocalMux I__4469 (
            .O(N__37048),
            .I(N__37039));
    Span4Mux_v I__4468 (
            .O(N__37045),
            .I(N__37036));
    Span4Mux_v I__4467 (
            .O(N__37042),
            .I(N__37033));
    Span4Mux_v I__4466 (
            .O(N__37039),
            .I(N__37030));
    Span4Mux_v I__4465 (
            .O(N__37036),
            .I(N__37025));
    Span4Mux_h I__4464 (
            .O(N__37033),
            .I(N__37025));
    Span4Mux_h I__4463 (
            .O(N__37030),
            .I(N__37022));
    Odrv4 I__4462 (
            .O(N__37025),
            .I(\pid_alt.error_12 ));
    Odrv4 I__4461 (
            .O(N__37022),
            .I(\pid_alt.error_12 ));
    InMux I__4460 (
            .O(N__37017),
            .I(\pid_alt.error_cry_11 ));
    InMux I__4459 (
            .O(N__37014),
            .I(N__37011));
    LocalMux I__4458 (
            .O(N__37011),
            .I(N__37006));
    InMux I__4457 (
            .O(N__37010),
            .I(N__37003));
    InMux I__4456 (
            .O(N__37009),
            .I(N__37000));
    Span4Mux_h I__4455 (
            .O(N__37006),
            .I(N__36997));
    LocalMux I__4454 (
            .O(N__37003),
            .I(N__36994));
    LocalMux I__4453 (
            .O(N__37000),
            .I(N__36991));
    Span4Mux_v I__4452 (
            .O(N__36997),
            .I(N__36988));
    Span4Mux_v I__4451 (
            .O(N__36994),
            .I(N__36985));
    Span4Mux_v I__4450 (
            .O(N__36991),
            .I(N__36982));
    Span4Mux_v I__4449 (
            .O(N__36988),
            .I(N__36977));
    Span4Mux_h I__4448 (
            .O(N__36985),
            .I(N__36977));
    Span4Mux_h I__4447 (
            .O(N__36982),
            .I(N__36974));
    Odrv4 I__4446 (
            .O(N__36977),
            .I(\pid_alt.error_13 ));
    Odrv4 I__4445 (
            .O(N__36974),
            .I(\pid_alt.error_13 ));
    InMux I__4444 (
            .O(N__36969),
            .I(\pid_alt.error_cry_12 ));
    InMux I__4443 (
            .O(N__36966),
            .I(N__36963));
    LocalMux I__4442 (
            .O(N__36963),
            .I(N__36960));
    Span4Mux_v I__4441 (
            .O(N__36960),
            .I(N__36956));
    InMux I__4440 (
            .O(N__36959),
            .I(N__36953));
    Span4Mux_v I__4439 (
            .O(N__36956),
            .I(N__36947));
    LocalMux I__4438 (
            .O(N__36953),
            .I(N__36947));
    InMux I__4437 (
            .O(N__36952),
            .I(N__36944));
    Span4Mux_h I__4436 (
            .O(N__36947),
            .I(N__36941));
    LocalMux I__4435 (
            .O(N__36944),
            .I(N__36938));
    Span4Mux_v I__4434 (
            .O(N__36941),
            .I(N__36935));
    Span12Mux_s4_h I__4433 (
            .O(N__36938),
            .I(N__36932));
    Odrv4 I__4432 (
            .O(N__36935),
            .I(\pid_alt.error_14 ));
    Odrv12 I__4431 (
            .O(N__36932),
            .I(\pid_alt.error_14 ));
    InMux I__4430 (
            .O(N__36927),
            .I(\pid_alt.error_cry_13 ));
    InMux I__4429 (
            .O(N__36924),
            .I(\pid_alt.error_cry_14 ));
    InMux I__4428 (
            .O(N__36921),
            .I(N__36918));
    LocalMux I__4427 (
            .O(N__36918),
            .I(N__36915));
    Span4Mux_v I__4426 (
            .O(N__36915),
            .I(N__36910));
    InMux I__4425 (
            .O(N__36914),
            .I(N__36907));
    InMux I__4424 (
            .O(N__36913),
            .I(N__36904));
    Span4Mux_v I__4423 (
            .O(N__36910),
            .I(N__36899));
    LocalMux I__4422 (
            .O(N__36907),
            .I(N__36899));
    LocalMux I__4421 (
            .O(N__36904),
            .I(N__36896));
    Span4Mux_h I__4420 (
            .O(N__36899),
            .I(N__36893));
    Span4Mux_v I__4419 (
            .O(N__36896),
            .I(N__36890));
    Span4Mux_v I__4418 (
            .O(N__36893),
            .I(N__36887));
    Span4Mux_h I__4417 (
            .O(N__36890),
            .I(N__36884));
    Odrv4 I__4416 (
            .O(N__36887),
            .I(\pid_alt.error_15 ));
    Odrv4 I__4415 (
            .O(N__36884),
            .I(\pid_alt.error_15 ));
    InMux I__4414 (
            .O(N__36879),
            .I(N__36876));
    LocalMux I__4413 (
            .O(N__36876),
            .I(\pid_alt.m21_e_0 ));
    InMux I__4412 (
            .O(N__36873),
            .I(N__36868));
    InMux I__4411 (
            .O(N__36872),
            .I(N__36865));
    InMux I__4410 (
            .O(N__36871),
            .I(N__36862));
    LocalMux I__4409 (
            .O(N__36868),
            .I(N__36859));
    LocalMux I__4408 (
            .O(N__36865),
            .I(N__36856));
    LocalMux I__4407 (
            .O(N__36862),
            .I(N__36853));
    Span4Mux_h I__4406 (
            .O(N__36859),
            .I(N__36850));
    Span4Mux_h I__4405 (
            .O(N__36856),
            .I(N__36847));
    Odrv12 I__4404 (
            .O(N__36853),
            .I(\pid_alt.error_i_acumm_esr_RNIQMD91Z0Z_1 ));
    Odrv4 I__4403 (
            .O(N__36850),
            .I(\pid_alt.error_i_acumm_esr_RNIQMD91Z0Z_1 ));
    Odrv4 I__4402 (
            .O(N__36847),
            .I(\pid_alt.error_i_acumm_esr_RNIQMD91Z0Z_1 ));
    InMux I__4401 (
            .O(N__36840),
            .I(N__36836));
    CascadeMux I__4400 (
            .O(N__36839),
            .I(N__36833));
    LocalMux I__4399 (
            .O(N__36836),
            .I(N__36830));
    InMux I__4398 (
            .O(N__36833),
            .I(N__36827));
    Span4Mux_v I__4397 (
            .O(N__36830),
            .I(N__36824));
    LocalMux I__4396 (
            .O(N__36827),
            .I(N__36821));
    Span4Mux_v I__4395 (
            .O(N__36824),
            .I(N__36818));
    Span4Mux_v I__4394 (
            .O(N__36821),
            .I(N__36815));
    Odrv4 I__4393 (
            .O(N__36818),
            .I(\pid_alt.error_i_regZ0Z_0 ));
    Odrv4 I__4392 (
            .O(N__36815),
            .I(\pid_alt.error_i_regZ0Z_0 ));
    InMux I__4391 (
            .O(N__36810),
            .I(\pid_alt.error_cry_1 ));
    InMux I__4390 (
            .O(N__36807),
            .I(N__36804));
    LocalMux I__4389 (
            .O(N__36804),
            .I(N__36799));
    InMux I__4388 (
            .O(N__36803),
            .I(N__36796));
    InMux I__4387 (
            .O(N__36802),
            .I(N__36793));
    Span4Mux_h I__4386 (
            .O(N__36799),
            .I(N__36790));
    LocalMux I__4385 (
            .O(N__36796),
            .I(N__36787));
    LocalMux I__4384 (
            .O(N__36793),
            .I(N__36784));
    Span4Mux_v I__4383 (
            .O(N__36790),
            .I(N__36781));
    Span4Mux_v I__4382 (
            .O(N__36787),
            .I(N__36778));
    Span4Mux_h I__4381 (
            .O(N__36784),
            .I(N__36775));
    Span4Mux_v I__4380 (
            .O(N__36781),
            .I(N__36770));
    Span4Mux_h I__4379 (
            .O(N__36778),
            .I(N__36770));
    Span4Mux_v I__4378 (
            .O(N__36775),
            .I(N__36767));
    Odrv4 I__4377 (
            .O(N__36770),
            .I(\pid_alt.error_3 ));
    Odrv4 I__4376 (
            .O(N__36767),
            .I(\pid_alt.error_3 ));
    InMux I__4375 (
            .O(N__36762),
            .I(\pid_alt.error_cry_2 ));
    CascadeMux I__4374 (
            .O(N__36759),
            .I(N__36756));
    InMux I__4373 (
            .O(N__36756),
            .I(N__36752));
    InMux I__4372 (
            .O(N__36755),
            .I(N__36749));
    LocalMux I__4371 (
            .O(N__36752),
            .I(N__36746));
    LocalMux I__4370 (
            .O(N__36749),
            .I(alt_command_0));
    Odrv12 I__4369 (
            .O(N__36746),
            .I(alt_command_0));
    InMux I__4368 (
            .O(N__36741),
            .I(N__36738));
    LocalMux I__4367 (
            .O(N__36738),
            .I(N__36733));
    InMux I__4366 (
            .O(N__36737),
            .I(N__36730));
    InMux I__4365 (
            .O(N__36736),
            .I(N__36727));
    Span4Mux_v I__4364 (
            .O(N__36733),
            .I(N__36722));
    LocalMux I__4363 (
            .O(N__36730),
            .I(N__36722));
    LocalMux I__4362 (
            .O(N__36727),
            .I(N__36719));
    Span4Mux_v I__4361 (
            .O(N__36722),
            .I(N__36716));
    Span4Mux_v I__4360 (
            .O(N__36719),
            .I(N__36713));
    Span4Mux_h I__4359 (
            .O(N__36716),
            .I(N__36710));
    Span4Mux_h I__4358 (
            .O(N__36713),
            .I(N__36707));
    Odrv4 I__4357 (
            .O(N__36710),
            .I(\pid_alt.error_4 ));
    Odrv4 I__4356 (
            .O(N__36707),
            .I(\pid_alt.error_4 ));
    InMux I__4355 (
            .O(N__36702),
            .I(\pid_alt.error_cry_3 ));
    CascadeMux I__4354 (
            .O(N__36699),
            .I(N__36696));
    InMux I__4353 (
            .O(N__36696),
            .I(N__36693));
    LocalMux I__4352 (
            .O(N__36693),
            .I(N__36689));
    InMux I__4351 (
            .O(N__36692),
            .I(N__36686));
    Span4Mux_v I__4350 (
            .O(N__36689),
            .I(N__36683));
    LocalMux I__4349 (
            .O(N__36686),
            .I(alt_command_1));
    Odrv4 I__4348 (
            .O(N__36683),
            .I(alt_command_1));
    InMux I__4347 (
            .O(N__36678),
            .I(N__36675));
    LocalMux I__4346 (
            .O(N__36675),
            .I(N__36671));
    InMux I__4345 (
            .O(N__36674),
            .I(N__36667));
    Span4Mux_v I__4344 (
            .O(N__36671),
            .I(N__36664));
    InMux I__4343 (
            .O(N__36670),
            .I(N__36661));
    LocalMux I__4342 (
            .O(N__36667),
            .I(N__36658));
    Span4Mux_v I__4341 (
            .O(N__36664),
            .I(N__36653));
    LocalMux I__4340 (
            .O(N__36661),
            .I(N__36653));
    Span4Mux_s1_h I__4339 (
            .O(N__36658),
            .I(N__36650));
    Span4Mux_h I__4338 (
            .O(N__36653),
            .I(N__36647));
    Span4Mux_h I__4337 (
            .O(N__36650),
            .I(N__36644));
    Span4Mux_v I__4336 (
            .O(N__36647),
            .I(N__36641));
    Span4Mux_v I__4335 (
            .O(N__36644),
            .I(N__36638));
    Odrv4 I__4334 (
            .O(N__36641),
            .I(\pid_alt.error_5 ));
    Odrv4 I__4333 (
            .O(N__36638),
            .I(\pid_alt.error_5 ));
    InMux I__4332 (
            .O(N__36633),
            .I(\pid_alt.error_cry_4 ));
    CascadeMux I__4331 (
            .O(N__36630),
            .I(N__36627));
    InMux I__4330 (
            .O(N__36627),
            .I(N__36623));
    InMux I__4329 (
            .O(N__36626),
            .I(N__36620));
    LocalMux I__4328 (
            .O(N__36623),
            .I(N__36617));
    LocalMux I__4327 (
            .O(N__36620),
            .I(alt_command_2));
    Odrv12 I__4326 (
            .O(N__36617),
            .I(alt_command_2));
    InMux I__4325 (
            .O(N__36612),
            .I(N__36609));
    LocalMux I__4324 (
            .O(N__36609),
            .I(N__36605));
    InMux I__4323 (
            .O(N__36608),
            .I(N__36601));
    Span4Mux_h I__4322 (
            .O(N__36605),
            .I(N__36598));
    InMux I__4321 (
            .O(N__36604),
            .I(N__36595));
    LocalMux I__4320 (
            .O(N__36601),
            .I(N__36592));
    Span4Mux_v I__4319 (
            .O(N__36598),
            .I(N__36589));
    LocalMux I__4318 (
            .O(N__36595),
            .I(N__36586));
    Span4Mux_h I__4317 (
            .O(N__36592),
            .I(N__36583));
    Span4Mux_v I__4316 (
            .O(N__36589),
            .I(N__36580));
    Span12Mux_s4_h I__4315 (
            .O(N__36586),
            .I(N__36577));
    Span4Mux_v I__4314 (
            .O(N__36583),
            .I(N__36574));
    Odrv4 I__4313 (
            .O(N__36580),
            .I(\pid_alt.error_6 ));
    Odrv12 I__4312 (
            .O(N__36577),
            .I(\pid_alt.error_6 ));
    Odrv4 I__4311 (
            .O(N__36574),
            .I(\pid_alt.error_6 ));
    InMux I__4310 (
            .O(N__36567),
            .I(\pid_alt.error_cry_5 ));
    CascadeMux I__4309 (
            .O(N__36564),
            .I(N__36561));
    InMux I__4308 (
            .O(N__36561),
            .I(N__36558));
    LocalMux I__4307 (
            .O(N__36558),
            .I(N__36554));
    InMux I__4306 (
            .O(N__36557),
            .I(N__36551));
    Span4Mux_v I__4305 (
            .O(N__36554),
            .I(N__36548));
    LocalMux I__4304 (
            .O(N__36551),
            .I(alt_command_3));
    Odrv4 I__4303 (
            .O(N__36548),
            .I(alt_command_3));
    InMux I__4302 (
            .O(N__36543),
            .I(N__36540));
    LocalMux I__4301 (
            .O(N__36540),
            .I(N__36537));
    Span4Mux_v I__4300 (
            .O(N__36537),
            .I(N__36532));
    InMux I__4299 (
            .O(N__36536),
            .I(N__36529));
    InMux I__4298 (
            .O(N__36535),
            .I(N__36526));
    Span4Mux_v I__4297 (
            .O(N__36532),
            .I(N__36521));
    LocalMux I__4296 (
            .O(N__36529),
            .I(N__36521));
    LocalMux I__4295 (
            .O(N__36526),
            .I(N__36518));
    Span4Mux_h I__4294 (
            .O(N__36521),
            .I(N__36515));
    Span4Mux_h I__4293 (
            .O(N__36518),
            .I(N__36512));
    Span4Mux_v I__4292 (
            .O(N__36515),
            .I(N__36509));
    Span4Mux_v I__4291 (
            .O(N__36512),
            .I(N__36506));
    Odrv4 I__4290 (
            .O(N__36509),
            .I(\pid_alt.error_7 ));
    Odrv4 I__4289 (
            .O(N__36506),
            .I(\pid_alt.error_7 ));
    InMux I__4288 (
            .O(N__36501),
            .I(\pid_alt.error_cry_6 ));
    InMux I__4287 (
            .O(N__36498),
            .I(N__36493));
    InMux I__4286 (
            .O(N__36497),
            .I(N__36490));
    InMux I__4285 (
            .O(N__36496),
            .I(N__36487));
    LocalMux I__4284 (
            .O(N__36493),
            .I(N__36484));
    LocalMux I__4283 (
            .O(N__36490),
            .I(N__36481));
    LocalMux I__4282 (
            .O(N__36487),
            .I(N__36478));
    Span12Mux_s4_h I__4281 (
            .O(N__36484),
            .I(N__36475));
    Span12Mux_v I__4280 (
            .O(N__36481),
            .I(N__36470));
    Span12Mux_s11_v I__4279 (
            .O(N__36478),
            .I(N__36470));
    Odrv12 I__4278 (
            .O(N__36475),
            .I(\pid_alt.error_8 ));
    Odrv12 I__4277 (
            .O(N__36470),
            .I(\pid_alt.error_8 ));
    InMux I__4276 (
            .O(N__36465),
            .I(bfn_4_19_0_));
    InMux I__4275 (
            .O(N__36462),
            .I(N__36459));
    LocalMux I__4274 (
            .O(N__36459),
            .I(N__36456));
    Span4Mux_v I__4273 (
            .O(N__36456),
            .I(N__36451));
    InMux I__4272 (
            .O(N__36455),
            .I(N__36448));
    InMux I__4271 (
            .O(N__36454),
            .I(N__36445));
    Span4Mux_v I__4270 (
            .O(N__36451),
            .I(N__36440));
    LocalMux I__4269 (
            .O(N__36448),
            .I(N__36440));
    LocalMux I__4268 (
            .O(N__36445),
            .I(N__36437));
    Span4Mux_h I__4267 (
            .O(N__36440),
            .I(N__36434));
    Span4Mux_h I__4266 (
            .O(N__36437),
            .I(N__36431));
    Span4Mux_v I__4265 (
            .O(N__36434),
            .I(N__36428));
    Span4Mux_v I__4264 (
            .O(N__36431),
            .I(N__36425));
    Odrv4 I__4263 (
            .O(N__36428),
            .I(\pid_alt.error_9 ));
    Odrv4 I__4262 (
            .O(N__36425),
            .I(\pid_alt.error_9 ));
    InMux I__4261 (
            .O(N__36420),
            .I(\pid_alt.error_cry_8 ));
    InMux I__4260 (
            .O(N__36417),
            .I(N__36414));
    LocalMux I__4259 (
            .O(N__36414),
            .I(N__36411));
    Span4Mux_v I__4258 (
            .O(N__36411),
            .I(N__36406));
    InMux I__4257 (
            .O(N__36410),
            .I(N__36403));
    InMux I__4256 (
            .O(N__36409),
            .I(N__36400));
    Span4Mux_v I__4255 (
            .O(N__36406),
            .I(N__36395));
    LocalMux I__4254 (
            .O(N__36403),
            .I(N__36395));
    LocalMux I__4253 (
            .O(N__36400),
            .I(N__36392));
    Span4Mux_h I__4252 (
            .O(N__36395),
            .I(N__36389));
    Span4Mux_v I__4251 (
            .O(N__36392),
            .I(N__36386));
    Span4Mux_v I__4250 (
            .O(N__36389),
            .I(N__36383));
    Span4Mux_h I__4249 (
            .O(N__36386),
            .I(N__36380));
    Odrv4 I__4248 (
            .O(N__36383),
            .I(\pid_alt.error_10 ));
    Odrv4 I__4247 (
            .O(N__36380),
            .I(\pid_alt.error_10 ));
    InMux I__4246 (
            .O(N__36375),
            .I(\pid_alt.error_cry_9 ));
    InMux I__4245 (
            .O(N__36372),
            .I(N__36365));
    InMux I__4244 (
            .O(N__36371),
            .I(N__36365));
    InMux I__4243 (
            .O(N__36370),
            .I(N__36362));
    LocalMux I__4242 (
            .O(N__36365),
            .I(N__36359));
    LocalMux I__4241 (
            .O(N__36362),
            .I(N__36356));
    Span4Mux_h I__4240 (
            .O(N__36359),
            .I(N__36353));
    Odrv4 I__4239 (
            .O(N__36356),
            .I(\pid_alt.error_i_reg_esr_RNI15KJZ0Z_14 ));
    Odrv4 I__4238 (
            .O(N__36353),
            .I(\pid_alt.error_i_reg_esr_RNI15KJZ0Z_14 ));
    CascadeMux I__4237 (
            .O(N__36348),
            .I(N__36344));
    CascadeMux I__4236 (
            .O(N__36347),
            .I(N__36341));
    InMux I__4235 (
            .O(N__36344),
            .I(N__36338));
    InMux I__4234 (
            .O(N__36341),
            .I(N__36335));
    LocalMux I__4233 (
            .O(N__36338),
            .I(\pid_alt.error_d_reg_prev_esr_RNIGFN02Z0Z_13 ));
    LocalMux I__4232 (
            .O(N__36335),
            .I(\pid_alt.error_d_reg_prev_esr_RNIGFN02Z0Z_13 ));
    CascadeMux I__4231 (
            .O(N__36330),
            .I(\uart_pc.N_126_li_cascade_ ));
    CascadeMux I__4230 (
            .O(N__36327),
            .I(\uart_pc.N_143_cascade_ ));
    InMux I__4229 (
            .O(N__36324),
            .I(N__36321));
    LocalMux I__4228 (
            .O(N__36321),
            .I(\uart_pc.timer_Count_RNO_0Z0Z_1 ));
    InMux I__4227 (
            .O(N__36318),
            .I(N__36314));
    InMux I__4226 (
            .O(N__36317),
            .I(N__36311));
    LocalMux I__4225 (
            .O(N__36314),
            .I(\pid_alt.drone_altitude_i_0 ));
    LocalMux I__4224 (
            .O(N__36311),
            .I(\pid_alt.drone_altitude_i_0 ));
    InMux I__4223 (
            .O(N__36306),
            .I(N__36303));
    LocalMux I__4222 (
            .O(N__36303),
            .I(\pid_alt.error_axbZ0Z_1 ));
    InMux I__4221 (
            .O(N__36300),
            .I(N__36296));
    InMux I__4220 (
            .O(N__36299),
            .I(N__36292));
    LocalMux I__4219 (
            .O(N__36296),
            .I(N__36289));
    InMux I__4218 (
            .O(N__36295),
            .I(N__36286));
    LocalMux I__4217 (
            .O(N__36292),
            .I(N__36283));
    Span4Mux_v I__4216 (
            .O(N__36289),
            .I(N__36280));
    LocalMux I__4215 (
            .O(N__36286),
            .I(N__36277));
    Span4Mux_v I__4214 (
            .O(N__36283),
            .I(N__36274));
    Span4Mux_v I__4213 (
            .O(N__36280),
            .I(N__36271));
    Span4Mux_v I__4212 (
            .O(N__36277),
            .I(N__36266));
    Span4Mux_v I__4211 (
            .O(N__36274),
            .I(N__36266));
    Span4Mux_h I__4210 (
            .O(N__36271),
            .I(N__36261));
    Span4Mux_h I__4209 (
            .O(N__36266),
            .I(N__36261));
    Odrv4 I__4208 (
            .O(N__36261),
            .I(\pid_alt.error_1 ));
    InMux I__4207 (
            .O(N__36258),
            .I(\pid_alt.error_cry_0 ));
    InMux I__4206 (
            .O(N__36255),
            .I(N__36252));
    LocalMux I__4205 (
            .O(N__36252),
            .I(N__36247));
    InMux I__4204 (
            .O(N__36251),
            .I(N__36244));
    InMux I__4203 (
            .O(N__36250),
            .I(N__36241));
    Span4Mux_v I__4202 (
            .O(N__36247),
            .I(N__36236));
    LocalMux I__4201 (
            .O(N__36244),
            .I(N__36236));
    LocalMux I__4200 (
            .O(N__36241),
            .I(N__36233));
    Span4Mux_v I__4199 (
            .O(N__36236),
            .I(N__36230));
    Span4Mux_h I__4198 (
            .O(N__36233),
            .I(N__36227));
    Span4Mux_h I__4197 (
            .O(N__36230),
            .I(N__36224));
    Span4Mux_v I__4196 (
            .O(N__36227),
            .I(N__36221));
    Odrv4 I__4195 (
            .O(N__36224),
            .I(\pid_alt.error_2 ));
    Odrv4 I__4194 (
            .O(N__36221),
            .I(\pid_alt.error_2 ));
    InMux I__4193 (
            .O(N__36216),
            .I(N__36213));
    LocalMux I__4192 (
            .O(N__36213),
            .I(N__36210));
    Span4Mux_h I__4191 (
            .O(N__36210),
            .I(N__36206));
    InMux I__4190 (
            .O(N__36209),
            .I(N__36203));
    Odrv4 I__4189 (
            .O(N__36206),
            .I(\pid_alt.error_d_reg_prev_esr_RNICISB3Z0Z_3 ));
    LocalMux I__4188 (
            .O(N__36203),
            .I(\pid_alt.error_d_reg_prev_esr_RNICISB3Z0Z_3 ));
    InMux I__4187 (
            .O(N__36198),
            .I(N__36192));
    InMux I__4186 (
            .O(N__36197),
            .I(N__36192));
    LocalMux I__4185 (
            .O(N__36192),
            .I(N__36189));
    Span4Mux_h I__4184 (
            .O(N__36189),
            .I(N__36186));
    Span4Mux_v I__4183 (
            .O(N__36186),
            .I(N__36183));
    Odrv4 I__4182 (
            .O(N__36183),
            .I(\pid_alt.error_d_reg_prev_esr_RNI6P511Z0Z_4 ));
    CascadeMux I__4181 (
            .O(N__36180),
            .I(\pid_alt.error_d_reg_prev_esr_RNI9S511_0Z0Z_5_cascade_ ));
    CascadeMux I__4180 (
            .O(N__36177),
            .I(N__36174));
    InMux I__4179 (
            .O(N__36174),
            .I(N__36171));
    LocalMux I__4178 (
            .O(N__36171),
            .I(\pid_alt.error_d_reg_prev_esr_RNIOGSO6Z0Z_4 ));
    InMux I__4177 (
            .O(N__36168),
            .I(N__36165));
    LocalMux I__4176 (
            .O(N__36165),
            .I(\pid_alt.error_d_reg_prev_esr_RNI88G14Z0Z_14 ));
    InMux I__4175 (
            .O(N__36162),
            .I(N__36159));
    LocalMux I__4174 (
            .O(N__36159),
            .I(\pid_alt.error_d_reg_prev_esr_RNIPMHMZ0Z_14 ));
    CascadeMux I__4173 (
            .O(N__36156),
            .I(\pid_alt.error_d_reg_prev_esr_RNIPMHMZ0Z_14_cascade_ ));
    InMux I__4172 (
            .O(N__36153),
            .I(N__36146));
    InMux I__4171 (
            .O(N__36152),
            .I(N__36146));
    InMux I__4170 (
            .O(N__36151),
            .I(N__36143));
    LocalMux I__4169 (
            .O(N__36146),
            .I(N__36140));
    LocalMux I__4168 (
            .O(N__36143),
            .I(N__36137));
    Span4Mux_h I__4167 (
            .O(N__36140),
            .I(N__36134));
    Odrv4 I__4166 (
            .O(N__36137),
            .I(\pid_alt.error_i_reg_esr_RNI38LJZ0Z_15 ));
    Odrv4 I__4165 (
            .O(N__36134),
            .I(\pid_alt.error_i_reg_esr_RNI38LJZ0Z_15 ));
    InMux I__4164 (
            .O(N__36129),
            .I(N__36126));
    LocalMux I__4163 (
            .O(N__36126),
            .I(N__36123));
    Span4Mux_v I__4162 (
            .O(N__36123),
            .I(N__36120));
    Span4Mux_h I__4161 (
            .O(N__36120),
            .I(N__36116));
    CascadeMux I__4160 (
            .O(N__36119),
            .I(N__36113));
    Span4Mux_v I__4159 (
            .O(N__36116),
            .I(N__36110));
    InMux I__4158 (
            .O(N__36113),
            .I(N__36107));
    Odrv4 I__4157 (
            .O(N__36110),
            .I(\pid_alt.error_d_reg_prev_esr_RNIOOO02Z0Z_14 ));
    LocalMux I__4156 (
            .O(N__36107),
            .I(\pid_alt.error_d_reg_prev_esr_RNIOOO02Z0Z_14 ));
    InMux I__4155 (
            .O(N__36102),
            .I(N__36096));
    InMux I__4154 (
            .O(N__36101),
            .I(N__36096));
    LocalMux I__4153 (
            .O(N__36096),
            .I(\pid_alt.error_d_reg_prev_esr_RNISPHM_0Z0Z_15 ));
    InMux I__4152 (
            .O(N__36093),
            .I(N__36087));
    InMux I__4151 (
            .O(N__36092),
            .I(N__36087));
    LocalMux I__4150 (
            .O(N__36087),
            .I(N__36084));
    Span4Mux_h I__4149 (
            .O(N__36084),
            .I(N__36081));
    Span4Mux_v I__4148 (
            .O(N__36081),
            .I(N__36078));
    Odrv4 I__4147 (
            .O(N__36078),
            .I(\pid_alt.error_p_regZ0Z_14 ));
    CascadeMux I__4146 (
            .O(N__36075),
            .I(\pid_alt.error_d_reg_prev_esr_RNIPMHM_0Z0Z_14_cascade_ ));
    InMux I__4145 (
            .O(N__36072),
            .I(N__36069));
    LocalMux I__4144 (
            .O(N__36069),
            .I(\pid_alt.error_d_reg_prev_esr_RNICQF44Z0Z_13 ));
    InMux I__4143 (
            .O(N__36066),
            .I(N__36057));
    InMux I__4142 (
            .O(N__36065),
            .I(N__36057));
    InMux I__4141 (
            .O(N__36064),
            .I(N__36057));
    LocalMux I__4140 (
            .O(N__36057),
            .I(N__36054));
    Span12Mux_h I__4139 (
            .O(N__36054),
            .I(N__36051));
    Span12Mux_v I__4138 (
            .O(N__36051),
            .I(N__36048));
    Odrv12 I__4137 (
            .O(N__36048),
            .I(\pid_alt.error_d_regZ0Z_14 ));
    CascadeMux I__4136 (
            .O(N__36045),
            .I(N__36042));
    InMux I__4135 (
            .O(N__36042),
            .I(N__36036));
    InMux I__4134 (
            .O(N__36041),
            .I(N__36036));
    LocalMux I__4133 (
            .O(N__36036),
            .I(\pid_alt.error_d_reg_prevZ0Z_14 ));
    InMux I__4132 (
            .O(N__36033),
            .I(N__36030));
    LocalMux I__4131 (
            .O(N__36030),
            .I(\pid_alt.error_d_reg_prev_esr_RNIPMHM_0Z0Z_14 ));
    InMux I__4130 (
            .O(N__36027),
            .I(N__36021));
    InMux I__4129 (
            .O(N__36026),
            .I(N__36021));
    LocalMux I__4128 (
            .O(N__36021),
            .I(N__36018));
    Span4Mux_h I__4127 (
            .O(N__36018),
            .I(N__36015));
    Odrv4 I__4126 (
            .O(N__36015),
            .I(\pid_alt.error_d_reg_prev_esr_RNIMJHMZ0Z_13 ));
    InMux I__4125 (
            .O(N__36012),
            .I(N__36009));
    LocalMux I__4124 (
            .O(N__36009),
            .I(N__36006));
    Span4Mux_h I__4123 (
            .O(N__36006),
            .I(N__36003));
    Odrv4 I__4122 (
            .O(N__36003),
            .I(\Commands_frame_decoder.state_ns_i_a2_0_2_0 ));
    CascadeMux I__4121 (
            .O(N__36000),
            .I(\pid_alt.error_d_reg_prev_esr_RNI9S511Z0Z_5_cascade_ ));
    InMux I__4120 (
            .O(N__35997),
            .I(N__35994));
    LocalMux I__4119 (
            .O(N__35994),
            .I(N__35991));
    Span4Mux_v I__4118 (
            .O(N__35991),
            .I(N__35987));
    InMux I__4117 (
            .O(N__35990),
            .I(N__35984));
    Odrv4 I__4116 (
            .O(N__35987),
            .I(\pid_alt.error_d_reg_prev_esr_RNIL81T2Z0Z_5 ));
    LocalMux I__4115 (
            .O(N__35984),
            .I(\pid_alt.error_d_reg_prev_esr_RNIL81T2Z0Z_5 ));
    InMux I__4114 (
            .O(N__35979),
            .I(N__35975));
    InMux I__4113 (
            .O(N__35978),
            .I(N__35972));
    LocalMux I__4112 (
            .O(N__35975),
            .I(N__35969));
    LocalMux I__4111 (
            .O(N__35972),
            .I(N__35966));
    Span4Mux_v I__4110 (
            .O(N__35969),
            .I(N__35961));
    Span4Mux_h I__4109 (
            .O(N__35966),
            .I(N__35961));
    Span4Mux_v I__4108 (
            .O(N__35961),
            .I(N__35958));
    Odrv4 I__4107 (
            .O(N__35958),
            .I(\pid_alt.error_p_regZ0Z_6 ));
    InMux I__4106 (
            .O(N__35955),
            .I(N__35952));
    LocalMux I__4105 (
            .O(N__35952),
            .I(N__35948));
    InMux I__4104 (
            .O(N__35951),
            .I(N__35945));
    Span4Mux_h I__4103 (
            .O(N__35948),
            .I(N__35942));
    LocalMux I__4102 (
            .O(N__35945),
            .I(\pid_alt.error_d_reg_prevZ0Z_6 ));
    Odrv4 I__4101 (
            .O(N__35942),
            .I(\pid_alt.error_d_reg_prevZ0Z_6 ));
    InMux I__4100 (
            .O(N__35937),
            .I(N__35932));
    InMux I__4099 (
            .O(N__35936),
            .I(N__35927));
    InMux I__4098 (
            .O(N__35935),
            .I(N__35927));
    LocalMux I__4097 (
            .O(N__35932),
            .I(N__35924));
    LocalMux I__4096 (
            .O(N__35927),
            .I(N__35921));
    Span4Mux_v I__4095 (
            .O(N__35924),
            .I(N__35918));
    Span4Mux_v I__4094 (
            .O(N__35921),
            .I(N__35915));
    Span4Mux_h I__4093 (
            .O(N__35918),
            .I(N__35912));
    Span4Mux_v I__4092 (
            .O(N__35915),
            .I(N__35909));
    Span4Mux_v I__4091 (
            .O(N__35912),
            .I(N__35906));
    Odrv4 I__4090 (
            .O(N__35909),
            .I(\pid_alt.error_d_regZ0Z_6 ));
    Odrv4 I__4089 (
            .O(N__35906),
            .I(\pid_alt.error_d_regZ0Z_6 ));
    InMux I__4088 (
            .O(N__35901),
            .I(N__35898));
    LocalMux I__4087 (
            .O(N__35898),
            .I(\pid_alt.error_d_reg_prev_esr_RNICV511_0Z0Z_6 ));
    InMux I__4086 (
            .O(N__35895),
            .I(N__35892));
    LocalMux I__4085 (
            .O(N__35892),
            .I(\pid_alt.error_d_reg_prev_esr_RNI9S511Z0Z_5 ));
    CascadeMux I__4084 (
            .O(N__35889),
            .I(\pid_alt.error_d_reg_prev_esr_RNICV511_0Z0Z_6_cascade_ ));
    InMux I__4083 (
            .O(N__35886),
            .I(N__35881));
    InMux I__4082 (
            .O(N__35885),
            .I(N__35876));
    InMux I__4081 (
            .O(N__35884),
            .I(N__35876));
    LocalMux I__4080 (
            .O(N__35881),
            .I(N__35873));
    LocalMux I__4079 (
            .O(N__35876),
            .I(N__35870));
    Span4Mux_v I__4078 (
            .O(N__35873),
            .I(N__35867));
    Span4Mux_h I__4077 (
            .O(N__35870),
            .I(N__35864));
    Odrv4 I__4076 (
            .O(N__35867),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_5_c_RNI0DLQ ));
    Odrv4 I__4075 (
            .O(N__35864),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_5_c_RNI0DLQ ));
    InMux I__4074 (
            .O(N__35859),
            .I(N__35856));
    LocalMux I__4073 (
            .O(N__35856),
            .I(\pid_alt.error_d_reg_prev_esr_RNI171A6Z0Z_5 ));
    CascadeMux I__4072 (
            .O(N__35853),
            .I(N__35849));
    InMux I__4071 (
            .O(N__35852),
            .I(N__35846));
    InMux I__4070 (
            .O(N__35849),
            .I(N__35843));
    LocalMux I__4069 (
            .O(N__35846),
            .I(\pid_alt.error_d_reg_prev_esr_RNICUVC3Z0Z_4 ));
    LocalMux I__4068 (
            .O(N__35843),
            .I(\pid_alt.error_d_reg_prev_esr_RNICUVC3Z0Z_4 ));
    InMux I__4067 (
            .O(N__35838),
            .I(N__35829));
    InMux I__4066 (
            .O(N__35837),
            .I(N__35829));
    InMux I__4065 (
            .O(N__35836),
            .I(N__35829));
    LocalMux I__4064 (
            .O(N__35829),
            .I(N__35826));
    Span4Mux_v I__4063 (
            .O(N__35826),
            .I(N__35823));
    Span4Mux_v I__4062 (
            .O(N__35823),
            .I(N__35820));
    Odrv4 I__4061 (
            .O(N__35820),
            .I(\pid_alt.error_d_regZ0Z_5 ));
    CascadeMux I__4060 (
            .O(N__35817),
            .I(N__35814));
    InMux I__4059 (
            .O(N__35814),
            .I(N__35808));
    InMux I__4058 (
            .O(N__35813),
            .I(N__35808));
    LocalMux I__4057 (
            .O(N__35808),
            .I(\pid_alt.error_d_reg_prevZ0Z_5 ));
    InMux I__4056 (
            .O(N__35805),
            .I(N__35799));
    InMux I__4055 (
            .O(N__35804),
            .I(N__35799));
    LocalMux I__4054 (
            .O(N__35799),
            .I(N__35796));
    Span4Mux_h I__4053 (
            .O(N__35796),
            .I(N__35793));
    Span4Mux_v I__4052 (
            .O(N__35793),
            .I(N__35790));
    Odrv4 I__4051 (
            .O(N__35790),
            .I(\pid_alt.error_p_regZ0Z_5 ));
    InMux I__4050 (
            .O(N__35787),
            .I(N__35784));
    LocalMux I__4049 (
            .O(N__35784),
            .I(\pid_alt.error_d_reg_prev_esr_RNI9S511_0Z0Z_5 ));
    CascadeMux I__4048 (
            .O(N__35781),
            .I(N__35774));
    InMux I__4047 (
            .O(N__35780),
            .I(N__35760));
    InMux I__4046 (
            .O(N__35779),
            .I(N__35760));
    InMux I__4045 (
            .O(N__35778),
            .I(N__35760));
    InMux I__4044 (
            .O(N__35777),
            .I(N__35760));
    InMux I__4043 (
            .O(N__35774),
            .I(N__35760));
    InMux I__4042 (
            .O(N__35773),
            .I(N__35760));
    LocalMux I__4041 (
            .O(N__35760),
            .I(\uart_pc.timer_Count_RNIMQ8T1Z0Z_2 ));
    InMux I__4040 (
            .O(N__35757),
            .I(N__35747));
    InMux I__4039 (
            .O(N__35756),
            .I(N__35734));
    InMux I__4038 (
            .O(N__35755),
            .I(N__35734));
    InMux I__4037 (
            .O(N__35754),
            .I(N__35734));
    InMux I__4036 (
            .O(N__35753),
            .I(N__35734));
    InMux I__4035 (
            .O(N__35752),
            .I(N__35734));
    InMux I__4034 (
            .O(N__35751),
            .I(N__35734));
    InMux I__4033 (
            .O(N__35750),
            .I(N__35731));
    LocalMux I__4032 (
            .O(N__35747),
            .I(N__35728));
    LocalMux I__4031 (
            .O(N__35734),
            .I(\uart_pc.timer_Count_RNILR1B2Z0Z_2 ));
    LocalMux I__4030 (
            .O(N__35731),
            .I(\uart_pc.timer_Count_RNILR1B2Z0Z_2 ));
    Odrv4 I__4029 (
            .O(N__35728),
            .I(\uart_pc.timer_Count_RNILR1B2Z0Z_2 ));
    CascadeMux I__4028 (
            .O(N__35721),
            .I(\uart_pc.timer_Count_RNIMQ8T1Z0Z_2_cascade_ ));
    CascadeMux I__4027 (
            .O(N__35718),
            .I(\Commands_frame_decoder.source_CH1data8lto7Z0Z_2_cascade_ ));
    CascadeMux I__4026 (
            .O(N__35715),
            .I(\Commands_frame_decoder.source_CH1data8_cascade_ ));
    CascadeMux I__4025 (
            .O(N__35712),
            .I(N__35708));
    InMux I__4024 (
            .O(N__35711),
            .I(N__35700));
    InMux I__4023 (
            .O(N__35708),
            .I(N__35700));
    InMux I__4022 (
            .O(N__35707),
            .I(N__35700));
    LocalMux I__4021 (
            .O(N__35700),
            .I(\Commands_frame_decoder.source_CH1data8 ));
    CascadeMux I__4020 (
            .O(N__35697),
            .I(N__35694));
    InMux I__4019 (
            .O(N__35694),
            .I(N__35688));
    InMux I__4018 (
            .O(N__35693),
            .I(N__35688));
    LocalMux I__4017 (
            .O(N__35688),
            .I(\pid_alt.source_pid_1_sqmuxa_0_a2_0_2 ));
    InMux I__4016 (
            .O(N__35685),
            .I(N__35682));
    LocalMux I__4015 (
            .O(N__35682),
            .I(\Commands_frame_decoder.state_ns_0_a3_0_1Z0Z_2 ));
    InMux I__4014 (
            .O(N__35679),
            .I(N__35675));
    InMux I__4013 (
            .O(N__35678),
            .I(N__35672));
    LocalMux I__4012 (
            .O(N__35675),
            .I(N__35669));
    LocalMux I__4011 (
            .O(N__35672),
            .I(N__35666));
    Odrv4 I__4010 (
            .O(N__35669),
            .I(\Commands_frame_decoder.source_CH4data_1_sqmuxa ));
    Odrv12 I__4009 (
            .O(N__35666),
            .I(\Commands_frame_decoder.source_CH4data_1_sqmuxa ));
    CascadeMux I__4008 (
            .O(N__35661),
            .I(N__35657));
    InMux I__4007 (
            .O(N__35660),
            .I(N__35654));
    InMux I__4006 (
            .O(N__35657),
            .I(N__35651));
    LocalMux I__4005 (
            .O(N__35654),
            .I(N__35648));
    LocalMux I__4004 (
            .O(N__35651),
            .I(\pid_alt.pid_preregZ0Z_5 ));
    Odrv4 I__4003 (
            .O(N__35648),
            .I(\pid_alt.pid_preregZ0Z_5 ));
    InMux I__4002 (
            .O(N__35643),
            .I(N__35637));
    InMux I__4001 (
            .O(N__35642),
            .I(N__35632));
    InMux I__4000 (
            .O(N__35641),
            .I(N__35632));
    InMux I__3999 (
            .O(N__35640),
            .I(N__35629));
    LocalMux I__3998 (
            .O(N__35637),
            .I(N__35624));
    LocalMux I__3997 (
            .O(N__35632),
            .I(N__35624));
    LocalMux I__3996 (
            .O(N__35629),
            .I(\pid_alt.N_154 ));
    Odrv4 I__3995 (
            .O(N__35624),
            .I(\pid_alt.N_154 ));
    CascadeMux I__3994 (
            .O(N__35619),
            .I(\pid_alt.N_57_cascade_ ));
    InMux I__3993 (
            .O(N__35616),
            .I(N__35613));
    LocalMux I__3992 (
            .O(N__35613),
            .I(\pid_alt.un1_reset_1 ));
    CascadeMux I__3991 (
            .O(N__35610),
            .I(N__35607));
    InMux I__3990 (
            .O(N__35607),
            .I(N__35604));
    LocalMux I__3989 (
            .O(N__35604),
            .I(\pid_alt.source_pid_1_sqmuxa_0_a2_1_7 ));
    InMux I__3988 (
            .O(N__35601),
            .I(N__35598));
    LocalMux I__3987 (
            .O(N__35598),
            .I(\pid_alt.N_51 ));
    InMux I__3986 (
            .O(N__35595),
            .I(N__35589));
    InMux I__3985 (
            .O(N__35594),
            .I(N__35589));
    LocalMux I__3984 (
            .O(N__35589),
            .I(N__35586));
    Span4Mux_v I__3983 (
            .O(N__35586),
            .I(N__35583));
    Odrv4 I__3982 (
            .O(N__35583),
            .I(\pid_alt.N_52 ));
    InMux I__3981 (
            .O(N__35580),
            .I(N__35575));
    InMux I__3980 (
            .O(N__35579),
            .I(N__35570));
    InMux I__3979 (
            .O(N__35578),
            .I(N__35570));
    LocalMux I__3978 (
            .O(N__35575),
            .I(N__35563));
    LocalMux I__3977 (
            .O(N__35570),
            .I(N__35563));
    InMux I__3976 (
            .O(N__35569),
            .I(N__35558));
    InMux I__3975 (
            .O(N__35568),
            .I(N__35558));
    Span4Mux_v I__3974 (
            .O(N__35563),
            .I(N__35555));
    LocalMux I__3973 (
            .O(N__35558),
            .I(\pid_alt.pid_preregZ0Z_4 ));
    Odrv4 I__3972 (
            .O(N__35555),
            .I(\pid_alt.pid_preregZ0Z_4 ));
    CascadeMux I__3971 (
            .O(N__35550),
            .I(\pid_alt.N_52_cascade_ ));
    CascadeMux I__3970 (
            .O(N__35547),
            .I(\pid_alt.N_54_cascade_ ));
    CascadeMux I__3969 (
            .O(N__35544),
            .I(N__35540));
    InMux I__3968 (
            .O(N__35543),
            .I(N__35532));
    InMux I__3967 (
            .O(N__35540),
            .I(N__35532));
    InMux I__3966 (
            .O(N__35539),
            .I(N__35532));
    LocalMux I__3965 (
            .O(N__35532),
            .I(\pid_alt.N_54 ));
    CEMux I__3964 (
            .O(N__35529),
            .I(N__35526));
    LocalMux I__3963 (
            .O(N__35526),
            .I(N__35521));
    CEMux I__3962 (
            .O(N__35525),
            .I(N__35518));
    CEMux I__3961 (
            .O(N__35524),
            .I(N__35515));
    Span4Mux_v I__3960 (
            .O(N__35521),
            .I(N__35510));
    LocalMux I__3959 (
            .O(N__35518),
            .I(N__35510));
    LocalMux I__3958 (
            .O(N__35515),
            .I(N__35507));
    Span4Mux_v I__3957 (
            .O(N__35510),
            .I(N__35504));
    Span4Mux_h I__3956 (
            .O(N__35507),
            .I(N__35501));
    Odrv4 I__3955 (
            .O(N__35504),
            .I(\pid_alt.N_72_i_1 ));
    Odrv4 I__3954 (
            .O(N__35501),
            .I(\pid_alt.N_72_i_1 ));
    InMux I__3953 (
            .O(N__35496),
            .I(N__35490));
    InMux I__3952 (
            .O(N__35495),
            .I(N__35490));
    LocalMux I__3951 (
            .O(N__35490),
            .I(N__35487));
    Span4Mux_h I__3950 (
            .O(N__35487),
            .I(N__35484));
    Odrv4 I__3949 (
            .O(N__35484),
            .I(\pid_alt.pid_preregZ0Z_2 ));
    CascadeMux I__3948 (
            .O(N__35481),
            .I(N__35478));
    InMux I__3947 (
            .O(N__35478),
            .I(N__35472));
    InMux I__3946 (
            .O(N__35477),
            .I(N__35472));
    LocalMux I__3945 (
            .O(N__35472),
            .I(N__35469));
    Span4Mux_h I__3944 (
            .O(N__35469),
            .I(N__35466));
    Odrv4 I__3943 (
            .O(N__35466),
            .I(\pid_alt.pid_preregZ0Z_1 ));
    CascadeMux I__3942 (
            .O(N__35463),
            .I(N__35459));
    InMux I__3941 (
            .O(N__35462),
            .I(N__35454));
    InMux I__3940 (
            .O(N__35459),
            .I(N__35454));
    LocalMux I__3939 (
            .O(N__35454),
            .I(N__35451));
    Span4Mux_h I__3938 (
            .O(N__35451),
            .I(N__35448));
    Odrv4 I__3937 (
            .O(N__35448),
            .I(\pid_alt.pid_preregZ0Z_3 ));
    InMux I__3936 (
            .O(N__35445),
            .I(N__35439));
    InMux I__3935 (
            .O(N__35444),
            .I(N__35439));
    LocalMux I__3934 (
            .O(N__35439),
            .I(N__35436));
    Span4Mux_h I__3933 (
            .O(N__35436),
            .I(N__35433));
    Odrv4 I__3932 (
            .O(N__35433),
            .I(\pid_alt.pid_preregZ0Z_0 ));
    InMux I__3931 (
            .O(N__35430),
            .I(N__35427));
    LocalMux I__3930 (
            .O(N__35427),
            .I(\pid_alt.error_i_acumm_preregZ0Z_15 ));
    CascadeMux I__3929 (
            .O(N__35424),
            .I(N__35421));
    InMux I__3928 (
            .O(N__35421),
            .I(N__35417));
    InMux I__3927 (
            .O(N__35420),
            .I(N__35414));
    LocalMux I__3926 (
            .O(N__35417),
            .I(N__35410));
    LocalMux I__3925 (
            .O(N__35414),
            .I(N__35407));
    InMux I__3924 (
            .O(N__35413),
            .I(N__35404));
    Span4Mux_v I__3923 (
            .O(N__35410),
            .I(N__35401));
    Span4Mux_v I__3922 (
            .O(N__35407),
            .I(N__35398));
    LocalMux I__3921 (
            .O(N__35404),
            .I(N__35393));
    Span4Mux_s3_h I__3920 (
            .O(N__35401),
            .I(N__35393));
    Odrv4 I__3919 (
            .O(N__35398),
            .I(\pid_alt.error_i_acumm_esr_RNI0VF91Z0Z_3 ));
    Odrv4 I__3918 (
            .O(N__35393),
            .I(\pid_alt.error_i_acumm_esr_RNI0VF91Z0Z_3 ));
    CascadeMux I__3917 (
            .O(N__35388),
            .I(\pid_alt.un1_reset_0_i_cascade_ ));
    CascadeMux I__3916 (
            .O(N__35385),
            .I(\pid_alt.source_pid_1_sqmuxa_0_o2_3_cascade_ ));
    CascadeMux I__3915 (
            .O(N__35382),
            .I(\pid_alt.N_51_cascade_ ));
    InMux I__3914 (
            .O(N__35379),
            .I(N__35376));
    LocalMux I__3913 (
            .O(N__35376),
            .I(\pid_alt.source_pid_1_sqmuxa_0_a2_0_3 ));
    CascadeMux I__3912 (
            .O(N__35373),
            .I(\pid_alt.error_d_reg_prev_esr_RNIVSHMZ0Z_16_cascade_ ));
    InMux I__3911 (
            .O(N__35370),
            .I(N__35365));
    InMux I__3910 (
            .O(N__35369),
            .I(N__35360));
    InMux I__3909 (
            .O(N__35368),
            .I(N__35360));
    LocalMux I__3908 (
            .O(N__35365),
            .I(\pid_alt.error_i_reg_esr_RNI7ENJZ0Z_17 ));
    LocalMux I__3907 (
            .O(N__35360),
            .I(\pid_alt.error_i_reg_esr_RNI7ENJZ0Z_17 ));
    CascadeMux I__3906 (
            .O(N__35355),
            .I(N__35352));
    InMux I__3905 (
            .O(N__35352),
            .I(N__35349));
    LocalMux I__3904 (
            .O(N__35349),
            .I(N__35346));
    Odrv12 I__3903 (
            .O(N__35346),
            .I(\pid_alt.error_d_reg_prev_esr_RNI8DL14Z0Z_16 ));
    InMux I__3902 (
            .O(N__35343),
            .I(N__35339));
    InMux I__3901 (
            .O(N__35342),
            .I(N__35336));
    LocalMux I__3900 (
            .O(N__35339),
            .I(N__35333));
    LocalMux I__3899 (
            .O(N__35336),
            .I(\pid_alt.error_d_reg_prev_esr_RNI02Q02Z0Z_15 ));
    Odrv12 I__3898 (
            .O(N__35333),
            .I(\pid_alt.error_d_reg_prev_esr_RNI02Q02Z0Z_15 ));
    InMux I__3897 (
            .O(N__35328),
            .I(N__35322));
    InMux I__3896 (
            .O(N__35327),
            .I(N__35322));
    LocalMux I__3895 (
            .O(N__35322),
            .I(N__35319));
    Span4Mux_h I__3894 (
            .O(N__35319),
            .I(N__35316));
    Odrv4 I__3893 (
            .O(N__35316),
            .I(\pid_alt.error_p_regZ0Z_16 ));
    CascadeMux I__3892 (
            .O(N__35313),
            .I(N__35310));
    InMux I__3891 (
            .O(N__35310),
            .I(N__35304));
    InMux I__3890 (
            .O(N__35309),
            .I(N__35304));
    LocalMux I__3889 (
            .O(N__35304),
            .I(\pid_alt.error_d_reg_prevZ0Z_16 ));
    InMux I__3888 (
            .O(N__35301),
            .I(N__35292));
    InMux I__3887 (
            .O(N__35300),
            .I(N__35292));
    InMux I__3886 (
            .O(N__35299),
            .I(N__35292));
    LocalMux I__3885 (
            .O(N__35292),
            .I(N__35289));
    Span4Mux_v I__3884 (
            .O(N__35289),
            .I(N__35286));
    Span4Mux_v I__3883 (
            .O(N__35286),
            .I(N__35283));
    Span4Mux_v I__3882 (
            .O(N__35283),
            .I(N__35280));
    Span4Mux_v I__3881 (
            .O(N__35280),
            .I(N__35277));
    Odrv4 I__3880 (
            .O(N__35277),
            .I(\pid_alt.error_d_regZ0Z_16 ));
    InMux I__3879 (
            .O(N__35274),
            .I(N__35271));
    LocalMux I__3878 (
            .O(N__35271),
            .I(\pid_alt.error_d_reg_prev_esr_RNIVSHM_0Z0Z_16 ));
    CascadeMux I__3877 (
            .O(N__35268),
            .I(\pid_alt.error_d_reg_prev_esr_RNIVSHM_0Z0Z_16_cascade_ ));
    InMux I__3876 (
            .O(N__35265),
            .I(N__35262));
    LocalMux I__3875 (
            .O(N__35262),
            .I(N__35257));
    InMux I__3874 (
            .O(N__35261),
            .I(N__35252));
    InMux I__3873 (
            .O(N__35260),
            .I(N__35252));
    Odrv4 I__3872 (
            .O(N__35257),
            .I(\pid_alt.error_i_reg_esr_RNI5BMJZ0Z_16 ));
    LocalMux I__3871 (
            .O(N__35252),
            .I(\pid_alt.error_i_reg_esr_RNI5BMJZ0Z_16 ));
    InMux I__3870 (
            .O(N__35247),
            .I(N__35244));
    LocalMux I__3869 (
            .O(N__35244),
            .I(N__35241));
    Odrv12 I__3868 (
            .O(N__35241),
            .I(\pid_alt.error_d_reg_prev_esr_RNIOQI14Z0Z_15 ));
    InMux I__3867 (
            .O(N__35238),
            .I(N__35235));
    LocalMux I__3866 (
            .O(N__35235),
            .I(N__35230));
    InMux I__3865 (
            .O(N__35234),
            .I(N__35225));
    InMux I__3864 (
            .O(N__35233),
            .I(N__35225));
    Span4Mux_v I__3863 (
            .O(N__35230),
            .I(N__35222));
    LocalMux I__3862 (
            .O(N__35225),
            .I(N__35219));
    Odrv4 I__3861 (
            .O(N__35222),
            .I(\pid_alt.error_i_acumm_esr_RNI33H91Z0Z_4 ));
    Odrv4 I__3860 (
            .O(N__35219),
            .I(\pid_alt.error_i_acumm_esr_RNI33H91Z0Z_4 ));
    CascadeMux I__3859 (
            .O(N__35214),
            .I(N__35209));
    InMux I__3858 (
            .O(N__35213),
            .I(N__35206));
    InMux I__3857 (
            .O(N__35212),
            .I(N__35203));
    InMux I__3856 (
            .O(N__35209),
            .I(N__35200));
    LocalMux I__3855 (
            .O(N__35206),
            .I(N__35197));
    LocalMux I__3854 (
            .O(N__35203),
            .I(N__35192));
    LocalMux I__3853 (
            .O(N__35200),
            .I(N__35192));
    Span4Mux_v I__3852 (
            .O(N__35197),
            .I(N__35189));
    Span4Mux_h I__3851 (
            .O(N__35192),
            .I(N__35186));
    Odrv4 I__3850 (
            .O(N__35189),
            .I(\pid_alt.error_i_acumm_esr_RNITQE91Z0Z_2 ));
    Odrv4 I__3849 (
            .O(N__35186),
            .I(\pid_alt.error_i_acumm_esr_RNITQE91Z0Z_2 ));
    CascadeMux I__3848 (
            .O(N__35181),
            .I(N__35174));
    InMux I__3847 (
            .O(N__35180),
            .I(N__35170));
    InMux I__3846 (
            .O(N__35179),
            .I(N__35165));
    InMux I__3845 (
            .O(N__35178),
            .I(N__35165));
    InMux I__3844 (
            .O(N__35177),
            .I(N__35158));
    InMux I__3843 (
            .O(N__35174),
            .I(N__35158));
    InMux I__3842 (
            .O(N__35173),
            .I(N__35158));
    LocalMux I__3841 (
            .O(N__35170),
            .I(\pid_alt.error_d_reg_prevZ0Z_20 ));
    LocalMux I__3840 (
            .O(N__35165),
            .I(\pid_alt.error_d_reg_prevZ0Z_20 ));
    LocalMux I__3839 (
            .O(N__35158),
            .I(\pid_alt.error_d_reg_prevZ0Z_20 ));
    InMux I__3838 (
            .O(N__35151),
            .I(N__35147));
    InMux I__3837 (
            .O(N__35150),
            .I(N__35144));
    LocalMux I__3836 (
            .O(N__35147),
            .I(N__35134));
    LocalMux I__3835 (
            .O(N__35144),
            .I(N__35134));
    InMux I__3834 (
            .O(N__35143),
            .I(N__35129));
    InMux I__3833 (
            .O(N__35142),
            .I(N__35129));
    InMux I__3832 (
            .O(N__35141),
            .I(N__35122));
    InMux I__3831 (
            .O(N__35140),
            .I(N__35122));
    InMux I__3830 (
            .O(N__35139),
            .I(N__35122));
    Sp12to4 I__3829 (
            .O(N__35134),
            .I(N__35115));
    LocalMux I__3828 (
            .O(N__35129),
            .I(N__35115));
    LocalMux I__3827 (
            .O(N__35122),
            .I(N__35115));
    Span12Mux_v I__3826 (
            .O(N__35115),
            .I(N__35112));
    Span12Mux_v I__3825 (
            .O(N__35112),
            .I(N__35109));
    Odrv12 I__3824 (
            .O(N__35109),
            .I(\pid_alt.error_d_regZ0Z_20 ));
    CascadeMux I__3823 (
            .O(N__35106),
            .I(N__35100));
    CascadeMux I__3822 (
            .O(N__35105),
            .I(N__35097));
    CascadeMux I__3821 (
            .O(N__35104),
            .I(N__35094));
    InMux I__3820 (
            .O(N__35103),
            .I(N__35089));
    InMux I__3819 (
            .O(N__35100),
            .I(N__35084));
    InMux I__3818 (
            .O(N__35097),
            .I(N__35084));
    InMux I__3817 (
            .O(N__35094),
            .I(N__35077));
    InMux I__3816 (
            .O(N__35093),
            .I(N__35077));
    InMux I__3815 (
            .O(N__35092),
            .I(N__35077));
    LocalMux I__3814 (
            .O(N__35089),
            .I(N__35072));
    LocalMux I__3813 (
            .O(N__35084),
            .I(N__35072));
    LocalMux I__3812 (
            .O(N__35077),
            .I(N__35069));
    Span4Mux_h I__3811 (
            .O(N__35072),
            .I(N__35066));
    Span4Mux_h I__3810 (
            .O(N__35069),
            .I(N__35063));
    Odrv4 I__3809 (
            .O(N__35066),
            .I(\pid_alt.error_p_regZ0Z_20 ));
    Odrv4 I__3808 (
            .O(N__35063),
            .I(\pid_alt.error_p_regZ0Z_20 ));
    InMux I__3807 (
            .O(N__35058),
            .I(N__35051));
    InMux I__3806 (
            .O(N__35057),
            .I(N__35046));
    InMux I__3805 (
            .O(N__35056),
            .I(N__35046));
    InMux I__3804 (
            .O(N__35055),
            .I(N__35041));
    InMux I__3803 (
            .O(N__35054),
            .I(N__35041));
    LocalMux I__3802 (
            .O(N__35051),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_20_c_RNISVKK ));
    LocalMux I__3801 (
            .O(N__35046),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_20_c_RNISVKK ));
    LocalMux I__3800 (
            .O(N__35041),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_20_c_RNISVKK ));
    CascadeMux I__3799 (
            .O(N__35034),
            .I(N__35031));
    InMux I__3798 (
            .O(N__35031),
            .I(N__35028));
    LocalMux I__3797 (
            .O(N__35028),
            .I(N__35025));
    Odrv4 I__3796 (
            .O(N__35025),
            .I(\pid_alt.error_d_reg_prev_esr_RNICG9B1_2Z0Z_20 ));
    InMux I__3795 (
            .O(N__35022),
            .I(N__35019));
    LocalMux I__3794 (
            .O(N__35019),
            .I(N__35015));
    InMux I__3793 (
            .O(N__35018),
            .I(N__35012));
    Span4Mux_h I__3792 (
            .O(N__35015),
            .I(N__35009));
    LocalMux I__3791 (
            .O(N__35012),
            .I(N__35006));
    Odrv4 I__3790 (
            .O(N__35009),
            .I(\pid_alt.error_p_regZ0Z_9 ));
    Odrv4 I__3789 (
            .O(N__35006),
            .I(\pid_alt.error_p_regZ0Z_9 ));
    InMux I__3788 (
            .O(N__35001),
            .I(N__34998));
    LocalMux I__3787 (
            .O(N__34998),
            .I(N__34994));
    InMux I__3786 (
            .O(N__34997),
            .I(N__34991));
    Odrv4 I__3785 (
            .O(N__34994),
            .I(\pid_alt.error_d_reg_prevZ0Z_9 ));
    LocalMux I__3784 (
            .O(N__34991),
            .I(\pid_alt.error_d_reg_prevZ0Z_9 ));
    InMux I__3783 (
            .O(N__34986),
            .I(N__34983));
    LocalMux I__3782 (
            .O(N__34983),
            .I(N__34978));
    InMux I__3781 (
            .O(N__34982),
            .I(N__34973));
    InMux I__3780 (
            .O(N__34981),
            .I(N__34973));
    Span12Mux_h I__3779 (
            .O(N__34978),
            .I(N__34968));
    LocalMux I__3778 (
            .O(N__34973),
            .I(N__34968));
    Span12Mux_v I__3777 (
            .O(N__34968),
            .I(N__34965));
    Odrv12 I__3776 (
            .O(N__34965),
            .I(\pid_alt.error_d_regZ0Z_9 ));
    CascadeMux I__3775 (
            .O(N__34962),
            .I(N__34959));
    InMux I__3774 (
            .O(N__34959),
            .I(N__34955));
    InMux I__3773 (
            .O(N__34958),
            .I(N__34952));
    LocalMux I__3772 (
            .O(N__34955),
            .I(N__34949));
    LocalMux I__3771 (
            .O(N__34952),
            .I(N__34946));
    Span4Mux_h I__3770 (
            .O(N__34949),
            .I(N__34943));
    Odrv12 I__3769 (
            .O(N__34946),
            .I(\pid_alt.error_d_reg_prev_esr_RNIG75T2Z0Z_8 ));
    Odrv4 I__3768 (
            .O(N__34943),
            .I(\pid_alt.error_d_reg_prev_esr_RNIG75T2Z0Z_8 ));
    CascadeMux I__3767 (
            .O(N__34938),
            .I(\pid_alt.error_d_reg_prev_esr_RNIL8611Z0Z_9_cascade_ ));
    InMux I__3766 (
            .O(N__34935),
            .I(N__34932));
    LocalMux I__3765 (
            .O(N__34932),
            .I(N__34929));
    Odrv12 I__3764 (
            .O(N__34929),
            .I(\pid_alt.error_d_reg_prev_esr_RNICI045Z0Z_9 ));
    InMux I__3763 (
            .O(N__34926),
            .I(N__34923));
    LocalMux I__3762 (
            .O(N__34923),
            .I(\pid_alt.error_d_reg_prev_esr_RNIL8611Z0Z_9 ));
    InMux I__3761 (
            .O(N__34920),
            .I(N__34914));
    InMux I__3760 (
            .O(N__34919),
            .I(N__34914));
    LocalMux I__3759 (
            .O(N__34914),
            .I(N__34911));
    Span4Mux_v I__3758 (
            .O(N__34911),
            .I(N__34908));
    Odrv4 I__3757 (
            .O(N__34908),
            .I(\pid_alt.error_d_reg_prev_esr_RNIDAHM_0Z0Z_10 ));
    InMux I__3756 (
            .O(N__34905),
            .I(N__34902));
    LocalMux I__3755 (
            .O(N__34902),
            .I(N__34898));
    CascadeMux I__3754 (
            .O(N__34901),
            .I(N__34895));
    Span4Mux_h I__3753 (
            .O(N__34898),
            .I(N__34892));
    InMux I__3752 (
            .O(N__34895),
            .I(N__34889));
    Span4Mux_v I__3751 (
            .O(N__34892),
            .I(N__34886));
    LocalMux I__3750 (
            .O(N__34889),
            .I(N__34883));
    Odrv4 I__3749 (
            .O(N__34886),
            .I(\pid_alt.error_d_reg_prev_esr_RNISAR62Z0Z_9 ));
    Odrv12 I__3748 (
            .O(N__34883),
            .I(\pid_alt.error_d_reg_prev_esr_RNISAR62Z0Z_9 ));
    CascadeMux I__3747 (
            .O(N__34878),
            .I(N__34874));
    InMux I__3746 (
            .O(N__34877),
            .I(N__34871));
    InMux I__3745 (
            .O(N__34874),
            .I(N__34868));
    LocalMux I__3744 (
            .O(N__34871),
            .I(N__34865));
    LocalMux I__3743 (
            .O(N__34868),
            .I(N__34862));
    Span4Mux_v I__3742 (
            .O(N__34865),
            .I(N__34859));
    Span4Mux_h I__3741 (
            .O(N__34862),
            .I(N__34856));
    Odrv4 I__3740 (
            .O(N__34859),
            .I(\pid_alt.error_d_reg_prev_esr_RNI8BR02Z0Z_16 ));
    Odrv4 I__3739 (
            .O(N__34856),
            .I(\pid_alt.error_d_reg_prev_esr_RNI8BR02Z0Z_16 ));
    InMux I__3738 (
            .O(N__34851),
            .I(N__34848));
    LocalMux I__3737 (
            .O(N__34848),
            .I(\pid_alt.error_d_reg_prev_esr_RNIVSHMZ0Z_16 ));
    InMux I__3736 (
            .O(N__34845),
            .I(N__34839));
    InMux I__3735 (
            .O(N__34844),
            .I(N__34839));
    LocalMux I__3734 (
            .O(N__34839),
            .I(\pid_alt.error_d_reg_prev_esr_RNI20IM_0Z0Z_17 ));
    InMux I__3733 (
            .O(N__34836),
            .I(N__34833));
    LocalMux I__3732 (
            .O(N__34833),
            .I(N__34830));
    Odrv12 I__3731 (
            .O(N__34830),
            .I(\pid_alt.error_d_reg_prev_esr_RNICG9B1_0Z0Z_20 ));
    InMux I__3730 (
            .O(N__34827),
            .I(N__34824));
    LocalMux I__3729 (
            .O(N__34824),
            .I(N__34821));
    Span4Mux_h I__3728 (
            .O(N__34821),
            .I(N__34817));
    InMux I__3727 (
            .O(N__34820),
            .I(N__34814));
    Span4Mux_v I__3726 (
            .O(N__34817),
            .I(N__34811));
    LocalMux I__3725 (
            .O(N__34814),
            .I(N__34808));
    Odrv4 I__3724 (
            .O(N__34811),
            .I(\pid_alt.error_p_regZ0Z_19 ));
    Odrv12 I__3723 (
            .O(N__34808),
            .I(\pid_alt.error_p_regZ0Z_19 ));
    CascadeMux I__3722 (
            .O(N__34803),
            .I(N__34799));
    InMux I__3721 (
            .O(N__34802),
            .I(N__34796));
    InMux I__3720 (
            .O(N__34799),
            .I(N__34793));
    LocalMux I__3719 (
            .O(N__34796),
            .I(N__34788));
    LocalMux I__3718 (
            .O(N__34793),
            .I(N__34788));
    Span4Mux_v I__3717 (
            .O(N__34788),
            .I(N__34785));
    Odrv4 I__3716 (
            .O(N__34785),
            .I(\pid_alt.error_d_reg_prev_esr_RNIOTT02Z0Z_18 ));
    CascadeMux I__3715 (
            .O(N__34782),
            .I(\pid_alt.error_d_reg_prev_esr_RNI86IMZ0Z_19_cascade_ ));
    InMux I__3714 (
            .O(N__34779),
            .I(N__34776));
    LocalMux I__3713 (
            .O(N__34776),
            .I(N__34773));
    Odrv4 I__3712 (
            .O(N__34773),
            .I(\pid_alt.error_d_reg_prev_esr_RNIK3024Z0Z_19 ));
    InMux I__3711 (
            .O(N__34770),
            .I(N__34767));
    LocalMux I__3710 (
            .O(N__34767),
            .I(\pid_alt.un1_pid_prereg_236_1 ));
    InMux I__3709 (
            .O(N__34764),
            .I(N__34761));
    LocalMux I__3708 (
            .O(N__34761),
            .I(\pid_alt.error_d_reg_prev_esr_RNI86IMZ0Z_19 ));
    CascadeMux I__3707 (
            .O(N__34758),
            .I(\pid_alt.un1_pid_prereg_236_1_cascade_ ));
    InMux I__3706 (
            .O(N__34755),
            .I(N__34750));
    InMux I__3705 (
            .O(N__34754),
            .I(N__34745));
    InMux I__3704 (
            .O(N__34753),
            .I(N__34745));
    LocalMux I__3703 (
            .O(N__34750),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_19_c_RNI4FRJ ));
    LocalMux I__3702 (
            .O(N__34745),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_19_c_RNI4FRJ ));
    CascadeMux I__3701 (
            .O(N__34740),
            .I(N__34737));
    InMux I__3700 (
            .O(N__34737),
            .I(N__34734));
    LocalMux I__3699 (
            .O(N__34734),
            .I(N__34731));
    Odrv4 I__3698 (
            .O(N__34731),
            .I(\pid_alt.error_d_reg_prev_esr_RNIS5212Z0Z_19 ));
    InMux I__3697 (
            .O(N__34728),
            .I(N__34722));
    InMux I__3696 (
            .O(N__34727),
            .I(N__34722));
    LocalMux I__3695 (
            .O(N__34722),
            .I(N__34718));
    InMux I__3694 (
            .O(N__34721),
            .I(N__34715));
    Span4Mux_v I__3693 (
            .O(N__34718),
            .I(N__34712));
    LocalMux I__3692 (
            .O(N__34715),
            .I(N__34709));
    Sp12to4 I__3691 (
            .O(N__34712),
            .I(N__34706));
    Span4Mux_v I__3690 (
            .O(N__34709),
            .I(N__34703));
    Span12Mux_h I__3689 (
            .O(N__34706),
            .I(N__34698));
    Sp12to4 I__3688 (
            .O(N__34703),
            .I(N__34698));
    Odrv12 I__3687 (
            .O(N__34698),
            .I(\pid_alt.error_d_regZ0Z_19 ));
    InMux I__3686 (
            .O(N__34695),
            .I(N__34691));
    InMux I__3685 (
            .O(N__34694),
            .I(N__34688));
    LocalMux I__3684 (
            .O(N__34691),
            .I(N__34685));
    LocalMux I__3683 (
            .O(N__34688),
            .I(\pid_alt.error_d_reg_prevZ0Z_19 ));
    Odrv12 I__3682 (
            .O(N__34685),
            .I(\pid_alt.error_d_reg_prevZ0Z_19 ));
    CascadeMux I__3681 (
            .O(N__34680),
            .I(N__34677));
    InMux I__3680 (
            .O(N__34677),
            .I(N__34674));
    LocalMux I__3679 (
            .O(N__34674),
            .I(N__34671));
    Odrv4 I__3678 (
            .O(N__34671),
            .I(\pid_alt.error_d_reg_prev_esr_RNICG9B1_1Z0Z_20 ));
    InMux I__3677 (
            .O(N__34668),
            .I(N__34664));
    InMux I__3676 (
            .O(N__34667),
            .I(N__34661));
    LocalMux I__3675 (
            .O(N__34664),
            .I(N__34656));
    LocalMux I__3674 (
            .O(N__34661),
            .I(N__34656));
    Odrv4 I__3673 (
            .O(N__34656),
            .I(\pid_alt.error_d_reg_prev_esr_RNICG9B1Z0Z_20 ));
    InMux I__3672 (
            .O(N__34653),
            .I(N__34650));
    LocalMux I__3671 (
            .O(N__34650),
            .I(N__34647));
    Span4Mux_h I__3670 (
            .O(N__34647),
            .I(N__34644));
    Odrv4 I__3669 (
            .O(N__34644),
            .I(\pid_alt.error_d_reg_prev_esr_RNIOVN14Z0Z_17 ));
    InMux I__3668 (
            .O(N__34641),
            .I(N__34638));
    LocalMux I__3667 (
            .O(N__34638),
            .I(N__34635));
    Odrv4 I__3666 (
            .O(N__34635),
            .I(\pid_alt.pid_preregZ0Z_18 ));
    InMux I__3665 (
            .O(N__34632),
            .I(\pid_alt.un1_pid_prereg_0_cry_17 ));
    InMux I__3664 (
            .O(N__34629),
            .I(N__34626));
    LocalMux I__3663 (
            .O(N__34626),
            .I(N__34623));
    Span4Mux_h I__3662 (
            .O(N__34623),
            .I(N__34620));
    Odrv4 I__3661 (
            .O(N__34620),
            .I(\pid_alt.error_d_reg_prev_esr_RNI8IQ14Z0Z_18 ));
    CascadeMux I__3660 (
            .O(N__34617),
            .I(N__34614));
    InMux I__3659 (
            .O(N__34614),
            .I(N__34611));
    LocalMux I__3658 (
            .O(N__34611),
            .I(N__34607));
    InMux I__3657 (
            .O(N__34610),
            .I(N__34604));
    Span4Mux_h I__3656 (
            .O(N__34607),
            .I(N__34601));
    LocalMux I__3655 (
            .O(N__34604),
            .I(\pid_alt.error_d_reg_prev_esr_RNIGKS02Z0Z_17 ));
    Odrv4 I__3654 (
            .O(N__34601),
            .I(\pid_alt.error_d_reg_prev_esr_RNIGKS02Z0Z_17 ));
    InMux I__3653 (
            .O(N__34596),
            .I(N__34593));
    LocalMux I__3652 (
            .O(N__34593),
            .I(N__34590));
    Odrv4 I__3651 (
            .O(N__34590),
            .I(\pid_alt.pid_preregZ0Z_19 ));
    InMux I__3650 (
            .O(N__34587),
            .I(\pid_alt.un1_pid_prereg_0_cry_18 ));
    InMux I__3649 (
            .O(N__34584),
            .I(N__34581));
    LocalMux I__3648 (
            .O(N__34581),
            .I(N__34578));
    Odrv4 I__3647 (
            .O(N__34578),
            .I(\pid_alt.pid_preregZ0Z_20 ));
    InMux I__3646 (
            .O(N__34575),
            .I(\pid_alt.un1_pid_prereg_0_cry_19 ));
    CascadeMux I__3645 (
            .O(N__34572),
            .I(N__34569));
    InMux I__3644 (
            .O(N__34569),
            .I(N__34566));
    LocalMux I__3643 (
            .O(N__34566),
            .I(N__34563));
    Odrv12 I__3642 (
            .O(N__34563),
            .I(\pid_alt.pid_preregZ0Z_21 ));
    InMux I__3641 (
            .O(N__34560),
            .I(\pid_alt.un1_pid_prereg_0_cry_20 ));
    CascadeMux I__3640 (
            .O(N__34557),
            .I(N__34554));
    InMux I__3639 (
            .O(N__34554),
            .I(N__34551));
    LocalMux I__3638 (
            .O(N__34551),
            .I(N__34548));
    Span4Mux_h I__3637 (
            .O(N__34548),
            .I(N__34545));
    Odrv4 I__3636 (
            .O(N__34545),
            .I(\pid_alt.pid_preregZ0Z_22 ));
    InMux I__3635 (
            .O(N__34542),
            .I(\pid_alt.un1_pid_prereg_0_cry_21 ));
    InMux I__3634 (
            .O(N__34539),
            .I(N__34536));
    LocalMux I__3633 (
            .O(N__34536),
            .I(N__34533));
    Odrv12 I__3632 (
            .O(N__34533),
            .I(\pid_alt.pid_preregZ0Z_23 ));
    InMux I__3631 (
            .O(N__34530),
            .I(bfn_3_18_0_));
    InMux I__3630 (
            .O(N__34527),
            .I(N__34524));
    LocalMux I__3629 (
            .O(N__34524),
            .I(N__34521));
    Span4Mux_h I__3628 (
            .O(N__34521),
            .I(N__34518));
    Odrv4 I__3627 (
            .O(N__34518),
            .I(\pid_alt.un1_pid_prereg_0_axb_24 ));
    InMux I__3626 (
            .O(N__34515),
            .I(\pid_alt.un1_pid_prereg_0_cry_23 ));
    InMux I__3625 (
            .O(N__34512),
            .I(N__34507));
    InMux I__3624 (
            .O(N__34511),
            .I(N__34502));
    InMux I__3623 (
            .O(N__34510),
            .I(N__34502));
    LocalMux I__3622 (
            .O(N__34507),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_6_c_RNI3HMQ ));
    LocalMux I__3621 (
            .O(N__34502),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_6_c_RNI3HMQ ));
    InMux I__3620 (
            .O(N__34497),
            .I(N__34493));
    CascadeMux I__3619 (
            .O(N__34496),
            .I(N__34490));
    LocalMux I__3618 (
            .O(N__34493),
            .I(N__34487));
    InMux I__3617 (
            .O(N__34490),
            .I(N__34484));
    Span4Mux_v I__3616 (
            .O(N__34487),
            .I(N__34481));
    LocalMux I__3615 (
            .O(N__34484),
            .I(N__34478));
    Odrv4 I__3614 (
            .O(N__34481),
            .I(\pid_alt.error_d_reg_prev_esr_RNI7T3T2Z0Z_7 ));
    Odrv4 I__3613 (
            .O(N__34478),
            .I(\pid_alt.error_d_reg_prev_esr_RNI7T3T2Z0Z_7 ));
    InMux I__3612 (
            .O(N__34473),
            .I(\pid_alt.un1_pid_prereg_0_cry_8 ));
    InMux I__3611 (
            .O(N__34470),
            .I(\pid_alt.un1_pid_prereg_0_cry_9 ));
    InMux I__3610 (
            .O(N__34467),
            .I(N__34464));
    LocalMux I__3609 (
            .O(N__34464),
            .I(N__34461));
    Odrv4 I__3608 (
            .O(N__34461),
            .I(\pid_alt.error_d_reg_prev_esr_RNITPKD4Z0Z_10 ));
    InMux I__3607 (
            .O(N__34458),
            .I(\pid_alt.un1_pid_prereg_0_cry_10 ));
    InMux I__3606 (
            .O(N__34455),
            .I(\pid_alt.un1_pid_prereg_0_cry_11 ));
    InMux I__3605 (
            .O(N__34452),
            .I(\pid_alt.un1_pid_prereg_0_cry_12 ));
    InMux I__3604 (
            .O(N__34449),
            .I(N__34446));
    LocalMux I__3603 (
            .O(N__34446),
            .I(N__34443));
    Odrv4 I__3602 (
            .O(N__34443),
            .I(\pid_alt.pid_preregZ0Z_14 ));
    InMux I__3601 (
            .O(N__34440),
            .I(\pid_alt.un1_pid_prereg_0_cry_13 ));
    InMux I__3600 (
            .O(N__34437),
            .I(N__34434));
    LocalMux I__3599 (
            .O(N__34434),
            .I(N__34431));
    Odrv4 I__3598 (
            .O(N__34431),
            .I(\pid_alt.pid_preregZ0Z_15 ));
    InMux I__3597 (
            .O(N__34428),
            .I(bfn_3_17_0_));
    InMux I__3596 (
            .O(N__34425),
            .I(N__34422));
    LocalMux I__3595 (
            .O(N__34422),
            .I(N__34419));
    Odrv4 I__3594 (
            .O(N__34419),
            .I(\pid_alt.pid_preregZ0Z_16 ));
    InMux I__3593 (
            .O(N__34416),
            .I(\pid_alt.un1_pid_prereg_0_cry_15 ));
    InMux I__3592 (
            .O(N__34413),
            .I(N__34410));
    LocalMux I__3591 (
            .O(N__34410),
            .I(N__34407));
    Odrv4 I__3590 (
            .O(N__34407),
            .I(\pid_alt.pid_preregZ0Z_17 ));
    InMux I__3589 (
            .O(N__34404),
            .I(\pid_alt.un1_pid_prereg_0_cry_16 ));
    CascadeMux I__3588 (
            .O(N__34401),
            .I(N__34398));
    InMux I__3587 (
            .O(N__34398),
            .I(N__34395));
    LocalMux I__3586 (
            .O(N__34395),
            .I(\pid_alt.error_d_reg_prev_esr_RNIFPN33Z0Z_1 ));
    InMux I__3585 (
            .O(N__34392),
            .I(\pid_alt.un1_pid_prereg_0_cry_0 ));
    InMux I__3584 (
            .O(N__34389),
            .I(N__34386));
    LocalMux I__3583 (
            .O(N__34386),
            .I(\pid_alt.error_d_reg_prev_esr_RNIF0465Z0Z_1 ));
    InMux I__3582 (
            .O(N__34383),
            .I(\pid_alt.un1_pid_prereg_0_cry_1 ));
    InMux I__3581 (
            .O(N__34380),
            .I(N__34377));
    LocalMux I__3580 (
            .O(N__34377),
            .I(\pid_alt.error_d_reg_prev_esr_RNILDG87Z0Z_2 ));
    InMux I__3579 (
            .O(N__34374),
            .I(\pid_alt.un1_pid_prereg_0_cry_2 ));
    CascadeMux I__3578 (
            .O(N__34371),
            .I(N__34368));
    InMux I__3577 (
            .O(N__34368),
            .I(N__34364));
    InMux I__3576 (
            .O(N__34367),
            .I(N__34361));
    LocalMux I__3575 (
            .O(N__34364),
            .I(\pid_alt.error_d_reg_prev_esr_RNILE0V5Z0Z_2 ));
    LocalMux I__3574 (
            .O(N__34361),
            .I(\pid_alt.error_d_reg_prev_esr_RNILE0V5Z0Z_2 ));
    CascadeMux I__3573 (
            .O(N__34356),
            .I(N__34353));
    InMux I__3572 (
            .O(N__34353),
            .I(N__34350));
    LocalMux I__3571 (
            .O(N__34350),
            .I(\pid_alt.error_d_reg_prev_esr_RNI11TA9Z0Z_3 ));
    InMux I__3570 (
            .O(N__34347),
            .I(\pid_alt.un1_pid_prereg_0_cry_3 ));
    InMux I__3569 (
            .O(N__34344),
            .I(\pid_alt.un1_pid_prereg_0_cry_4 ));
    InMux I__3568 (
            .O(N__34341),
            .I(\pid_alt.un1_pid_prereg_0_cry_5 ));
    CascadeMux I__3567 (
            .O(N__34338),
            .I(N__34335));
    InMux I__3566 (
            .O(N__34335),
            .I(N__34332));
    LocalMux I__3565 (
            .O(N__34332),
            .I(\pid_alt.error_d_reg_prev_esr_RNIJR3Q5Z0Z_6 ));
    InMux I__3564 (
            .O(N__34329),
            .I(bfn_3_16_0_));
    InMux I__3563 (
            .O(N__34326),
            .I(N__34323));
    LocalMux I__3562 (
            .O(N__34323),
            .I(\pid_alt.error_d_reg_prev_esr_RNI5G6Q5Z0Z_7 ));
    CascadeMux I__3561 (
            .O(N__34320),
            .I(N__34316));
    InMux I__3560 (
            .O(N__34319),
            .I(N__34313));
    InMux I__3559 (
            .O(N__34316),
            .I(N__34310));
    LocalMux I__3558 (
            .O(N__34313),
            .I(\pid_alt.error_d_reg_prev_esr_RNIUI2T2Z0Z_6 ));
    LocalMux I__3557 (
            .O(N__34310),
            .I(\pid_alt.error_d_reg_prev_esr_RNIUI2T2Z0Z_6 ));
    InMux I__3556 (
            .O(N__34305),
            .I(\pid_alt.un1_pid_prereg_0_cry_7 ));
    InMux I__3555 (
            .O(N__34302),
            .I(N__34299));
    LocalMux I__3554 (
            .O(N__34299),
            .I(N__34296));
    Span4Mux_h I__3553 (
            .O(N__34296),
            .I(N__34293));
    Odrv4 I__3552 (
            .O(N__34293),
            .I(\pid_alt.error_d_reg_prev_esr_RNIN49Q5Z0Z_8 ));
    CascadeMux I__3551 (
            .O(N__34290),
            .I(\pid_alt.source_pid_1_sqmuxa_0_a2_2_5_cascade_ ));
    CascadeMux I__3550 (
            .O(N__34287),
            .I(\pid_alt.N_539_cascade_ ));
    CascadeMux I__3549 (
            .O(N__34284),
            .I(\pid_alt.source_pid_9_0_0_4_cascade_ ));
    InMux I__3548 (
            .O(N__34281),
            .I(N__34278));
    LocalMux I__3547 (
            .O(N__34278),
            .I(\pid_alt.source_pid_1_sqmuxa_0_a2_2_6 ));
    CascadeMux I__3546 (
            .O(N__34275),
            .I(N__34272));
    InMux I__3545 (
            .O(N__34272),
            .I(N__34269));
    LocalMux I__3544 (
            .O(N__34269),
            .I(N__34266));
    Span4Mux_v I__3543 (
            .O(N__34266),
            .I(N__34262));
    InMux I__3542 (
            .O(N__34265),
            .I(N__34259));
    Span4Mux_s3_h I__3541 (
            .O(N__34262),
            .I(N__34254));
    LocalMux I__3540 (
            .O(N__34259),
            .I(N__34254));
    Odrv4 I__3539 (
            .O(N__34254),
            .I(\pid_alt.error_d_reg_prev_i_0 ));
    InMux I__3538 (
            .O(N__34251),
            .I(N__34248));
    LocalMux I__3537 (
            .O(N__34248),
            .I(\pid_alt.error_p_reg_esr_RNI3SMI1Z0Z_0 ));
    CascadeMux I__3536 (
            .O(N__34245),
            .I(N__34242));
    InMux I__3535 (
            .O(N__34242),
            .I(N__34239));
    LocalMux I__3534 (
            .O(N__34239),
            .I(N__34235));
    InMux I__3533 (
            .O(N__34238),
            .I(N__34232));
    Span4Mux_v I__3532 (
            .O(N__34235),
            .I(N__34229));
    LocalMux I__3531 (
            .O(N__34232),
            .I(N__34226));
    Span4Mux_h I__3530 (
            .O(N__34229),
            .I(N__34223));
    Odrv12 I__3529 (
            .O(N__34226),
            .I(\pid_alt.un1_pid_prereg_0 ));
    Odrv4 I__3528 (
            .O(N__34223),
            .I(\pid_alt.un1_pid_prereg_0 ));
    InMux I__3527 (
            .O(N__34218),
            .I(\pid_alt.un1_pid_prereg_un1_pid_prereg_0_cry_0_c_THRU_CO ));
    CascadeMux I__3526 (
            .O(N__34215),
            .I(N__34211));
    InMux I__3525 (
            .O(N__34214),
            .I(N__34207));
    InMux I__3524 (
            .O(N__34211),
            .I(N__34202));
    InMux I__3523 (
            .O(N__34210),
            .I(N__34202));
    LocalMux I__3522 (
            .O(N__34207),
            .I(\Commands_frame_decoder.stateZ0Z_13 ));
    LocalMux I__3521 (
            .O(N__34202),
            .I(\Commands_frame_decoder.stateZ0Z_13 ));
    InMux I__3520 (
            .O(N__34197),
            .I(N__34191));
    InMux I__3519 (
            .O(N__34196),
            .I(N__34191));
    LocalMux I__3518 (
            .O(N__34191),
            .I(\Commands_frame_decoder.N_410 ));
    CascadeMux I__3517 (
            .O(N__34188),
            .I(N__34185));
    InMux I__3516 (
            .O(N__34185),
            .I(N__34181));
    InMux I__3515 (
            .O(N__34184),
            .I(N__34178));
    LocalMux I__3514 (
            .O(N__34181),
            .I(\Commands_frame_decoder.N_406 ));
    LocalMux I__3513 (
            .O(N__34178),
            .I(\Commands_frame_decoder.N_406 ));
    InMux I__3512 (
            .O(N__34173),
            .I(N__34170));
    LocalMux I__3511 (
            .O(N__34170),
            .I(N__34167));
    Odrv4 I__3510 (
            .O(N__34167),
            .I(\Commands_frame_decoder.WDT8lt14_0 ));
    InMux I__3509 (
            .O(N__34164),
            .I(N__34160));
    InMux I__3508 (
            .O(N__34163),
            .I(N__34154));
    LocalMux I__3507 (
            .O(N__34160),
            .I(N__34151));
    InMux I__3506 (
            .O(N__34159),
            .I(N__34148));
    InMux I__3505 (
            .O(N__34158),
            .I(N__34143));
    InMux I__3504 (
            .O(N__34157),
            .I(N__34143));
    LocalMux I__3503 (
            .O(N__34154),
            .I(\Commands_frame_decoder.WDTZ0Z_14 ));
    Odrv4 I__3502 (
            .O(N__34151),
            .I(\Commands_frame_decoder.WDTZ0Z_14 ));
    LocalMux I__3501 (
            .O(N__34148),
            .I(\Commands_frame_decoder.WDTZ0Z_14 ));
    LocalMux I__3500 (
            .O(N__34143),
            .I(\Commands_frame_decoder.WDTZ0Z_14 ));
    InMux I__3499 (
            .O(N__34134),
            .I(N__34130));
    InMux I__3498 (
            .O(N__34133),
            .I(N__34124));
    LocalMux I__3497 (
            .O(N__34130),
            .I(N__34121));
    InMux I__3496 (
            .O(N__34129),
            .I(N__34118));
    InMux I__3495 (
            .O(N__34128),
            .I(N__34113));
    InMux I__3494 (
            .O(N__34127),
            .I(N__34113));
    LocalMux I__3493 (
            .O(N__34124),
            .I(\Commands_frame_decoder.WDTZ0Z_15 ));
    Odrv4 I__3492 (
            .O(N__34121),
            .I(\Commands_frame_decoder.WDTZ0Z_15 ));
    LocalMux I__3491 (
            .O(N__34118),
            .I(\Commands_frame_decoder.WDTZ0Z_15 ));
    LocalMux I__3490 (
            .O(N__34113),
            .I(\Commands_frame_decoder.WDTZ0Z_15 ));
    CascadeMux I__3489 (
            .O(N__34104),
            .I(\Commands_frame_decoder.N_403_cascade_ ));
    CascadeMux I__3488 (
            .O(N__34101),
            .I(N__34097));
    InMux I__3487 (
            .O(N__34100),
            .I(N__34091));
    InMux I__3486 (
            .O(N__34097),
            .I(N__34091));
    InMux I__3485 (
            .O(N__34096),
            .I(N__34088));
    LocalMux I__3484 (
            .O(N__34091),
            .I(\Commands_frame_decoder.stateZ0Z_11 ));
    LocalMux I__3483 (
            .O(N__34088),
            .I(\Commands_frame_decoder.stateZ0Z_11 ));
    CascadeMux I__3482 (
            .O(N__34083),
            .I(N__34080));
    InMux I__3481 (
            .O(N__34080),
            .I(N__34074));
    InMux I__3480 (
            .O(N__34079),
            .I(N__34074));
    LocalMux I__3479 (
            .O(N__34074),
            .I(\Commands_frame_decoder.stateZ0Z_8 ));
    InMux I__3478 (
            .O(N__34071),
            .I(N__34067));
    InMux I__3477 (
            .O(N__34070),
            .I(N__34064));
    LocalMux I__3476 (
            .O(N__34067),
            .I(\Commands_frame_decoder.stateZ0Z_9 ));
    LocalMux I__3475 (
            .O(N__34064),
            .I(\Commands_frame_decoder.stateZ0Z_9 ));
    CascadeMux I__3474 (
            .O(N__34059),
            .I(N__34053));
    InMux I__3473 (
            .O(N__34058),
            .I(N__34050));
    InMux I__3472 (
            .O(N__34057),
            .I(N__34045));
    InMux I__3471 (
            .O(N__34056),
            .I(N__34045));
    InMux I__3470 (
            .O(N__34053),
            .I(N__34042));
    LocalMux I__3469 (
            .O(N__34050),
            .I(N__34039));
    LocalMux I__3468 (
            .O(N__34045),
            .I(\Commands_frame_decoder.stateZ0Z_7 ));
    LocalMux I__3467 (
            .O(N__34042),
            .I(\Commands_frame_decoder.stateZ0Z_7 ));
    Odrv12 I__3466 (
            .O(N__34039),
            .I(\Commands_frame_decoder.stateZ0Z_7 ));
    SRMux I__3465 (
            .O(N__34032),
            .I(N__34029));
    LocalMux I__3464 (
            .O(N__34029),
            .I(N__34026));
    Sp12to4 I__3463 (
            .O(N__34026),
            .I(N__34022));
    SRMux I__3462 (
            .O(N__34025),
            .I(N__34019));
    Odrv12 I__3461 (
            .O(N__34022),
            .I(\Commands_frame_decoder.un1_state57_iZ0 ));
    LocalMux I__3460 (
            .O(N__34019),
            .I(\Commands_frame_decoder.un1_state57_iZ0 ));
    CascadeMux I__3459 (
            .O(N__34014),
            .I(N__34011));
    InMux I__3458 (
            .O(N__34011),
            .I(N__34002));
    InMux I__3457 (
            .O(N__34010),
            .I(N__34002));
    InMux I__3456 (
            .O(N__34009),
            .I(N__34002));
    LocalMux I__3455 (
            .O(N__34002),
            .I(\Commands_frame_decoder.countZ0Z_0 ));
    InMux I__3454 (
            .O(N__33999),
            .I(N__33996));
    LocalMux I__3453 (
            .O(N__33996),
            .I(\Commands_frame_decoder.N_370_2 ));
    InMux I__3452 (
            .O(N__33993),
            .I(N__33990));
    LocalMux I__3451 (
            .O(N__33990),
            .I(\Commands_frame_decoder.N_371 ));
    CascadeMux I__3450 (
            .O(N__33987),
            .I(\Commands_frame_decoder.N_370_2_cascade_ ));
    InMux I__3449 (
            .O(N__33984),
            .I(N__33981));
    LocalMux I__3448 (
            .O(N__33981),
            .I(N__33977));
    InMux I__3447 (
            .O(N__33980),
            .I(N__33974));
    Odrv4 I__3446 (
            .O(N__33977),
            .I(\Commands_frame_decoder.N_365_0 ));
    LocalMux I__3445 (
            .O(N__33974),
            .I(\Commands_frame_decoder.N_365_0 ));
    CascadeMux I__3444 (
            .O(N__33969),
            .I(\Commands_frame_decoder.state_ns_i_0_0_cascade_ ));
    InMux I__3443 (
            .O(N__33966),
            .I(N__33962));
    InMux I__3442 (
            .O(N__33965),
            .I(N__33959));
    LocalMux I__3441 (
            .O(N__33962),
            .I(\Commands_frame_decoder.stateZ0Z_0 ));
    LocalMux I__3440 (
            .O(N__33959),
            .I(\Commands_frame_decoder.stateZ0Z_0 ));
    CascadeMux I__3439 (
            .O(N__33954),
            .I(N__33951));
    InMux I__3438 (
            .O(N__33951),
            .I(N__33948));
    LocalMux I__3437 (
            .O(N__33948),
            .I(N__33945));
    Odrv4 I__3436 (
            .O(N__33945),
            .I(\Commands_frame_decoder.state_ns_0_a3_3_1 ));
    InMux I__3435 (
            .O(N__33942),
            .I(N__33936));
    InMux I__3434 (
            .O(N__33941),
            .I(N__33929));
    InMux I__3433 (
            .O(N__33940),
            .I(N__33929));
    InMux I__3432 (
            .O(N__33939),
            .I(N__33929));
    LocalMux I__3431 (
            .O(N__33936),
            .I(\Commands_frame_decoder.stateZ0Z_1 ));
    LocalMux I__3430 (
            .O(N__33929),
            .I(\Commands_frame_decoder.stateZ0Z_1 ));
    InMux I__3429 (
            .O(N__33924),
            .I(N__33918));
    InMux I__3428 (
            .O(N__33923),
            .I(N__33918));
    LocalMux I__3427 (
            .O(N__33918),
            .I(\Commands_frame_decoder.N_372 ));
    CascadeMux I__3426 (
            .O(N__33915),
            .I(N__33912));
    InMux I__3425 (
            .O(N__33912),
            .I(N__33906));
    InMux I__3424 (
            .O(N__33911),
            .I(N__33901));
    InMux I__3423 (
            .O(N__33910),
            .I(N__33901));
    InMux I__3422 (
            .O(N__33909),
            .I(N__33898));
    LocalMux I__3421 (
            .O(N__33906),
            .I(\Commands_frame_decoder.stateZ0Z_14 ));
    LocalMux I__3420 (
            .O(N__33901),
            .I(\Commands_frame_decoder.stateZ0Z_14 ));
    LocalMux I__3419 (
            .O(N__33898),
            .I(\Commands_frame_decoder.stateZ0Z_14 ));
    InMux I__3418 (
            .O(N__33891),
            .I(N__33886));
    InMux I__3417 (
            .O(N__33890),
            .I(N__33883));
    InMux I__3416 (
            .O(N__33889),
            .I(N__33880));
    LocalMux I__3415 (
            .O(N__33886),
            .I(\Commands_frame_decoder.WDTZ0Z_10 ));
    LocalMux I__3414 (
            .O(N__33883),
            .I(\Commands_frame_decoder.WDTZ0Z_10 ));
    LocalMux I__3413 (
            .O(N__33880),
            .I(\Commands_frame_decoder.WDTZ0Z_10 ));
    InMux I__3412 (
            .O(N__33873),
            .I(N__33867));
    InMux I__3411 (
            .O(N__33872),
            .I(N__33864));
    InMux I__3410 (
            .O(N__33871),
            .I(N__33859));
    InMux I__3409 (
            .O(N__33870),
            .I(N__33859));
    LocalMux I__3408 (
            .O(N__33867),
            .I(\Commands_frame_decoder.WDTZ0Z_13 ));
    LocalMux I__3407 (
            .O(N__33864),
            .I(\Commands_frame_decoder.WDTZ0Z_13 ));
    LocalMux I__3406 (
            .O(N__33859),
            .I(\Commands_frame_decoder.WDTZ0Z_13 ));
    CascadeMux I__3405 (
            .O(N__33852),
            .I(N__33848));
    InMux I__3404 (
            .O(N__33851),
            .I(N__33843));
    InMux I__3403 (
            .O(N__33848),
            .I(N__33838));
    InMux I__3402 (
            .O(N__33847),
            .I(N__33838));
    InMux I__3401 (
            .O(N__33846),
            .I(N__33835));
    LocalMux I__3400 (
            .O(N__33843),
            .I(\Commands_frame_decoder.WDTZ0Z_12 ));
    LocalMux I__3399 (
            .O(N__33838),
            .I(\Commands_frame_decoder.WDTZ0Z_12 ));
    LocalMux I__3398 (
            .O(N__33835),
            .I(\Commands_frame_decoder.WDTZ0Z_12 ));
    InMux I__3397 (
            .O(N__33828),
            .I(N__33822));
    InMux I__3396 (
            .O(N__33827),
            .I(N__33817));
    InMux I__3395 (
            .O(N__33826),
            .I(N__33817));
    InMux I__3394 (
            .O(N__33825),
            .I(N__33814));
    LocalMux I__3393 (
            .O(N__33822),
            .I(\Commands_frame_decoder.WDTZ0Z_11 ));
    LocalMux I__3392 (
            .O(N__33817),
            .I(\Commands_frame_decoder.WDTZ0Z_11 ));
    LocalMux I__3391 (
            .O(N__33814),
            .I(\Commands_frame_decoder.WDTZ0Z_11 ));
    InMux I__3390 (
            .O(N__33807),
            .I(N__33802));
    InMux I__3389 (
            .O(N__33806),
            .I(N__33799));
    InMux I__3388 (
            .O(N__33805),
            .I(N__33796));
    LocalMux I__3387 (
            .O(N__33802),
            .I(\Commands_frame_decoder.WDTZ0Z_6 ));
    LocalMux I__3386 (
            .O(N__33799),
            .I(\Commands_frame_decoder.WDTZ0Z_6 ));
    LocalMux I__3385 (
            .O(N__33796),
            .I(\Commands_frame_decoder.WDTZ0Z_6 ));
    InMux I__3384 (
            .O(N__33789),
            .I(N__33784));
    InMux I__3383 (
            .O(N__33788),
            .I(N__33781));
    InMux I__3382 (
            .O(N__33787),
            .I(N__33778));
    LocalMux I__3381 (
            .O(N__33784),
            .I(\Commands_frame_decoder.WDTZ0Z_5 ));
    LocalMux I__3380 (
            .O(N__33781),
            .I(\Commands_frame_decoder.WDTZ0Z_5 ));
    LocalMux I__3379 (
            .O(N__33778),
            .I(\Commands_frame_decoder.WDTZ0Z_5 ));
    CascadeMux I__3378 (
            .O(N__33771),
            .I(N__33766));
    CascadeMux I__3377 (
            .O(N__33770),
            .I(N__33763));
    InMux I__3376 (
            .O(N__33769),
            .I(N__33760));
    InMux I__3375 (
            .O(N__33766),
            .I(N__33757));
    InMux I__3374 (
            .O(N__33763),
            .I(N__33754));
    LocalMux I__3373 (
            .O(N__33760),
            .I(\Commands_frame_decoder.WDTZ0Z_7 ));
    LocalMux I__3372 (
            .O(N__33757),
            .I(\Commands_frame_decoder.WDTZ0Z_7 ));
    LocalMux I__3371 (
            .O(N__33754),
            .I(\Commands_frame_decoder.WDTZ0Z_7 ));
    InMux I__3370 (
            .O(N__33747),
            .I(N__33742));
    InMux I__3369 (
            .O(N__33746),
            .I(N__33739));
    InMux I__3368 (
            .O(N__33745),
            .I(N__33736));
    LocalMux I__3367 (
            .O(N__33742),
            .I(\Commands_frame_decoder.WDTZ0Z_4 ));
    LocalMux I__3366 (
            .O(N__33739),
            .I(\Commands_frame_decoder.WDTZ0Z_4 ));
    LocalMux I__3365 (
            .O(N__33736),
            .I(\Commands_frame_decoder.WDTZ0Z_4 ));
    InMux I__3364 (
            .O(N__33729),
            .I(N__33726));
    LocalMux I__3363 (
            .O(N__33726),
            .I(\Commands_frame_decoder.WDT_RNI2VDI1Z0Z_10 ));
    InMux I__3362 (
            .O(N__33723),
            .I(N__33720));
    LocalMux I__3361 (
            .O(N__33720),
            .I(\Commands_frame_decoder.WDT_RNITK4LZ0Z_8 ));
    CascadeMux I__3360 (
            .O(N__33717),
            .I(\Commands_frame_decoder.WDT_RNIET8A1Z0Z_4_cascade_ ));
    InMux I__3359 (
            .O(N__33714),
            .I(N__33711));
    LocalMux I__3358 (
            .O(N__33711),
            .I(\Commands_frame_decoder.WDT_RNIHV6PZ0Z_11 ));
    CascadeMux I__3357 (
            .O(N__33708),
            .I(\Commands_frame_decoder.WDT8lt14_0_cascade_ ));
    CEMux I__3356 (
            .O(N__33705),
            .I(N__33702));
    LocalMux I__3355 (
            .O(N__33702),
            .I(N__33699));
    Odrv4 I__3354 (
            .O(N__33699),
            .I(\Commands_frame_decoder.state_RNIQRI31Z0Z_10 ));
    InMux I__3353 (
            .O(N__33696),
            .I(N__33693));
    LocalMux I__3352 (
            .O(N__33693),
            .I(N__33690));
    Odrv12 I__3351 (
            .O(N__33690),
            .I(\Commands_frame_decoder.count_1_sqmuxa ));
    CascadeMux I__3350 (
            .O(N__33687),
            .I(\Commands_frame_decoder.WDT8lto9_3_cascade_ ));
    CascadeMux I__3349 (
            .O(N__33684),
            .I(N__33681));
    InMux I__3348 (
            .O(N__33681),
            .I(N__33678));
    LocalMux I__3347 (
            .O(N__33678),
            .I(\Commands_frame_decoder.state_0_sqmuxacf0_1 ));
    InMux I__3346 (
            .O(N__33675),
            .I(N__33672));
    LocalMux I__3345 (
            .O(N__33672),
            .I(\Commands_frame_decoder.state_0_sqmuxacf1 ));
    CascadeMux I__3344 (
            .O(N__33669),
            .I(\Commands_frame_decoder.state_0_sqmuxacf0_cascade_ ));
    InMux I__3343 (
            .O(N__33666),
            .I(N__33663));
    LocalMux I__3342 (
            .O(N__33663),
            .I(\Commands_frame_decoder.WDT8lt12_0 ));
    CascadeMux I__3341 (
            .O(N__33660),
            .I(N__33656));
    InMux I__3340 (
            .O(N__33659),
            .I(N__33653));
    InMux I__3339 (
            .O(N__33656),
            .I(N__33650));
    LocalMux I__3338 (
            .O(N__33653),
            .I(\Commands_frame_decoder.state_0_sqmuxa ));
    LocalMux I__3337 (
            .O(N__33650),
            .I(\Commands_frame_decoder.state_0_sqmuxa ));
    CascadeMux I__3336 (
            .O(N__33645),
            .I(N__33639));
    InMux I__3335 (
            .O(N__33644),
            .I(N__33630));
    InMux I__3334 (
            .O(N__33643),
            .I(N__33630));
    InMux I__3333 (
            .O(N__33642),
            .I(N__33630));
    InMux I__3332 (
            .O(N__33639),
            .I(N__33630));
    LocalMux I__3331 (
            .O(N__33630),
            .I(\Commands_frame_decoder.preinitZ0 ));
    InMux I__3330 (
            .O(N__33627),
            .I(N__33622));
    InMux I__3329 (
            .O(N__33626),
            .I(N__33619));
    InMux I__3328 (
            .O(N__33625),
            .I(N__33616));
    LocalMux I__3327 (
            .O(N__33622),
            .I(\Commands_frame_decoder.WDTZ0Z_8 ));
    LocalMux I__3326 (
            .O(N__33619),
            .I(\Commands_frame_decoder.WDTZ0Z_8 ));
    LocalMux I__3325 (
            .O(N__33616),
            .I(\Commands_frame_decoder.WDTZ0Z_8 ));
    InMux I__3324 (
            .O(N__33609),
            .I(N__33604));
    InMux I__3323 (
            .O(N__33608),
            .I(N__33601));
    InMux I__3322 (
            .O(N__33607),
            .I(N__33598));
    LocalMux I__3321 (
            .O(N__33604),
            .I(\Commands_frame_decoder.WDTZ0Z_9 ));
    LocalMux I__3320 (
            .O(N__33601),
            .I(\Commands_frame_decoder.WDTZ0Z_9 ));
    LocalMux I__3319 (
            .O(N__33598),
            .I(\Commands_frame_decoder.WDTZ0Z_9 ));
    CascadeMux I__3318 (
            .O(N__33591),
            .I(\pid_alt.N_545_cascade_ ));
    InMux I__3317 (
            .O(N__33588),
            .I(N__33585));
    LocalMux I__3316 (
            .O(N__33585),
            .I(\pid_alt.error_i_acumm_preregZ0Z_16 ));
    InMux I__3315 (
            .O(N__33582),
            .I(N__33579));
    LocalMux I__3314 (
            .O(N__33579),
            .I(N__33574));
    InMux I__3313 (
            .O(N__33578),
            .I(N__33569));
    InMux I__3312 (
            .O(N__33577),
            .I(N__33569));
    Odrv4 I__3311 (
            .O(N__33574),
            .I(\pid_alt.error_i_reg_esr_RNIBKPJZ0Z_19 ));
    LocalMux I__3310 (
            .O(N__33569),
            .I(\pid_alt.error_i_reg_esr_RNIBKPJZ0Z_19 ));
    InMux I__3309 (
            .O(N__33564),
            .I(N__33561));
    LocalMux I__3308 (
            .O(N__33561),
            .I(\pid_alt.error_i_acumm_preregZ0Z_19 ));
    InMux I__3307 (
            .O(N__33558),
            .I(N__33555));
    LocalMux I__3306 (
            .O(N__33555),
            .I(\pid_alt.error_i_acumm_preregZ0Z_14 ));
    InMux I__3305 (
            .O(N__33552),
            .I(N__33549));
    LocalMux I__3304 (
            .O(N__33549),
            .I(N__33546));
    Span4Mux_h I__3303 (
            .O(N__33546),
            .I(N__33543));
    Odrv4 I__3302 (
            .O(N__33543),
            .I(\pid_alt.O_5_12 ));
    InMux I__3301 (
            .O(N__33540),
            .I(N__33537));
    LocalMux I__3300 (
            .O(N__33537),
            .I(N__33533));
    InMux I__3299 (
            .O(N__33536),
            .I(N__33530));
    Span4Mux_s2_h I__3298 (
            .O(N__33533),
            .I(N__33527));
    LocalMux I__3297 (
            .O(N__33530),
            .I(N__33524));
    Odrv4 I__3296 (
            .O(N__33527),
            .I(\pid_alt.error_p_regZ0Z_8 ));
    Odrv12 I__3295 (
            .O(N__33524),
            .I(\pid_alt.error_p_regZ0Z_8 ));
    InMux I__3294 (
            .O(N__33519),
            .I(N__33516));
    LocalMux I__3293 (
            .O(N__33516),
            .I(N__33513));
    Odrv4 I__3292 (
            .O(N__33513),
            .I(\pid_alt.O_5_5 ));
    InMux I__3291 (
            .O(N__33510),
            .I(N__33501));
    InMux I__3290 (
            .O(N__33509),
            .I(N__33501));
    InMux I__3289 (
            .O(N__33508),
            .I(N__33501));
    LocalMux I__3288 (
            .O(N__33501),
            .I(N__33498));
    Sp12to4 I__3287 (
            .O(N__33498),
            .I(N__33495));
    Odrv12 I__3286 (
            .O(N__33495),
            .I(\pid_alt.error_p_regZ0Z_1 ));
    InMux I__3285 (
            .O(N__33492),
            .I(N__33489));
    LocalMux I__3284 (
            .O(N__33489),
            .I(N__33486));
    Odrv4 I__3283 (
            .O(N__33486),
            .I(\pid_alt.O_5_7 ));
    InMux I__3282 (
            .O(N__33483),
            .I(N__33477));
    InMux I__3281 (
            .O(N__33482),
            .I(N__33477));
    LocalMux I__3280 (
            .O(N__33477),
            .I(N__33474));
    Span12Mux_v I__3279 (
            .O(N__33474),
            .I(N__33471));
    Odrv12 I__3278 (
            .O(N__33471),
            .I(\pid_alt.error_p_regZ0Z_3 ));
    CEMux I__3277 (
            .O(N__33468),
            .I(N__33423));
    CEMux I__3276 (
            .O(N__33467),
            .I(N__33423));
    CEMux I__3275 (
            .O(N__33466),
            .I(N__33423));
    CEMux I__3274 (
            .O(N__33465),
            .I(N__33423));
    CEMux I__3273 (
            .O(N__33464),
            .I(N__33423));
    CEMux I__3272 (
            .O(N__33463),
            .I(N__33423));
    CEMux I__3271 (
            .O(N__33462),
            .I(N__33423));
    CEMux I__3270 (
            .O(N__33461),
            .I(N__33423));
    CEMux I__3269 (
            .O(N__33460),
            .I(N__33423));
    CEMux I__3268 (
            .O(N__33459),
            .I(N__33423));
    CEMux I__3267 (
            .O(N__33458),
            .I(N__33423));
    CEMux I__3266 (
            .O(N__33457),
            .I(N__33423));
    CEMux I__3265 (
            .O(N__33456),
            .I(N__33423));
    CEMux I__3264 (
            .O(N__33455),
            .I(N__33423));
    CEMux I__3263 (
            .O(N__33454),
            .I(N__33423));
    GlobalMux I__3262 (
            .O(N__33423),
            .I(N__33420));
    gio2CtrlBuf I__3261 (
            .O(N__33420),
            .I(\pid_alt.N_939_0_g ));
    InMux I__3260 (
            .O(N__33417),
            .I(N__33414));
    LocalMux I__3259 (
            .O(N__33414),
            .I(N__33411));
    Odrv12 I__3258 (
            .O(N__33411),
            .I(alt_kd_0));
    CEMux I__3257 (
            .O(N__33408),
            .I(N__33405));
    LocalMux I__3256 (
            .O(N__33405),
            .I(N__33400));
    CEMux I__3255 (
            .O(N__33404),
            .I(N__33397));
    CEMux I__3254 (
            .O(N__33403),
            .I(N__33394));
    Span4Mux_h I__3253 (
            .O(N__33400),
            .I(N__33389));
    LocalMux I__3252 (
            .O(N__33397),
            .I(N__33389));
    LocalMux I__3251 (
            .O(N__33394),
            .I(N__33386));
    Span4Mux_v I__3250 (
            .O(N__33389),
            .I(N__33381));
    Span4Mux_v I__3249 (
            .O(N__33386),
            .I(N__33381));
    Odrv4 I__3248 (
            .O(N__33381),
            .I(\Commands_frame_decoder.state_RNIRSI31Z0Z_11 ));
    CascadeMux I__3247 (
            .O(N__33378),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_20_c_RNISVKK_cascade_ ));
    InMux I__3246 (
            .O(N__33375),
            .I(N__33371));
    InMux I__3245 (
            .O(N__33374),
            .I(N__33368));
    LocalMux I__3244 (
            .O(N__33371),
            .I(\pid_alt.error_p_regZ0Z_17 ));
    LocalMux I__3243 (
            .O(N__33368),
            .I(\pid_alt.error_p_regZ0Z_17 ));
    InMux I__3242 (
            .O(N__33363),
            .I(N__33358));
    InMux I__3241 (
            .O(N__33362),
            .I(N__33353));
    InMux I__3240 (
            .O(N__33361),
            .I(N__33353));
    LocalMux I__3239 (
            .O(N__33358),
            .I(N__33350));
    LocalMux I__3238 (
            .O(N__33353),
            .I(N__33347));
    Odrv4 I__3237 (
            .O(N__33350),
            .I(\pid_alt.error_i_reg_esr_RNI4NMPZ0Z_11 ));
    Odrv4 I__3236 (
            .O(N__33347),
            .I(\pid_alt.error_i_reg_esr_RNI4NMPZ0Z_11 ));
    InMux I__3235 (
            .O(N__33342),
            .I(N__33337));
    InMux I__3234 (
            .O(N__33341),
            .I(N__33332));
    InMux I__3233 (
            .O(N__33340),
            .I(N__33332));
    LocalMux I__3232 (
            .O(N__33337),
            .I(\pid_alt.error_i_reg_esr_RNI9HOJZ0Z_18 ));
    LocalMux I__3231 (
            .O(N__33332),
            .I(\pid_alt.error_i_reg_esr_RNI9HOJZ0Z_18 ));
    InMux I__3230 (
            .O(N__33327),
            .I(N__33324));
    LocalMux I__3229 (
            .O(N__33324),
            .I(N__33320));
    InMux I__3228 (
            .O(N__33323),
            .I(N__33317));
    Span4Mux_v I__3227 (
            .O(N__33320),
            .I(N__33313));
    LocalMux I__3226 (
            .O(N__33317),
            .I(N__33310));
    InMux I__3225 (
            .O(N__33316),
            .I(N__33307));
    Span4Mux_v I__3224 (
            .O(N__33313),
            .I(N__33304));
    Span12Mux_h I__3223 (
            .O(N__33310),
            .I(N__33299));
    LocalMux I__3222 (
            .O(N__33307),
            .I(N__33299));
    Span4Mux_v I__3221 (
            .O(N__33304),
            .I(N__33296));
    Span12Mux_v I__3220 (
            .O(N__33299),
            .I(N__33293));
    Span4Mux_v I__3219 (
            .O(N__33296),
            .I(N__33290));
    Odrv12 I__3218 (
            .O(N__33293),
            .I(\pid_alt.error_d_regZ0Z_17 ));
    Odrv4 I__3217 (
            .O(N__33290),
            .I(\pid_alt.error_d_regZ0Z_17 ));
    InMux I__3216 (
            .O(N__33285),
            .I(N__33281));
    InMux I__3215 (
            .O(N__33284),
            .I(N__33278));
    LocalMux I__3214 (
            .O(N__33281),
            .I(\pid_alt.error_d_reg_prevZ0Z_17 ));
    LocalMux I__3213 (
            .O(N__33278),
            .I(\pid_alt.error_d_reg_prevZ0Z_17 ));
    InMux I__3212 (
            .O(N__33273),
            .I(N__33270));
    LocalMux I__3211 (
            .O(N__33270),
            .I(\pid_alt.error_i_acumm_preregZ0Z_18 ));
    CascadeMux I__3210 (
            .O(N__33267),
            .I(N__33264));
    InMux I__3209 (
            .O(N__33264),
            .I(N__33261));
    LocalMux I__3208 (
            .O(N__33261),
            .I(\pid_alt.error_i_acumm_preregZ0Z_20 ));
    InMux I__3207 (
            .O(N__33258),
            .I(N__33255));
    LocalMux I__3206 (
            .O(N__33255),
            .I(\pid_alt.error_i_acumm_preregZ0Z_17 ));
    CascadeMux I__3205 (
            .O(N__33252),
            .I(\pid_alt.m7_e_4_cascade_ ));
    InMux I__3204 (
            .O(N__33249),
            .I(N__33246));
    LocalMux I__3203 (
            .O(N__33246),
            .I(N__33243));
    Span4Mux_v I__3202 (
            .O(N__33243),
            .I(N__33240));
    Span4Mux_v I__3201 (
            .O(N__33240),
            .I(N__33237));
    Odrv4 I__3200 (
            .O(N__33237),
            .I(\pid_alt.error_i_regZ0Z_14 ));
    InMux I__3199 (
            .O(N__33234),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_13 ));
    InMux I__3198 (
            .O(N__33231),
            .I(N__33228));
    LocalMux I__3197 (
            .O(N__33228),
            .I(N__33225));
    Span4Mux_v I__3196 (
            .O(N__33225),
            .I(N__33222));
    Span4Mux_v I__3195 (
            .O(N__33222),
            .I(N__33219));
    Odrv4 I__3194 (
            .O(N__33219),
            .I(\pid_alt.error_i_regZ0Z_15 ));
    InMux I__3193 (
            .O(N__33216),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_14 ));
    InMux I__3192 (
            .O(N__33213),
            .I(N__33210));
    LocalMux I__3191 (
            .O(N__33210),
            .I(N__33207));
    Span4Mux_v I__3190 (
            .O(N__33207),
            .I(N__33204));
    Span4Mux_v I__3189 (
            .O(N__33204),
            .I(N__33201));
    Odrv4 I__3188 (
            .O(N__33201),
            .I(\pid_alt.error_i_regZ0Z_16 ));
    InMux I__3187 (
            .O(N__33198),
            .I(bfn_2_20_0_));
    InMux I__3186 (
            .O(N__33195),
            .I(N__33192));
    LocalMux I__3185 (
            .O(N__33192),
            .I(N__33189));
    Span4Mux_v I__3184 (
            .O(N__33189),
            .I(N__33186));
    Span4Mux_v I__3183 (
            .O(N__33186),
            .I(N__33183));
    Odrv4 I__3182 (
            .O(N__33183),
            .I(\pid_alt.error_i_regZ0Z_17 ));
    InMux I__3181 (
            .O(N__33180),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_16 ));
    InMux I__3180 (
            .O(N__33177),
            .I(N__33174));
    LocalMux I__3179 (
            .O(N__33174),
            .I(N__33171));
    Span4Mux_v I__3178 (
            .O(N__33171),
            .I(N__33168));
    Span4Mux_v I__3177 (
            .O(N__33168),
            .I(N__33165));
    Odrv4 I__3176 (
            .O(N__33165),
            .I(\pid_alt.error_i_regZ0Z_18 ));
    InMux I__3175 (
            .O(N__33162),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_17 ));
    InMux I__3174 (
            .O(N__33159),
            .I(N__33156));
    LocalMux I__3173 (
            .O(N__33156),
            .I(N__33153));
    Span4Mux_v I__3172 (
            .O(N__33153),
            .I(N__33150));
    Span4Mux_v I__3171 (
            .O(N__33150),
            .I(N__33147));
    Odrv4 I__3170 (
            .O(N__33147),
            .I(\pid_alt.error_i_regZ0Z_19 ));
    InMux I__3169 (
            .O(N__33144),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_18 ));
    InMux I__3168 (
            .O(N__33141),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_19 ));
    InMux I__3167 (
            .O(N__33138),
            .I(N__33132));
    InMux I__3166 (
            .O(N__33137),
            .I(N__33132));
    LocalMux I__3165 (
            .O(N__33132),
            .I(N__33129));
    Span12Mux_v I__3164 (
            .O(N__33129),
            .I(N__33126));
    Odrv12 I__3163 (
            .O(N__33126),
            .I(\pid_alt.error_i_regZ0Z_20 ));
    InMux I__3162 (
            .O(N__33123),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_20 ));
    CascadeMux I__3161 (
            .O(N__33120),
            .I(N__33117));
    InMux I__3160 (
            .O(N__33117),
            .I(N__33114));
    LocalMux I__3159 (
            .O(N__33114),
            .I(N__33111));
    Span4Mux_v I__3158 (
            .O(N__33111),
            .I(N__33108));
    Span4Mux_v I__3157 (
            .O(N__33108),
            .I(N__33105));
    Odrv4 I__3156 (
            .O(N__33105),
            .I(\pid_alt.error_i_regZ0Z_6 ));
    InMux I__3155 (
            .O(N__33102),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_5 ));
    CascadeMux I__3154 (
            .O(N__33099),
            .I(N__33096));
    InMux I__3153 (
            .O(N__33096),
            .I(N__33093));
    LocalMux I__3152 (
            .O(N__33093),
            .I(N__33090));
    Span4Mux_v I__3151 (
            .O(N__33090),
            .I(N__33087));
    Span4Mux_v I__3150 (
            .O(N__33087),
            .I(N__33084));
    Span4Mux_v I__3149 (
            .O(N__33084),
            .I(N__33081));
    Odrv4 I__3148 (
            .O(N__33081),
            .I(\pid_alt.error_i_regZ0Z_7 ));
    InMux I__3147 (
            .O(N__33078),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_6 ));
    CascadeMux I__3146 (
            .O(N__33075),
            .I(N__33072));
    InMux I__3145 (
            .O(N__33072),
            .I(N__33069));
    LocalMux I__3144 (
            .O(N__33069),
            .I(N__33066));
    Span4Mux_v I__3143 (
            .O(N__33066),
            .I(N__33063));
    Span4Mux_v I__3142 (
            .O(N__33063),
            .I(N__33060));
    Odrv4 I__3141 (
            .O(N__33060),
            .I(\pid_alt.error_i_regZ0Z_8 ));
    InMux I__3140 (
            .O(N__33057),
            .I(bfn_2_19_0_));
    CascadeMux I__3139 (
            .O(N__33054),
            .I(N__33051));
    InMux I__3138 (
            .O(N__33051),
            .I(N__33048));
    LocalMux I__3137 (
            .O(N__33048),
            .I(N__33045));
    Span4Mux_v I__3136 (
            .O(N__33045),
            .I(N__33042));
    Span4Mux_v I__3135 (
            .O(N__33042),
            .I(N__33039));
    Odrv4 I__3134 (
            .O(N__33039),
            .I(\pid_alt.error_i_regZ0Z_9 ));
    InMux I__3133 (
            .O(N__33036),
            .I(N__33027));
    InMux I__3132 (
            .O(N__33035),
            .I(N__33027));
    InMux I__3131 (
            .O(N__33034),
            .I(N__33027));
    LocalMux I__3130 (
            .O(N__33027),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_8_c_RNI9POQ ));
    InMux I__3129 (
            .O(N__33024),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_8 ));
    CascadeMux I__3128 (
            .O(N__33021),
            .I(N__33018));
    InMux I__3127 (
            .O(N__33018),
            .I(N__33015));
    LocalMux I__3126 (
            .O(N__33015),
            .I(N__33012));
    Span4Mux_v I__3125 (
            .O(N__33012),
            .I(N__33009));
    Odrv4 I__3124 (
            .O(N__33009),
            .I(\pid_alt.error_i_regZ0Z_10 ));
    InMux I__3123 (
            .O(N__33006),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_9 ));
    CascadeMux I__3122 (
            .O(N__33003),
            .I(N__33000));
    InMux I__3121 (
            .O(N__33000),
            .I(N__32997));
    LocalMux I__3120 (
            .O(N__32997),
            .I(N__32994));
    Span4Mux_v I__3119 (
            .O(N__32994),
            .I(N__32991));
    Span4Mux_v I__3118 (
            .O(N__32991),
            .I(N__32988));
    Odrv4 I__3117 (
            .O(N__32988),
            .I(\pid_alt.error_i_regZ0Z_11 ));
    InMux I__3116 (
            .O(N__32985),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_10 ));
    CascadeMux I__3115 (
            .O(N__32982),
            .I(N__32979));
    InMux I__3114 (
            .O(N__32979),
            .I(N__32976));
    LocalMux I__3113 (
            .O(N__32976),
            .I(N__32973));
    Span4Mux_v I__3112 (
            .O(N__32973),
            .I(N__32970));
    Span4Mux_v I__3111 (
            .O(N__32970),
            .I(N__32967));
    Odrv4 I__3110 (
            .O(N__32967),
            .I(\pid_alt.error_i_regZ0Z_12 ));
    InMux I__3109 (
            .O(N__32964),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_11 ));
    CascadeMux I__3108 (
            .O(N__32961),
            .I(N__32958));
    InMux I__3107 (
            .O(N__32958),
            .I(N__32955));
    LocalMux I__3106 (
            .O(N__32955),
            .I(N__32952));
    Span12Mux_v I__3105 (
            .O(N__32952),
            .I(N__32949));
    Odrv12 I__3104 (
            .O(N__32949),
            .I(\pid_alt.error_i_regZ0Z_13 ));
    InMux I__3103 (
            .O(N__32946),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_12 ));
    InMux I__3102 (
            .O(N__32943),
            .I(N__32937));
    InMux I__3101 (
            .O(N__32942),
            .I(N__32937));
    LocalMux I__3100 (
            .O(N__32937),
            .I(N__32934));
    Span4Mux_v I__3099 (
            .O(N__32934),
            .I(N__32931));
    Odrv4 I__3098 (
            .O(N__32931),
            .I(\pid_alt.error_p_regZ0Z_7 ));
    CascadeMux I__3097 (
            .O(N__32928),
            .I(N__32925));
    InMux I__3096 (
            .O(N__32925),
            .I(N__32919));
    InMux I__3095 (
            .O(N__32924),
            .I(N__32919));
    LocalMux I__3094 (
            .O(N__32919),
            .I(\pid_alt.error_d_reg_prevZ0Z_7 ));
    InMux I__3093 (
            .O(N__32916),
            .I(N__32907));
    InMux I__3092 (
            .O(N__32915),
            .I(N__32907));
    InMux I__3091 (
            .O(N__32914),
            .I(N__32907));
    LocalMux I__3090 (
            .O(N__32907),
            .I(N__32904));
    Span12Mux_s7_h I__3089 (
            .O(N__32904),
            .I(N__32901));
    Span12Mux_v I__3088 (
            .O(N__32901),
            .I(N__32898));
    Odrv12 I__3087 (
            .O(N__32898),
            .I(\pid_alt.error_d_regZ0Z_7 ));
    InMux I__3086 (
            .O(N__32895),
            .I(N__32892));
    LocalMux I__3085 (
            .O(N__32892),
            .I(\pid_alt.error_d_reg_prev_esr_RNIF2611_0Z0Z_7 ));
    InMux I__3084 (
            .O(N__32889),
            .I(N__32883));
    InMux I__3083 (
            .O(N__32888),
            .I(N__32883));
    LocalMux I__3082 (
            .O(N__32883),
            .I(N__32880));
    Span4Mux_v I__3081 (
            .O(N__32880),
            .I(N__32877));
    Odrv4 I__3080 (
            .O(N__32877),
            .I(\pid_alt.error_d_reg_prev_esr_RNICV511Z0Z_6 ));
    CascadeMux I__3079 (
            .O(N__32874),
            .I(\pid_alt.error_d_reg_prev_esr_RNIF2611_0Z0Z_7_cascade_ ));
    CascadeMux I__3078 (
            .O(N__32871),
            .I(N__32868));
    InMux I__3077 (
            .O(N__32868),
            .I(N__32865));
    LocalMux I__3076 (
            .O(N__32865),
            .I(N__32862));
    Span4Mux_v I__3075 (
            .O(N__32862),
            .I(N__32859));
    Odrv4 I__3074 (
            .O(N__32859),
            .I(\pid_alt.error_i_regZ0Z_1 ));
    InMux I__3073 (
            .O(N__32856),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_0 ));
    CascadeMux I__3072 (
            .O(N__32853),
            .I(N__32850));
    InMux I__3071 (
            .O(N__32850),
            .I(N__32847));
    LocalMux I__3070 (
            .O(N__32847),
            .I(N__32844));
    Span4Mux_v I__3069 (
            .O(N__32844),
            .I(N__32841));
    Odrv4 I__3068 (
            .O(N__32841),
            .I(\pid_alt.error_i_regZ0Z_2 ));
    InMux I__3067 (
            .O(N__32838),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_1 ));
    CascadeMux I__3066 (
            .O(N__32835),
            .I(N__32832));
    InMux I__3065 (
            .O(N__32832),
            .I(N__32829));
    LocalMux I__3064 (
            .O(N__32829),
            .I(N__32826));
    Span4Mux_v I__3063 (
            .O(N__32826),
            .I(N__32823));
    Odrv4 I__3062 (
            .O(N__32823),
            .I(\pid_alt.error_i_regZ0Z_3 ));
    InMux I__3061 (
            .O(N__32820),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_2 ));
    CascadeMux I__3060 (
            .O(N__32817),
            .I(N__32814));
    InMux I__3059 (
            .O(N__32814),
            .I(N__32811));
    LocalMux I__3058 (
            .O(N__32811),
            .I(N__32808));
    Span4Mux_v I__3057 (
            .O(N__32808),
            .I(N__32805));
    Odrv4 I__3056 (
            .O(N__32805),
            .I(\pid_alt.error_i_regZ0Z_4 ));
    InMux I__3055 (
            .O(N__32802),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_3 ));
    CascadeMux I__3054 (
            .O(N__32799),
            .I(N__32796));
    InMux I__3053 (
            .O(N__32796),
            .I(N__32793));
    LocalMux I__3052 (
            .O(N__32793),
            .I(N__32790));
    Span4Mux_v I__3051 (
            .O(N__32790),
            .I(N__32787));
    Span4Mux_v I__3050 (
            .O(N__32787),
            .I(N__32784));
    Odrv4 I__3049 (
            .O(N__32784),
            .I(\pid_alt.error_i_regZ0Z_5 ));
    InMux I__3048 (
            .O(N__32781),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_4 ));
    InMux I__3047 (
            .O(N__32778),
            .I(N__32769));
    InMux I__3046 (
            .O(N__32777),
            .I(N__32769));
    InMux I__3045 (
            .O(N__32776),
            .I(N__32769));
    LocalMux I__3044 (
            .O(N__32769),
            .I(N__32766));
    Span4Mux_v I__3043 (
            .O(N__32766),
            .I(N__32763));
    Span4Mux_v I__3042 (
            .O(N__32763),
            .I(N__32760));
    Odrv4 I__3041 (
            .O(N__32760),
            .I(\pid_alt.error_d_regZ0Z_3 ));
    CascadeMux I__3040 (
            .O(N__32757),
            .I(N__32754));
    InMux I__3039 (
            .O(N__32754),
            .I(N__32748));
    InMux I__3038 (
            .O(N__32753),
            .I(N__32748));
    LocalMux I__3037 (
            .O(N__32748),
            .I(\pid_alt.error_d_reg_prevZ0Z_3 ));
    InMux I__3036 (
            .O(N__32745),
            .I(N__32742));
    LocalMux I__3035 (
            .O(N__32742),
            .I(\pid_alt.error_d_reg_prev_esr_RNI3M511_0Z0Z_3 ));
    InMux I__3034 (
            .O(N__32739),
            .I(N__32733));
    InMux I__3033 (
            .O(N__32738),
            .I(N__32733));
    LocalMux I__3032 (
            .O(N__32733),
            .I(\pid_alt.error_d_reg_prev_esr_RNI0J511Z0Z_2 ));
    CascadeMux I__3031 (
            .O(N__32730),
            .I(\pid_alt.error_d_reg_prev_esr_RNI3M511_0Z0Z_3_cascade_ ));
    InMux I__3030 (
            .O(N__32727),
            .I(N__32721));
    InMux I__3029 (
            .O(N__32726),
            .I(N__32721));
    LocalMux I__3028 (
            .O(N__32721),
            .I(\pid_alt.error_d_reg_prev_esr_RNII5LS3Z0Z_1 ));
    InMux I__3027 (
            .O(N__32718),
            .I(N__32712));
    InMux I__3026 (
            .O(N__32717),
            .I(N__32712));
    LocalMux I__3025 (
            .O(N__32712),
            .I(N__32708));
    InMux I__3024 (
            .O(N__32711),
            .I(N__32705));
    Span4Mux_v I__3023 (
            .O(N__32708),
            .I(N__32700));
    LocalMux I__3022 (
            .O(N__32705),
            .I(N__32700));
    Span4Mux_v I__3021 (
            .O(N__32700),
            .I(N__32697));
    Span4Mux_v I__3020 (
            .O(N__32697),
            .I(N__32694));
    Odrv4 I__3019 (
            .O(N__32694),
            .I(\pid_alt.error_d_regZ0Z_8 ));
    InMux I__3018 (
            .O(N__32691),
            .I(N__32688));
    LocalMux I__3017 (
            .O(N__32688),
            .I(N__32684));
    InMux I__3016 (
            .O(N__32687),
            .I(N__32681));
    Span4Mux_v I__3015 (
            .O(N__32684),
            .I(N__32678));
    LocalMux I__3014 (
            .O(N__32681),
            .I(\pid_alt.error_d_reg_prevZ0Z_8 ));
    Odrv4 I__3013 (
            .O(N__32678),
            .I(\pid_alt.error_d_reg_prevZ0Z_8 ));
    CascadeMux I__3012 (
            .O(N__32673),
            .I(\pid_alt.error_d_reg_prev_esr_RNII5611_0Z0Z_8_cascade_ ));
    InMux I__3011 (
            .O(N__32670),
            .I(N__32667));
    LocalMux I__3010 (
            .O(N__32667),
            .I(\pid_alt.error_d_reg_prev_esr_RNIF2611Z0Z_7 ));
    InMux I__3009 (
            .O(N__32664),
            .I(N__32661));
    LocalMux I__3008 (
            .O(N__32661),
            .I(\pid_alt.error_d_reg_prev_esr_RNII5611_0Z0Z_8 ));
    CascadeMux I__3007 (
            .O(N__32658),
            .I(\pid_alt.error_d_reg_prev_esr_RNIF2611Z0Z_7_cascade_ ));
    InMux I__3006 (
            .O(N__32655),
            .I(N__32651));
    InMux I__3005 (
            .O(N__32654),
            .I(N__32648));
    LocalMux I__3004 (
            .O(N__32651),
            .I(N__32645));
    LocalMux I__3003 (
            .O(N__32648),
            .I(N__32642));
    Span4Mux_v I__3002 (
            .O(N__32645),
            .I(N__32639));
    Odrv12 I__3001 (
            .O(N__32642),
            .I(\pid_alt.error_p_regZ0Z_2 ));
    Odrv4 I__3000 (
            .O(N__32639),
            .I(\pid_alt.error_p_regZ0Z_2 ));
    InMux I__2999 (
            .O(N__32634),
            .I(N__32631));
    LocalMux I__2998 (
            .O(N__32631),
            .I(\pid_alt.error_d_reg_prev_esr_RNI0J511_0Z0Z_2 ));
    InMux I__2997 (
            .O(N__32628),
            .I(N__32616));
    InMux I__2996 (
            .O(N__32627),
            .I(N__32616));
    InMux I__2995 (
            .O(N__32626),
            .I(N__32616));
    InMux I__2994 (
            .O(N__32625),
            .I(N__32616));
    LocalMux I__2993 (
            .O(N__32616),
            .I(N__32613));
    Span4Mux_v I__2992 (
            .O(N__32613),
            .I(N__32610));
    Odrv4 I__2991 (
            .O(N__32610),
            .I(\pid_alt.error_d_regZ0Z_1 ));
    InMux I__2990 (
            .O(N__32607),
            .I(N__32602));
    InMux I__2989 (
            .O(N__32606),
            .I(N__32597));
    InMux I__2988 (
            .O(N__32605),
            .I(N__32597));
    LocalMux I__2987 (
            .O(N__32602),
            .I(\pid_alt.error_d_reg_prevZ0Z_1 ));
    LocalMux I__2986 (
            .O(N__32597),
            .I(\pid_alt.error_d_reg_prevZ0Z_1 ));
    CascadeMux I__2985 (
            .O(N__32592),
            .I(\pid_alt.error_d_reg_prev_esr_RNI0J511_0Z0Z_2_cascade_ ));
    InMux I__2984 (
            .O(N__32589),
            .I(N__32583));
    InMux I__2983 (
            .O(N__32588),
            .I(N__32583));
    LocalMux I__2982 (
            .O(N__32583),
            .I(\pid_alt.error_p_reg_esr_RNIOI4PZ0Z_0 ));
    CascadeMux I__2981 (
            .O(N__32580),
            .I(\pid_alt.un1_pid_prereg_16_0_cascade_ ));
    InMux I__2980 (
            .O(N__32577),
            .I(N__32573));
    InMux I__2979 (
            .O(N__32576),
            .I(N__32570));
    LocalMux I__2978 (
            .O(N__32573),
            .I(\pid_alt.error_d_reg_prev_esr_RNITF511_0Z0Z_1 ));
    LocalMux I__2977 (
            .O(N__32570),
            .I(\pid_alt.error_d_reg_prev_esr_RNITF511_0Z0Z_1 ));
    InMux I__2976 (
            .O(N__32565),
            .I(N__32558));
    InMux I__2975 (
            .O(N__32564),
            .I(N__32558));
    InMux I__2974 (
            .O(N__32563),
            .I(N__32555));
    LocalMux I__2973 (
            .O(N__32558),
            .I(N__32552));
    LocalMux I__2972 (
            .O(N__32555),
            .I(N__32549));
    Span4Mux_v I__2971 (
            .O(N__32552),
            .I(N__32546));
    Odrv12 I__2970 (
            .O(N__32549),
            .I(\pid_alt.error_d_regZ0Z_2 ));
    Odrv4 I__2969 (
            .O(N__32546),
            .I(\pid_alt.error_d_regZ0Z_2 ));
    InMux I__2968 (
            .O(N__32541),
            .I(N__32538));
    LocalMux I__2967 (
            .O(N__32538),
            .I(N__32534));
    InMux I__2966 (
            .O(N__32537),
            .I(N__32531));
    Odrv4 I__2965 (
            .O(N__32534),
            .I(\pid_alt.error_d_reg_prevZ0Z_2 ));
    LocalMux I__2964 (
            .O(N__32531),
            .I(\pid_alt.error_d_reg_prevZ0Z_2 ));
    InMux I__2963 (
            .O(N__32526),
            .I(N__32523));
    LocalMux I__2962 (
            .O(N__32523),
            .I(\pid_alt.error_d_reg_prev_esr_RNI3M511Z0Z_3 ));
    CascadeMux I__2961 (
            .O(N__32520),
            .I(\pid_alt.error_d_reg_prev_esr_RNI3M511Z0Z_3_cascade_ ));
    InMux I__2960 (
            .O(N__32517),
            .I(N__32514));
    LocalMux I__2959 (
            .O(N__32514),
            .I(N__32510));
    InMux I__2958 (
            .O(N__32513),
            .I(N__32507));
    Span4Mux_v I__2957 (
            .O(N__32510),
            .I(N__32504));
    LocalMux I__2956 (
            .O(N__32507),
            .I(\pid_alt.error_p_regZ0Z_4 ));
    Odrv4 I__2955 (
            .O(N__32504),
            .I(\pid_alt.error_p_regZ0Z_4 ));
    InMux I__2954 (
            .O(N__32499),
            .I(N__32495));
    InMux I__2953 (
            .O(N__32498),
            .I(N__32492));
    LocalMux I__2952 (
            .O(N__32495),
            .I(N__32489));
    LocalMux I__2951 (
            .O(N__32492),
            .I(N__32486));
    Span4Mux_v I__2950 (
            .O(N__32489),
            .I(N__32483));
    Odrv12 I__2949 (
            .O(N__32486),
            .I(\pid_alt.error_d_reg_prevZ0Z_4 ));
    Odrv4 I__2948 (
            .O(N__32483),
            .I(\pid_alt.error_d_reg_prevZ0Z_4 ));
    InMux I__2947 (
            .O(N__32478),
            .I(N__32473));
    InMux I__2946 (
            .O(N__32477),
            .I(N__32470));
    InMux I__2945 (
            .O(N__32476),
            .I(N__32467));
    LocalMux I__2944 (
            .O(N__32473),
            .I(N__32464));
    LocalMux I__2943 (
            .O(N__32470),
            .I(N__32459));
    LocalMux I__2942 (
            .O(N__32467),
            .I(N__32459));
    Span4Mux_v I__2941 (
            .O(N__32464),
            .I(N__32456));
    Span12Mux_v I__2940 (
            .O(N__32459),
            .I(N__32453));
    Span4Mux_v I__2939 (
            .O(N__32456),
            .I(N__32450));
    Odrv12 I__2938 (
            .O(N__32453),
            .I(\pid_alt.error_d_regZ0Z_4 ));
    Odrv4 I__2937 (
            .O(N__32450),
            .I(\pid_alt.error_d_regZ0Z_4 ));
    InMux I__2936 (
            .O(N__32445),
            .I(N__32439));
    InMux I__2935 (
            .O(N__32444),
            .I(N__32439));
    LocalMux I__2934 (
            .O(N__32439),
            .I(\pid_alt.error_d_reg_prev_esr_RNI6P511_0Z0Z_4 ));
    CascadeMux I__2933 (
            .O(N__32436),
            .I(\pid_alt.error_p_reg_esr_RNIOI4PZ0Z_0_cascade_ ));
    InMux I__2932 (
            .O(N__32433),
            .I(N__32430));
    LocalMux I__2931 (
            .O(N__32430),
            .I(\pid_alt.error_d_reg_prevZ0Z_0 ));
    InMux I__2930 (
            .O(N__32427),
            .I(N__32418));
    InMux I__2929 (
            .O(N__32426),
            .I(N__32418));
    InMux I__2928 (
            .O(N__32425),
            .I(N__32418));
    LocalMux I__2927 (
            .O(N__32418),
            .I(\pid_alt.error_d_regZ0Z_0 ));
    CascadeMux I__2926 (
            .O(N__32415),
            .I(N__32412));
    InMux I__2925 (
            .O(N__32412),
            .I(N__32406));
    InMux I__2924 (
            .O(N__32411),
            .I(N__32406));
    LocalMux I__2923 (
            .O(N__32406),
            .I(N__32403));
    Odrv4 I__2922 (
            .O(N__32403),
            .I(\pid_alt.error_p_regZ0Z_0 ));
    InMux I__2921 (
            .O(N__32400),
            .I(N__32397));
    LocalMux I__2920 (
            .O(N__32397),
            .I(\pid_alt.error_d_reg_prev_esr_RNITF511Z0Z_1 ));
    CascadeMux I__2919 (
            .O(N__32394),
            .I(\pid_alt.error_d_reg_prev_esr_RNITF511_0Z0Z_1_cascade_ ));
    CascadeMux I__2918 (
            .O(N__32391),
            .I(\Commands_frame_decoder.N_410_cascade_ ));
    InMux I__2917 (
            .O(N__32388),
            .I(N__32385));
    LocalMux I__2916 (
            .O(N__32385),
            .I(N__32382));
    Span4Mux_v I__2915 (
            .O(N__32382),
            .I(N__32379));
    Sp12to4 I__2914 (
            .O(N__32379),
            .I(N__32375));
    InMux I__2913 (
            .O(N__32378),
            .I(N__32372));
    Span12Mux_s3_h I__2912 (
            .O(N__32375),
            .I(N__32368));
    LocalMux I__2911 (
            .O(N__32372),
            .I(N__32365));
    InMux I__2910 (
            .O(N__32371),
            .I(N__32362));
    Span12Mux_h I__2909 (
            .O(N__32368),
            .I(N__32359));
    Span4Mux_v I__2908 (
            .O(N__32365),
            .I(N__32356));
    LocalMux I__2907 (
            .O(N__32362),
            .I(xy_kp_4));
    Odrv12 I__2906 (
            .O(N__32359),
            .I(xy_kp_4));
    Odrv4 I__2905 (
            .O(N__32356),
            .I(xy_kp_4));
    CascadeMux I__2904 (
            .O(N__32349),
            .I(\Commands_frame_decoder.source_CH3data_1_sqmuxa_cascade_ ));
    InMux I__2903 (
            .O(N__32346),
            .I(N__32340));
    InMux I__2902 (
            .O(N__32345),
            .I(N__32340));
    LocalMux I__2901 (
            .O(N__32340),
            .I(\Commands_frame_decoder.stateZ0Z_5 ));
    InMux I__2900 (
            .O(N__32337),
            .I(N__32334));
    LocalMux I__2899 (
            .O(N__32334),
            .I(N__32331));
    Odrv4 I__2898 (
            .O(N__32331),
            .I(alt_ki_2));
    InMux I__2897 (
            .O(N__32328),
            .I(N__32325));
    LocalMux I__2896 (
            .O(N__32325),
            .I(N__32322));
    Odrv4 I__2895 (
            .O(N__32322),
            .I(alt_ki_3));
    InMux I__2894 (
            .O(N__32319),
            .I(N__32316));
    LocalMux I__2893 (
            .O(N__32316),
            .I(N__32313));
    Span4Mux_s2_h I__2892 (
            .O(N__32313),
            .I(N__32310));
    Odrv4 I__2891 (
            .O(N__32310),
            .I(alt_ki_4));
    InMux I__2890 (
            .O(N__32307),
            .I(N__32304));
    LocalMux I__2889 (
            .O(N__32304),
            .I(N__32301));
    Span4Mux_s2_h I__2888 (
            .O(N__32301),
            .I(N__32298));
    Odrv4 I__2887 (
            .O(N__32298),
            .I(alt_ki_5));
    InMux I__2886 (
            .O(N__32295),
            .I(N__32292));
    LocalMux I__2885 (
            .O(N__32292),
            .I(N__32289));
    Span4Mux_s1_h I__2884 (
            .O(N__32289),
            .I(N__32286));
    Odrv4 I__2883 (
            .O(N__32286),
            .I(alt_ki_6));
    InMux I__2882 (
            .O(N__32283),
            .I(N__32280));
    LocalMux I__2881 (
            .O(N__32280),
            .I(N__32277));
    Sp12to4 I__2880 (
            .O(N__32277),
            .I(N__32274));
    Odrv12 I__2879 (
            .O(N__32274),
            .I(alt_ki_7));
    CascadeMux I__2878 (
            .O(N__32271),
            .I(\Commands_frame_decoder.state_ns_0_a3_0_1_cascade_ ));
    CascadeMux I__2877 (
            .O(N__32268),
            .I(\Commands_frame_decoder.state_ns_i_a2_2_1Z0Z_0_cascade_ ));
    InMux I__2876 (
            .O(N__32265),
            .I(\Commands_frame_decoder.un1_WDT_cry_8 ));
    InMux I__2875 (
            .O(N__32262),
            .I(\Commands_frame_decoder.un1_WDT_cry_9 ));
    InMux I__2874 (
            .O(N__32259),
            .I(\Commands_frame_decoder.un1_WDT_cry_10 ));
    InMux I__2873 (
            .O(N__32256),
            .I(\Commands_frame_decoder.un1_WDT_cry_11 ));
    InMux I__2872 (
            .O(N__32253),
            .I(\Commands_frame_decoder.un1_WDT_cry_12 ));
    InMux I__2871 (
            .O(N__32250),
            .I(\Commands_frame_decoder.un1_WDT_cry_13 ));
    InMux I__2870 (
            .O(N__32247),
            .I(\Commands_frame_decoder.un1_WDT_cry_14 ));
    InMux I__2869 (
            .O(N__32244),
            .I(N__32241));
    LocalMux I__2868 (
            .O(N__32241),
            .I(N__32238));
    Odrv4 I__2867 (
            .O(N__32238),
            .I(alt_ki_0));
    InMux I__2866 (
            .O(N__32235),
            .I(N__32232));
    LocalMux I__2865 (
            .O(N__32232),
            .I(N__32229));
    Odrv4 I__2864 (
            .O(N__32229),
            .I(alt_ki_1));
    InMux I__2863 (
            .O(N__32226),
            .I(N__32223));
    LocalMux I__2862 (
            .O(N__32223),
            .I(\Commands_frame_decoder.WDTZ0Z_0 ));
    InMux I__2861 (
            .O(N__32220),
            .I(N__32217));
    LocalMux I__2860 (
            .O(N__32217),
            .I(\Commands_frame_decoder.WDTZ0Z_1 ));
    InMux I__2859 (
            .O(N__32214),
            .I(\Commands_frame_decoder.un1_WDT_cry_0 ));
    InMux I__2858 (
            .O(N__32211),
            .I(N__32208));
    LocalMux I__2857 (
            .O(N__32208),
            .I(\Commands_frame_decoder.WDTZ0Z_2 ));
    InMux I__2856 (
            .O(N__32205),
            .I(\Commands_frame_decoder.un1_WDT_cry_1 ));
    InMux I__2855 (
            .O(N__32202),
            .I(N__32199));
    LocalMux I__2854 (
            .O(N__32199),
            .I(\Commands_frame_decoder.WDTZ0Z_3 ));
    InMux I__2853 (
            .O(N__32196),
            .I(\Commands_frame_decoder.un1_WDT_cry_2 ));
    InMux I__2852 (
            .O(N__32193),
            .I(\Commands_frame_decoder.un1_WDT_cry_3 ));
    InMux I__2851 (
            .O(N__32190),
            .I(\Commands_frame_decoder.un1_WDT_cry_4 ));
    InMux I__2850 (
            .O(N__32187),
            .I(\Commands_frame_decoder.un1_WDT_cry_5 ));
    InMux I__2849 (
            .O(N__32184),
            .I(\Commands_frame_decoder.un1_WDT_cry_6 ));
    InMux I__2848 (
            .O(N__32181),
            .I(bfn_2_10_0_));
    InMux I__2847 (
            .O(N__32178),
            .I(N__32175));
    LocalMux I__2846 (
            .O(N__32175),
            .I(N__32172));
    Odrv4 I__2845 (
            .O(N__32172),
            .I(\pid_alt.O_5_20 ));
    InMux I__2844 (
            .O(N__32169),
            .I(N__32166));
    LocalMux I__2843 (
            .O(N__32166),
            .I(N__32163));
    Span4Mux_h I__2842 (
            .O(N__32163),
            .I(N__32160));
    Odrv4 I__2841 (
            .O(N__32160),
            .I(\pid_alt.O_3_16 ));
    InMux I__2840 (
            .O(N__32157),
            .I(N__32154));
    LocalMux I__2839 (
            .O(N__32154),
            .I(N__32151));
    Span4Mux_v I__2838 (
            .O(N__32151),
            .I(N__32148));
    Odrv4 I__2837 (
            .O(N__32148),
            .I(alt_kd_1));
    InMux I__2836 (
            .O(N__32145),
            .I(N__32142));
    LocalMux I__2835 (
            .O(N__32142),
            .I(N__32139));
    Span4Mux_s2_h I__2834 (
            .O(N__32139),
            .I(N__32136));
    Odrv4 I__2833 (
            .O(N__32136),
            .I(alt_kd_4));
    InMux I__2832 (
            .O(N__32133),
            .I(N__32130));
    LocalMux I__2831 (
            .O(N__32130),
            .I(N__32127));
    Span4Mux_s2_h I__2830 (
            .O(N__32127),
            .I(N__32124));
    Odrv4 I__2829 (
            .O(N__32124),
            .I(alt_kd_3));
    InMux I__2828 (
            .O(N__32121),
            .I(N__32118));
    LocalMux I__2827 (
            .O(N__32118),
            .I(N__32115));
    Sp12to4 I__2826 (
            .O(N__32115),
            .I(N__32112));
    Span12Mux_s6_v I__2825 (
            .O(N__32112),
            .I(N__32109));
    Odrv12 I__2824 (
            .O(N__32109),
            .I(alt_kd_5));
    InMux I__2823 (
            .O(N__32106),
            .I(N__32103));
    LocalMux I__2822 (
            .O(N__32103),
            .I(N__32100));
    Span4Mux_s2_h I__2821 (
            .O(N__32100),
            .I(N__32097));
    Odrv4 I__2820 (
            .O(N__32097),
            .I(alt_kd_6));
    InMux I__2819 (
            .O(N__32094),
            .I(N__32091));
    LocalMux I__2818 (
            .O(N__32091),
            .I(N__32088));
    Span4Mux_s2_h I__2817 (
            .O(N__32088),
            .I(N__32085));
    Odrv4 I__2816 (
            .O(N__32085),
            .I(alt_kd_2));
    InMux I__2815 (
            .O(N__32082),
            .I(N__32079));
    LocalMux I__2814 (
            .O(N__32079),
            .I(N__32076));
    Span4Mux_s2_h I__2813 (
            .O(N__32076),
            .I(N__32073));
    Odrv4 I__2812 (
            .O(N__32073),
            .I(alt_kd_7));
    InMux I__2811 (
            .O(N__32070),
            .I(N__32067));
    LocalMux I__2810 (
            .O(N__32067),
            .I(N__32064));
    Odrv4 I__2809 (
            .O(N__32064),
            .I(\pid_alt.O_5_19 ));
    InMux I__2808 (
            .O(N__32061),
            .I(N__32058));
    LocalMux I__2807 (
            .O(N__32058),
            .I(N__32055));
    Odrv4 I__2806 (
            .O(N__32055),
            .I(\pid_alt.O_5_13 ));
    InMux I__2805 (
            .O(N__32052),
            .I(N__32049));
    LocalMux I__2804 (
            .O(N__32049),
            .I(N__32046));
    Odrv4 I__2803 (
            .O(N__32046),
            .I(\pid_alt.O_5_17 ));
    InMux I__2802 (
            .O(N__32043),
            .I(N__32040));
    LocalMux I__2801 (
            .O(N__32040),
            .I(N__32037));
    Odrv4 I__2800 (
            .O(N__32037),
            .I(\pid_alt.O_5_18 ));
    InMux I__2799 (
            .O(N__32034),
            .I(N__32031));
    LocalMux I__2798 (
            .O(N__32031),
            .I(N__32028));
    Odrv4 I__2797 (
            .O(N__32028),
            .I(\pid_alt.O_5_22 ));
    InMux I__2796 (
            .O(N__32025),
            .I(N__32019));
    InMux I__2795 (
            .O(N__32024),
            .I(N__32019));
    LocalMux I__2794 (
            .O(N__32019),
            .I(N__32016));
    Odrv12 I__2793 (
            .O(N__32016),
            .I(\pid_alt.error_p_regZ0Z_18 ));
    InMux I__2792 (
            .O(N__32013),
            .I(N__32010));
    LocalMux I__2791 (
            .O(N__32010),
            .I(\pid_alt.O_5_9 ));
    InMux I__2790 (
            .O(N__32007),
            .I(N__32004));
    LocalMux I__2789 (
            .O(N__32004),
            .I(\pid_alt.O_5_10 ));
    InMux I__2788 (
            .O(N__32001),
            .I(N__31998));
    LocalMux I__2787 (
            .O(N__31998),
            .I(\pid_alt.O_5_11 ));
    InMux I__2786 (
            .O(N__31995),
            .I(N__31992));
    LocalMux I__2785 (
            .O(N__31992),
            .I(N__31989));
    Odrv4 I__2784 (
            .O(N__31989),
            .I(\pid_alt.O_5_23 ));
    InMux I__2783 (
            .O(N__31986),
            .I(N__31983));
    LocalMux I__2782 (
            .O(N__31983),
            .I(N__31980));
    Odrv4 I__2781 (
            .O(N__31980),
            .I(\pid_alt.O_5_6 ));
    InMux I__2780 (
            .O(N__31977),
            .I(N__31971));
    InMux I__2779 (
            .O(N__31976),
            .I(N__31971));
    LocalMux I__2778 (
            .O(N__31971),
            .I(N__31968));
    Odrv4 I__2777 (
            .O(N__31968),
            .I(\pid_alt.error_d_reg_prev_esr_RNI20IMZ0Z_17 ));
    InMux I__2776 (
            .O(N__31965),
            .I(N__31962));
    LocalMux I__2775 (
            .O(N__31962),
            .I(N__31959));
    Span4Mux_h I__2774 (
            .O(N__31959),
            .I(N__31956));
    Odrv4 I__2773 (
            .O(N__31956),
            .I(\pid_alt.O_5_21 ));
    InMux I__2772 (
            .O(N__31953),
            .I(N__31950));
    LocalMux I__2771 (
            .O(N__31950),
            .I(N__31947));
    Odrv4 I__2770 (
            .O(N__31947),
            .I(\pid_alt.O_5_8 ));
    InMux I__2769 (
            .O(N__31944),
            .I(N__31941));
    LocalMux I__2768 (
            .O(N__31941),
            .I(N__31938));
    Span4Mux_h I__2767 (
            .O(N__31938),
            .I(N__31935));
    Odrv4 I__2766 (
            .O(N__31935),
            .I(\pid_alt.O_5_24 ));
    InMux I__2765 (
            .O(N__31932),
            .I(N__31929));
    LocalMux I__2764 (
            .O(N__31929),
            .I(N__31926));
    Odrv4 I__2763 (
            .O(N__31926),
            .I(\pid_alt.O_5_16 ));
    InMux I__2762 (
            .O(N__31923),
            .I(N__31920));
    LocalMux I__2761 (
            .O(N__31920),
            .I(N__31917));
    Odrv4 I__2760 (
            .O(N__31917),
            .I(\pid_alt.O_5_14 ));
    InMux I__2759 (
            .O(N__31914),
            .I(N__31908));
    InMux I__2758 (
            .O(N__31913),
            .I(N__31908));
    LocalMux I__2757 (
            .O(N__31908),
            .I(N__31905));
    Odrv12 I__2756 (
            .O(N__31905),
            .I(\pid_alt.error_p_regZ0Z_10 ));
    InMux I__2755 (
            .O(N__31902),
            .I(N__31899));
    LocalMux I__2754 (
            .O(N__31899),
            .I(N__31896));
    Odrv4 I__2753 (
            .O(N__31896),
            .I(\pid_alt.O_5_15 ));
    InMux I__2752 (
            .O(N__31893),
            .I(N__31887));
    InMux I__2751 (
            .O(N__31892),
            .I(N__31887));
    LocalMux I__2750 (
            .O(N__31887),
            .I(N__31884));
    Odrv12 I__2749 (
            .O(N__31884),
            .I(\pid_alt.error_p_regZ0Z_11 ));
    InMux I__2748 (
            .O(N__31881),
            .I(N__31878));
    LocalMux I__2747 (
            .O(N__31878),
            .I(\pid_alt.error_d_reg_prev_esr_RNI53IM_0Z0Z_18 ));
    CascadeMux I__2746 (
            .O(N__31875),
            .I(\pid_alt.error_d_reg_prev_esr_RNI53IM_0Z0Z_18_cascade_ ));
    CascadeMux I__2745 (
            .O(N__31872),
            .I(\pid_alt.error_d_reg_prev_esr_RNII5611Z0Z_8_cascade_ ));
    InMux I__2744 (
            .O(N__31869),
            .I(N__31866));
    LocalMux I__2743 (
            .O(N__31866),
            .I(\pid_alt.error_d_reg_prev_esr_RNIL8611_0Z0Z_9 ));
    InMux I__2742 (
            .O(N__31863),
            .I(N__31860));
    LocalMux I__2741 (
            .O(N__31860),
            .I(\pid_alt.error_d_reg_prev_esr_RNII5611Z0Z_8 ));
    CascadeMux I__2740 (
            .O(N__31857),
            .I(\pid_alt.error_d_reg_prev_esr_RNIL8611_0Z0Z_9_cascade_ ));
    InMux I__2739 (
            .O(N__31854),
            .I(N__31848));
    InMux I__2738 (
            .O(N__31853),
            .I(N__31848));
    LocalMux I__2737 (
            .O(N__31848),
            .I(\pid_alt.error_d_reg_prevZ0Z_11 ));
    InMux I__2736 (
            .O(N__31845),
            .I(N__31840));
    InMux I__2735 (
            .O(N__31844),
            .I(N__31835));
    InMux I__2734 (
            .O(N__31843),
            .I(N__31835));
    LocalMux I__2733 (
            .O(N__31840),
            .I(N__31830));
    LocalMux I__2732 (
            .O(N__31835),
            .I(N__31830));
    Odrv12 I__2731 (
            .O(N__31830),
            .I(\pid_alt.error_d_regZ0Z_11 ));
    CascadeMux I__2730 (
            .O(N__31827),
            .I(\pid_alt.error_d_reg_prev_esr_RNI86IM_0Z0Z_19_cascade_ ));
    InMux I__2729 (
            .O(N__31824),
            .I(N__31821));
    LocalMux I__2728 (
            .O(N__31821),
            .I(\pid_alt.error_d_reg_prev_esr_RNI53IMZ0Z_18 ));
    InMux I__2727 (
            .O(N__31818),
            .I(N__31815));
    LocalMux I__2726 (
            .O(N__31815),
            .I(\pid_alt.error_d_reg_prev_esr_RNI86IM_0Z0Z_19 ));
    CascadeMux I__2725 (
            .O(N__31812),
            .I(\pid_alt.error_d_reg_prev_esr_RNI53IMZ0Z_18_cascade_ ));
    CascadeMux I__2724 (
            .O(N__31809),
            .I(N__31806));
    InMux I__2723 (
            .O(N__31806),
            .I(N__31800));
    InMux I__2722 (
            .O(N__31805),
            .I(N__31800));
    LocalMux I__2721 (
            .O(N__31800),
            .I(\pid_alt.error_d_reg_prevZ0Z_18 ));
    InMux I__2720 (
            .O(N__31797),
            .I(N__31788));
    InMux I__2719 (
            .O(N__31796),
            .I(N__31788));
    InMux I__2718 (
            .O(N__31795),
            .I(N__31788));
    LocalMux I__2717 (
            .O(N__31788),
            .I(N__31785));
    Span4Mux_v I__2716 (
            .O(N__31785),
            .I(N__31782));
    Span4Mux_v I__2715 (
            .O(N__31782),
            .I(N__31779));
    Span4Mux_v I__2714 (
            .O(N__31779),
            .I(N__31776));
    Odrv4 I__2713 (
            .O(N__31776),
            .I(\pid_alt.error_d_regZ0Z_18 ));
    InMux I__2712 (
            .O(N__31773),
            .I(N__31770));
    LocalMux I__2711 (
            .O(N__31770),
            .I(\pid_front.O_0_8 ));
    InMux I__2710 (
            .O(N__31767),
            .I(N__31764));
    LocalMux I__2709 (
            .O(N__31764),
            .I(\pid_front.O_0_9 ));
    CascadeMux I__2708 (
            .O(N__31761),
            .I(\pid_alt.error_d_reg_prev_esr_RNIGDHM_0Z0Z_11_cascade_ ));
    InMux I__2707 (
            .O(N__31758),
            .I(N__31755));
    LocalMux I__2706 (
            .O(N__31755),
            .I(\pid_alt.error_d_reg_prev_esr_RNIDAHMZ0Z_10 ));
    InMux I__2705 (
            .O(N__31752),
            .I(N__31749));
    LocalMux I__2704 (
            .O(N__31749),
            .I(\pid_alt.error_d_reg_prev_esr_RNIGDHM_0Z0Z_11 ));
    CascadeMux I__2703 (
            .O(N__31746),
            .I(\pid_alt.error_d_reg_prev_esr_RNIDAHMZ0Z_10_cascade_ ));
    InMux I__2702 (
            .O(N__31743),
            .I(N__31737));
    InMux I__2701 (
            .O(N__31742),
            .I(N__31737));
    LocalMux I__2700 (
            .O(N__31737),
            .I(\pid_alt.error_d_reg_prevZ0Z_10 ));
    InMux I__2699 (
            .O(N__31734),
            .I(N__31725));
    InMux I__2698 (
            .O(N__31733),
            .I(N__31725));
    InMux I__2697 (
            .O(N__31732),
            .I(N__31725));
    LocalMux I__2696 (
            .O(N__31725),
            .I(N__31722));
    Odrv12 I__2695 (
            .O(N__31722),
            .I(\pid_alt.error_d_regZ0Z_10 ));
    InMux I__2694 (
            .O(N__31719),
            .I(N__31716));
    LocalMux I__2693 (
            .O(N__31716),
            .I(N__31713));
    Odrv4 I__2692 (
            .O(N__31713),
            .I(\pid_front.O_0_19 ));
    InMux I__2691 (
            .O(N__31710),
            .I(N__31707));
    LocalMux I__2690 (
            .O(N__31707),
            .I(N__31704));
    Odrv4 I__2689 (
            .O(N__31704),
            .I(\pid_front.O_0_10 ));
    InMux I__2688 (
            .O(N__31701),
            .I(N__31698));
    LocalMux I__2687 (
            .O(N__31698),
            .I(N__31695));
    Odrv4 I__2686 (
            .O(N__31695),
            .I(\pid_front.O_0_21 ));
    InMux I__2685 (
            .O(N__31692),
            .I(N__31689));
    LocalMux I__2684 (
            .O(N__31689),
            .I(N__31686));
    Odrv4 I__2683 (
            .O(N__31686),
            .I(\pid_front.O_0_22 ));
    InMux I__2682 (
            .O(N__31683),
            .I(N__31680));
    LocalMux I__2681 (
            .O(N__31680),
            .I(\pid_front.O_0_5 ));
    InMux I__2680 (
            .O(N__31677),
            .I(N__31674));
    LocalMux I__2679 (
            .O(N__31674),
            .I(N__31671));
    Odrv4 I__2678 (
            .O(N__31671),
            .I(\pid_front.O_0_23 ));
    InMux I__2677 (
            .O(N__31668),
            .I(N__31665));
    LocalMux I__2676 (
            .O(N__31665),
            .I(N__31662));
    Odrv4 I__2675 (
            .O(N__31662),
            .I(\pid_front.O_0_24 ));
    InMux I__2674 (
            .O(N__31659),
            .I(N__31656));
    LocalMux I__2673 (
            .O(N__31656),
            .I(\pid_front.O_0_11 ));
    InMux I__2672 (
            .O(N__31653),
            .I(N__31650));
    LocalMux I__2671 (
            .O(N__31650),
            .I(\pid_front.O_0_7 ));
    InMux I__2670 (
            .O(N__31647),
            .I(N__31644));
    LocalMux I__2669 (
            .O(N__31644),
            .I(N__31641));
    Odrv4 I__2668 (
            .O(N__31641),
            .I(\pid_alt.O_4_4 ));
    InMux I__2667 (
            .O(N__31638),
            .I(N__31635));
    LocalMux I__2666 (
            .O(N__31635),
            .I(N__31632));
    Span4Mux_v I__2665 (
            .O(N__31632),
            .I(N__31629));
    Span4Mux_v I__2664 (
            .O(N__31629),
            .I(N__31626));
    Span4Mux_v I__2663 (
            .O(N__31626),
            .I(N__31623));
    Odrv4 I__2662 (
            .O(N__31623),
            .I(\pid_alt.O_5_4 ));
    InMux I__2661 (
            .O(N__31620),
            .I(N__31617));
    LocalMux I__2660 (
            .O(N__31617),
            .I(N__31614));
    Span4Mux_h I__2659 (
            .O(N__31614),
            .I(N__31611));
    Odrv4 I__2658 (
            .O(N__31611),
            .I(\pid_alt.O_4_5 ));
    InMux I__2657 (
            .O(N__31608),
            .I(N__31605));
    LocalMux I__2656 (
            .O(N__31605),
            .I(N__31602));
    Span4Mux_v I__2655 (
            .O(N__31602),
            .I(N__31599));
    Span4Mux_v I__2654 (
            .O(N__31599),
            .I(N__31596));
    Odrv4 I__2653 (
            .O(N__31596),
            .I(\pid_alt.O_3_4 ));
    InMux I__2652 (
            .O(N__31593),
            .I(N__31590));
    LocalMux I__2651 (
            .O(N__31590),
            .I(N__31587));
    Odrv4 I__2650 (
            .O(N__31587),
            .I(\pid_front.O_0_14 ));
    InMux I__2649 (
            .O(N__31584),
            .I(N__31581));
    LocalMux I__2648 (
            .O(N__31581),
            .I(N__31578));
    Odrv4 I__2647 (
            .O(N__31578),
            .I(\pid_front.O_0_15 ));
    InMux I__2646 (
            .O(N__31575),
            .I(N__31572));
    LocalMux I__2645 (
            .O(N__31572),
            .I(N__31569));
    Span4Mux_h I__2644 (
            .O(N__31569),
            .I(N__31566));
    Odrv4 I__2643 (
            .O(N__31566),
            .I(\pid_front.O_0_16 ));
    InMux I__2642 (
            .O(N__31563),
            .I(N__31560));
    LocalMux I__2641 (
            .O(N__31560),
            .I(N__31557));
    Odrv4 I__2640 (
            .O(N__31557),
            .I(\pid_front.O_0_17 ));
    InMux I__2639 (
            .O(N__31554),
            .I(N__31551));
    LocalMux I__2638 (
            .O(N__31551),
            .I(N__31548));
    Odrv4 I__2637 (
            .O(N__31548),
            .I(\pid_front.O_0_18 ));
    InMux I__2636 (
            .O(N__31545),
            .I(N__31542));
    LocalMux I__2635 (
            .O(N__31542),
            .I(\pid_alt.O_4_20 ));
    InMux I__2634 (
            .O(N__31539),
            .I(N__31536));
    LocalMux I__2633 (
            .O(N__31536),
            .I(\pid_alt.O_4_21 ));
    InMux I__2632 (
            .O(N__31533),
            .I(N__31530));
    LocalMux I__2631 (
            .O(N__31530),
            .I(\pid_alt.O_4_22 ));
    InMux I__2630 (
            .O(N__31527),
            .I(N__31524));
    LocalMux I__2629 (
            .O(N__31524),
            .I(\pid_alt.O_4_23 ));
    InMux I__2628 (
            .O(N__31521),
            .I(N__31518));
    LocalMux I__2627 (
            .O(N__31518),
            .I(\pid_alt.O_4_6 ));
    InMux I__2626 (
            .O(N__31515),
            .I(N__31512));
    LocalMux I__2625 (
            .O(N__31512),
            .I(N__31509));
    Odrv4 I__2624 (
            .O(N__31509),
            .I(\pid_alt.O_4_24 ));
    InMux I__2623 (
            .O(N__31506),
            .I(N__31503));
    LocalMux I__2622 (
            .O(N__31503),
            .I(N__31500));
    Odrv4 I__2621 (
            .O(N__31500),
            .I(\pid_alt.O_4_7 ));
    InMux I__2620 (
            .O(N__31497),
            .I(N__31494));
    LocalMux I__2619 (
            .O(N__31494),
            .I(\pid_alt.O_4_8 ));
    InMux I__2618 (
            .O(N__31491),
            .I(N__31488));
    LocalMux I__2617 (
            .O(N__31488),
            .I(\pid_alt.O_4_9 ));
    InMux I__2616 (
            .O(N__31485),
            .I(N__31482));
    LocalMux I__2615 (
            .O(N__31482),
            .I(\pid_alt.O_4_14 ));
    InMux I__2614 (
            .O(N__31479),
            .I(N__31476));
    LocalMux I__2613 (
            .O(N__31476),
            .I(N__31473));
    Odrv4 I__2612 (
            .O(N__31473),
            .I(\pid_alt.O_3_12 ));
    InMux I__2611 (
            .O(N__31470),
            .I(N__31467));
    LocalMux I__2610 (
            .O(N__31467),
            .I(\pid_alt.O_4_12 ));
    InMux I__2609 (
            .O(N__31464),
            .I(N__31461));
    LocalMux I__2608 (
            .O(N__31461),
            .I(\pid_alt.O_4_13 ));
    InMux I__2607 (
            .O(N__31458),
            .I(N__31455));
    LocalMux I__2606 (
            .O(N__31455),
            .I(\pid_alt.O_4_10 ));
    InMux I__2605 (
            .O(N__31452),
            .I(N__31449));
    LocalMux I__2604 (
            .O(N__31449),
            .I(\pid_alt.O_4_15 ));
    InMux I__2603 (
            .O(N__31446),
            .I(N__31443));
    LocalMux I__2602 (
            .O(N__31443),
            .I(N__31440));
    Odrv4 I__2601 (
            .O(N__31440),
            .I(\pid_alt.O_4_16 ));
    InMux I__2600 (
            .O(N__31437),
            .I(N__31434));
    LocalMux I__2599 (
            .O(N__31434),
            .I(N__31431));
    Odrv4 I__2598 (
            .O(N__31431),
            .I(\pid_alt.O_4_17 ));
    InMux I__2597 (
            .O(N__31428),
            .I(N__31425));
    LocalMux I__2596 (
            .O(N__31425),
            .I(\pid_alt.O_4_18 ));
    InMux I__2595 (
            .O(N__31422),
            .I(N__31419));
    LocalMux I__2594 (
            .O(N__31419),
            .I(\pid_alt.O_4_19 ));
    InMux I__2593 (
            .O(N__31416),
            .I(N__31413));
    LocalMux I__2592 (
            .O(N__31413),
            .I(\pid_alt.O_3_19 ));
    InMux I__2591 (
            .O(N__31410),
            .I(N__31407));
    LocalMux I__2590 (
            .O(N__31407),
            .I(\pid_alt.O_3_8 ));
    InMux I__2589 (
            .O(N__31404),
            .I(N__31401));
    LocalMux I__2588 (
            .O(N__31401),
            .I(\pid_alt.O_3_7 ));
    InMux I__2587 (
            .O(N__31398),
            .I(N__31395));
    LocalMux I__2586 (
            .O(N__31395),
            .I(\pid_alt.O_3_10 ));
    InMux I__2585 (
            .O(N__31392),
            .I(N__31389));
    LocalMux I__2584 (
            .O(N__31389),
            .I(\pid_alt.O_3_9 ));
    InMux I__2583 (
            .O(N__31386),
            .I(N__31383));
    LocalMux I__2582 (
            .O(N__31383),
            .I(\pid_alt.O_3_14 ));
    InMux I__2581 (
            .O(N__31380),
            .I(N__31377));
    LocalMux I__2580 (
            .O(N__31377),
            .I(N__31374));
    Odrv4 I__2579 (
            .O(N__31374),
            .I(\pid_alt.O_3_13 ));
    InMux I__2578 (
            .O(N__31371),
            .I(N__31368));
    LocalMux I__2577 (
            .O(N__31368),
            .I(N__31365));
    Odrv4 I__2576 (
            .O(N__31365),
            .I(\pid_alt.O_3_6 ));
    InMux I__2575 (
            .O(N__31362),
            .I(N__31359));
    LocalMux I__2574 (
            .O(N__31359),
            .I(N__31356));
    Span4Mux_v I__2573 (
            .O(N__31356),
            .I(N__31353));
    Odrv4 I__2572 (
            .O(N__31353),
            .I(\pid_alt.O_3_5 ));
    InMux I__2571 (
            .O(N__31350),
            .I(N__31347));
    LocalMux I__2570 (
            .O(N__31347),
            .I(N__31344));
    Odrv4 I__2569 (
            .O(N__31344),
            .I(\pid_alt.O_3_21 ));
    InMux I__2568 (
            .O(N__31341),
            .I(N__31338));
    LocalMux I__2567 (
            .O(N__31338),
            .I(N__31335));
    Odrv4 I__2566 (
            .O(N__31335),
            .I(\pid_alt.O_3_18 ));
    InMux I__2565 (
            .O(N__31332),
            .I(N__31329));
    LocalMux I__2564 (
            .O(N__31329),
            .I(\pid_alt.O_3_11 ));
    InMux I__2563 (
            .O(N__31326),
            .I(N__31323));
    LocalMux I__2562 (
            .O(N__31323),
            .I(\pid_alt.O_3_15 ));
    InMux I__2561 (
            .O(N__31320),
            .I(N__31317));
    LocalMux I__2560 (
            .O(N__31317),
            .I(N__31314));
    Odrv4 I__2559 (
            .O(N__31314),
            .I(\pid_alt.O_3_17 ));
    InMux I__2558 (
            .O(N__31311),
            .I(N__31308));
    LocalMux I__2557 (
            .O(N__31308),
            .I(N__31305));
    Odrv4 I__2556 (
            .O(N__31305),
            .I(\pid_alt.O_3_24 ));
    InMux I__2555 (
            .O(N__31302),
            .I(N__31299));
    LocalMux I__2554 (
            .O(N__31299),
            .I(\pid_alt.O_3_20 ));
    InMux I__2553 (
            .O(N__31296),
            .I(N__31293));
    LocalMux I__2552 (
            .O(N__31293),
            .I(\pid_alt.O_3_22 ));
    InMux I__2551 (
            .O(N__31290),
            .I(N__31287));
    LocalMux I__2550 (
            .O(N__31287),
            .I(\pid_alt.O_3_23 ));
    InMux I__2549 (
            .O(N__31284),
            .I(N__31281));
    LocalMux I__2548 (
            .O(N__31281),
            .I(N__31278));
    Span4Mux_h I__2547 (
            .O(N__31278),
            .I(N__31275));
    Span4Mux_v I__2546 (
            .O(N__31275),
            .I(N__31272));
    Odrv4 I__2545 (
            .O(N__31272),
            .I(\pid_alt.O_4_11 ));
    IoInMux I__2544 (
            .O(N__31269),
            .I(N__31266));
    LocalMux I__2543 (
            .O(N__31266),
            .I(N__31263));
    Span4Mux_s0_v I__2542 (
            .O(N__31263),
            .I(N__31260));
    Sp12to4 I__2541 (
            .O(N__31260),
            .I(N__31257));
    Span12Mux_h I__2540 (
            .O(N__31257),
            .I(N__31254));
    Span12Mux_v I__2539 (
            .O(N__31254),
            .I(N__31251));
    Span12Mux_v I__2538 (
            .O(N__31251),
            .I(N__31248));
    Span12Mux_h I__2537 (
            .O(N__31248),
            .I(N__31245));
    Odrv12 I__2536 (
            .O(N__31245),
            .I(\Pc2drone_pll_inst.clk_system_pll ));
    defparam IN_MUX_bfv_17_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_11_0_));
    defparam IN_MUX_bfv_17_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_12_0_ (
            .carryinitin(\pid_side.un1_pid_prereg_0_cry_6 ),
            .carryinitout(bfn_17_12_0_));
    defparam IN_MUX_bfv_17_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_13_0_ (
            .carryinitin(\pid_side.un1_pid_prereg_0_cry_14 ),
            .carryinitout(bfn_17_13_0_));
    defparam IN_MUX_bfv_17_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_14_0_ (
            .carryinitin(\pid_side.un1_pid_prereg_0_cry_22 ),
            .carryinitout(bfn_17_14_0_));
    defparam IN_MUX_bfv_9_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_17_0_));
    defparam IN_MUX_bfv_9_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_18_0_ (
            .carryinitin(\pid_front.un1_pid_prereg_0_cry_6 ),
            .carryinitout(bfn_9_18_0_));
    defparam IN_MUX_bfv_9_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_19_0_ (
            .carryinitin(\pid_front.un1_pid_prereg_0_cry_14 ),
            .carryinitout(bfn_9_19_0_));
    defparam IN_MUX_bfv_9_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_20_0_ (
            .carryinitin(\pid_front.un1_pid_prereg_0_cry_22 ),
            .carryinitout(bfn_9_20_0_));
    defparam IN_MUX_bfv_3_15_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_15_0_));
    defparam IN_MUX_bfv_3_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_16_0_ (
            .carryinitin(\pid_alt.un1_pid_prereg_0_cry_6 ),
            .carryinitout(bfn_3_16_0_));
    defparam IN_MUX_bfv_3_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_17_0_ (
            .carryinitin(\pid_alt.un1_pid_prereg_0_cry_14 ),
            .carryinitout(bfn_3_17_0_));
    defparam IN_MUX_bfv_3_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_18_0_ (
            .carryinitin(\pid_alt.un1_pid_prereg_0_cry_22 ),
            .carryinitout(bfn_3_18_0_));
    defparam IN_MUX_bfv_9_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_11_0_));
    defparam IN_MUX_bfv_9_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_12_0_ (
            .carryinitin(\scaler_4.un3_source_data_0_cry_7 ),
            .carryinitout(bfn_9_12_0_));
    defparam IN_MUX_bfv_9_8_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_8_0_));
    defparam IN_MUX_bfv_9_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_9_0_ (
            .carryinitin(\scaler_4.un2_source_data_0_cry_8 ),
            .carryinitout(bfn_9_9_0_));
    defparam IN_MUX_bfv_8_1_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_1_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_1_0_));
    defparam IN_MUX_bfv_8_2_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_2_0_ (
            .carryinitin(\reset_module_System.count_1_cry_8 ),
            .carryinitout(bfn_8_2_0_));
    defparam IN_MUX_bfv_8_3_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_3_0_ (
            .carryinitin(\reset_module_System.count_1_cry_16 ),
            .carryinitout(bfn_8_3_0_));
    defparam IN_MUX_bfv_8_8_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_8_0_));
    defparam IN_MUX_bfv_8_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_9_0_ (
            .carryinitin(\ppm_encoder_1.un1_throttle_cry_7 ),
            .carryinitout(bfn_8_9_0_));
    defparam IN_MUX_bfv_9_6_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_6_0_));
    defparam IN_MUX_bfv_9_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_7_0_ (
            .carryinitin(\ppm_encoder_1.un1_rudder_cry_13 ),
            .carryinitout(bfn_9_7_0_));
    defparam IN_MUX_bfv_10_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_11_0_));
    defparam IN_MUX_bfv_10_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_12_0_ (
            .carryinitin(\ppm_encoder_1.un1_elevator_cry_7 ),
            .carryinitout(bfn_10_12_0_));
    defparam IN_MUX_bfv_11_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_9_0_));
    defparam IN_MUX_bfv_11_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_10_0_ (
            .carryinitin(\ppm_encoder_1.un1_aileron_cry_7 ),
            .carryinitout(bfn_11_10_0_));
    defparam IN_MUX_bfv_10_3_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_3_0_));
    defparam IN_MUX_bfv_10_4_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_4_0_ (
            .carryinitin(\ppm_encoder_1.un1_init_pulses_0_cry_7 ),
            .carryinitout(bfn_10_4_0_));
    defparam IN_MUX_bfv_10_5_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_5_0_ (
            .carryinitin(\ppm_encoder_1.un1_init_pulses_0_cry_15 ),
            .carryinitout(bfn_10_5_0_));
    defparam IN_MUX_bfv_14_2_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_2_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_2_0_));
    defparam IN_MUX_bfv_14_3_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_3_0_ (
            .carryinitin(\ppm_encoder_1.counter24_0_data_tmp_7 ),
            .carryinitout(bfn_14_3_0_));
    defparam IN_MUX_bfv_15_8_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_8_0_));
    defparam IN_MUX_bfv_15_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_9_0_ (
            .carryinitin(\pid_side.un11lto30_i_a2_6 ),
            .carryinitout(bfn_15_9_0_));
    defparam IN_MUX_bfv_8_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_15_0_));
    defparam IN_MUX_bfv_8_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_16_0_ (
            .carryinitin(\pid_front.un11lto30_i_a2_6 ),
            .carryinitout(bfn_8_16_0_));
    defparam IN_MUX_bfv_4_18_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_18_0_));
    defparam IN_MUX_bfv_4_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_19_0_ (
            .carryinitin(\pid_alt.error_cry_7 ),
            .carryinitout(bfn_4_19_0_));
    defparam IN_MUX_bfv_7_15_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_15_0_));
    defparam IN_MUX_bfv_5_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_9_0_));
    defparam IN_MUX_bfv_16_4_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_4_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_4_0_));
    defparam IN_MUX_bfv_16_5_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_5_0_ (
            .carryinitin(\ppm_encoder_1.un1_counter_13_cry_7 ),
            .carryinitout(bfn_16_5_0_));
    defparam IN_MUX_bfv_16_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_6_0_ (
            .carryinitin(\ppm_encoder_1.un1_counter_13_cry_15 ),
            .carryinitout(bfn_16_6_0_));
    defparam IN_MUX_bfv_11_1_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_1_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_1_0_));
    defparam IN_MUX_bfv_11_2_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_2_0_ (
            .carryinitin(\ppm_encoder_1.un1_init_pulses_3_cry_7 ),
            .carryinitout(bfn_11_2_0_));
    defparam IN_MUX_bfv_11_3_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_3_0_ (
            .carryinitin(\ppm_encoder_1.un1_init_pulses_3_cry_15 ),
            .carryinitout(bfn_11_3_0_));
    defparam IN_MUX_bfv_16_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_13_0_));
    defparam IN_MUX_bfv_16_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_14_0_ (
            .carryinitin(\pid_side.un1_error_i_acumm_prereg_cry_7 ),
            .carryinitout(bfn_16_14_0_));
    defparam IN_MUX_bfv_16_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_15_0_ (
            .carryinitin(\pid_side.un1_error_i_acumm_prereg_cry_15 ),
            .carryinitout(bfn_16_15_0_));
    defparam IN_MUX_bfv_16_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_16_0_ (
            .carryinitin(\pid_side.un1_error_i_acumm_prereg_cry_23 ),
            .carryinitout(bfn_16_16_0_));
    defparam IN_MUX_bfv_18_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_17_0_));
    defparam IN_MUX_bfv_18_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_18_0_ (
            .carryinitin(\pid_side.error_cry_3_0 ),
            .carryinitout(bfn_18_18_0_));
    defparam IN_MUX_bfv_13_23_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_23_0_));
    defparam IN_MUX_bfv_13_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_24_0_ (
            .carryinitin(\pid_front.un1_error_i_acumm_prereg_cry_7 ),
            .carryinitout(bfn_13_24_0_));
    defparam IN_MUX_bfv_13_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_25_0_ (
            .carryinitin(\pid_front.un1_error_i_acumm_prereg_cry_15 ),
            .carryinitout(bfn_13_25_0_));
    defparam IN_MUX_bfv_13_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_26_0_ (
            .carryinitin(\pid_front.un1_error_i_acumm_prereg_cry_23 ),
            .carryinitout(bfn_13_26_0_));
    defparam IN_MUX_bfv_13_21_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_21_0_));
    defparam IN_MUX_bfv_13_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_22_0_ (
            .carryinitin(\pid_front.error_cry_3_0 ),
            .carryinitout(bfn_13_22_0_));
    defparam IN_MUX_bfv_2_18_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_18_0_));
    defparam IN_MUX_bfv_2_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_19_0_ (
            .carryinitin(\pid_alt.un1_error_i_acumm_prereg_cry_7 ),
            .carryinitout(bfn_2_19_0_));
    defparam IN_MUX_bfv_2_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_20_0_ (
            .carryinitin(\pid_alt.un1_error_i_acumm_prereg_cry_15 ),
            .carryinitout(bfn_2_20_0_));
    defparam IN_MUX_bfv_8_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_13_0_));
    defparam IN_MUX_bfv_8_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_14_0_ (
            .carryinitin(\dron_frame_decoder_1.un1_WDT_cry_7 ),
            .carryinitout(bfn_8_14_0_));
    defparam IN_MUX_bfv_2_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_9_0_));
    defparam IN_MUX_bfv_2_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_10_0_ (
            .carryinitin(\Commands_frame_decoder.un1_WDT_cry_7 ),
            .carryinitout(bfn_2_10_0_));
    ICE_GB \reset_module_System.reset_RNITC69  (
            .USERSIGNALTOGLOBALBUFFER(N__65943),
            .GLOBALBUFFEROUTPUT(reset_system_g));
    ICE_GB \pid_side.state_RNIL5IF_0_0  (
            .USERSIGNALTOGLOBALBUFFER(N__50652),
            .GLOBALBUFFEROUTPUT(\pid_side.N_838_g ));
    ICE_GB \pid_alt.state_RNICP2N1_0_0  (
            .USERSIGNALTOGLOBALBUFFER(N__71850),
            .GLOBALBUFFEROUTPUT(\pid_alt.N_939_0_g ));
    ICE_GB \pid_front.state_RNIM14N_0_0  (
            .USERSIGNALTOGLOBALBUFFER(N__51417),
            .GLOBALBUFFEROUTPUT(\pid_front.N_1705_g ));
    ICE_GB \Pc2drone_pll_inst.PLLOUTCORE_derived_clock_RNI5FOA  (
            .USERSIGNALTOGLOBALBUFFER(N__31269),
            .GLOBALBUFFEROUTPUT(clk_system_pll_g));
    ICE_GB \reset_module_System.reset_RNITC69_0  (
            .USERSIGNALTOGLOBALBUFFER(N__62646),
            .GLOBALBUFFEROUTPUT(N_940_g));
    ICE_GB \pid_front.state_RNIPKTD_0_0  (
            .USERSIGNALTOGLOBALBUFFER(N__46833),
            .GLOBALBUFFEROUTPUT(\pid_front.N_764_g ));
    ICE_GB \pid_alt.state_RNIH1EN_0_0  (
            .USERSIGNALTOGLOBALBUFFER(N__55989),
            .GLOBALBUFFEROUTPUT(\pid_alt.state_0_g_0 ));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \pid_alt.error_i_reg_esr_7_LC_1_4_0 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_7_LC_1_4_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_7_LC_1_4_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_7_LC_1_4_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31284),
            .lcout(\pid_alt.error_i_regZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87070),
            .ce(N__33454),
            .sr(N__86044));
    defparam \pid_alt.error_d_reg_esr_17_LC_1_4_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_17_LC_1_4_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_17_LC_1_4_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_17_LC_1_4_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31350),
            .lcout(\pid_alt.error_d_regZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87070),
            .ce(N__33454),
            .sr(N__86044));
    defparam \pid_alt.error_d_reg_esr_14_LC_1_4_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_14_LC_1_4_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_14_LC_1_4_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_14_LC_1_4_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31341),
            .lcout(\pid_alt.error_d_regZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87070),
            .ce(N__33454),
            .sr(N__86044));
    defparam \pid_alt.error_d_reg_esr_7_LC_1_5_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_7_LC_1_5_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_7_LC_1_5_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_d_reg_esr_7_LC_1_5_2  (
            .in0(N__31332),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_d_regZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87083),
            .ce(N__33456),
            .sr(N__86043));
    defparam \pid_alt.error_d_reg_esr_11_LC_1_5_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_11_LC_1_5_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_11_LC_1_5_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_11_LC_1_5_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31326),
            .lcout(\pid_alt.error_d_regZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87083),
            .ce(N__33456),
            .sr(N__86043));
    defparam \pid_alt.error_d_reg_esr_13_LC_1_5_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_13_LC_1_5_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_13_LC_1_5_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_13_LC_1_5_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31320),
            .lcout(\pid_alt.error_d_regZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87083),
            .ce(N__33456),
            .sr(N__86043));
    defparam \pid_alt.error_d_reg_esr_20_LC_1_5_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_20_LC_1_5_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_20_LC_1_5_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_20_LC_1_5_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31311),
            .lcout(\pid_alt.error_d_regZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87083),
            .ce(N__33456),
            .sr(N__86043));
    defparam \pid_alt.error_d_reg_esr_16_LC_1_6_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_16_LC_1_6_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_16_LC_1_6_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_16_LC_1_6_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31302),
            .lcout(\pid_alt.error_d_regZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87097),
            .ce(N__33457),
            .sr(N__86041));
    defparam \pid_alt.error_d_reg_esr_18_LC_1_6_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_18_LC_1_6_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_18_LC_1_6_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_18_LC_1_6_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31296),
            .lcout(\pid_alt.error_d_regZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87097),
            .ce(N__33457),
            .sr(N__86041));
    defparam \pid_alt.error_d_reg_esr_19_LC_1_6_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_19_LC_1_6_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_19_LC_1_6_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_19_LC_1_6_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31290),
            .lcout(\pid_alt.error_d_regZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87097),
            .ce(N__33457),
            .sr(N__86041));
    defparam \pid_alt.error_d_reg_esr_15_LC_1_6_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_15_LC_1_6_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_15_LC_1_6_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_15_LC_1_6_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31416),
            .lcout(\pid_alt.error_d_regZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87097),
            .ce(N__33457),
            .sr(N__86041));
    defparam \pid_alt.error_d_reg_esr_4_LC_1_6_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_4_LC_1_6_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_4_LC_1_6_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_4_LC_1_6_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31410),
            .lcout(\pid_alt.error_d_regZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87097),
            .ce(N__33457),
            .sr(N__86041));
    defparam \pid_alt.error_d_reg_esr_3_LC_1_6_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_3_LC_1_6_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_3_LC_1_6_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_3_LC_1_6_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31404),
            .lcout(\pid_alt.error_d_regZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87097),
            .ce(N__33457),
            .sr(N__86041));
    defparam \pid_alt.error_d_reg_esr_6_LC_1_6_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_6_LC_1_6_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_6_LC_1_6_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_6_LC_1_6_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31398),
            .lcout(\pid_alt.error_d_regZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87097),
            .ce(N__33457),
            .sr(N__86041));
    defparam \pid_alt.error_d_reg_esr_5_LC_1_7_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_5_LC_1_7_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_5_LC_1_7_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_5_LC_1_7_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31392),
            .lcout(\pid_alt.error_d_regZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87112),
            .ce(N__33458),
            .sr(N__86040));
    defparam \pid_alt.error_d_reg_esr_10_LC_1_7_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_10_LC_1_7_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_10_LC_1_7_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_10_LC_1_7_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31386),
            .lcout(\pid_alt.error_d_regZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87112),
            .ce(N__33458),
            .sr(N__86040));
    defparam \pid_alt.error_d_reg_esr_9_LC_1_8_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_9_LC_1_8_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_9_LC_1_8_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_9_LC_1_8_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31380),
            .lcout(\pid_alt.error_d_regZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87126),
            .ce(N__33459),
            .sr(N__86039));
    defparam \pid_alt.error_d_reg_esr_2_LC_1_8_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_2_LC_1_8_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_2_LC_1_8_3 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \pid_alt.error_d_reg_esr_2_LC_1_8_3  (
            .in0(_gnd_net_),
            .in1(N__31371),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_d_regZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87126),
            .ce(N__33459),
            .sr(N__86039));
    defparam \pid_alt.error_d_reg_esr_1_LC_1_9_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_1_LC_1_9_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_1_LC_1_9_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_1_LC_1_9_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31362),
            .lcout(\pid_alt.error_d_regZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87141),
            .ce(N__33460),
            .sr(N__86038));
    defparam \pid_alt.error_d_reg_esr_8_LC_1_9_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_8_LC_1_9_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_8_LC_1_9_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_8_LC_1_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31479),
            .lcout(\pid_alt.error_d_regZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87141),
            .ce(N__33460),
            .sr(N__86038));
    defparam \pid_alt.error_i_reg_esr_8_LC_1_10_0 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_8_LC_1_10_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_8_LC_1_10_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_8_LC_1_10_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31470),
            .lcout(\pid_alt.error_i_regZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87159),
            .ce(N__33461),
            .sr(N__86037));
    defparam \pid_alt.error_i_reg_esr_9_LC_1_10_2 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_9_LC_1_10_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_9_LC_1_10_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_9_LC_1_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31464),
            .lcout(\pid_alt.error_i_regZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87159),
            .ce(N__33461),
            .sr(N__86037));
    defparam \pid_alt.error_i_reg_esr_6_LC_1_10_4 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_6_LC_1_10_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_6_LC_1_10_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_6_LC_1_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31458),
            .lcout(\pid_alt.error_i_regZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87159),
            .ce(N__33461),
            .sr(N__86037));
    defparam \pid_alt.error_i_reg_esr_11_LC_1_10_5 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_11_LC_1_10_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_11_LC_1_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_11_LC_1_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31452),
            .lcout(\pid_alt.error_i_regZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87159),
            .ce(N__33461),
            .sr(N__86037));
    defparam \pid_alt.error_i_reg_esr_12_LC_1_10_6 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_12_LC_1_10_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_12_LC_1_10_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_12_LC_1_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31446),
            .lcout(\pid_alt.error_i_regZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87159),
            .ce(N__33461),
            .sr(N__86037));
    defparam \pid_alt.error_i_reg_esr_13_LC_1_10_7 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_13_LC_1_10_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_13_LC_1_10_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_13_LC_1_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31437),
            .lcout(\pid_alt.error_i_regZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87159),
            .ce(N__33461),
            .sr(N__86037));
    defparam \pid_alt.error_i_reg_esr_14_LC_1_11_0 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_14_LC_1_11_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_14_LC_1_11_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_14_LC_1_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31428),
            .lcout(\pid_alt.error_i_regZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87173),
            .ce(N__33462),
            .sr(N__86036));
    defparam \pid_alt.error_i_reg_esr_15_LC_1_11_1 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_15_LC_1_11_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_15_LC_1_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_15_LC_1_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31422),
            .lcout(\pid_alt.error_i_regZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87173),
            .ce(N__33462),
            .sr(N__86036));
    defparam \pid_alt.error_i_reg_esr_16_LC_1_11_2 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_16_LC_1_11_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_16_LC_1_11_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_16_LC_1_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31545),
            .lcout(\pid_alt.error_i_regZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87173),
            .ce(N__33462),
            .sr(N__86036));
    defparam \pid_alt.error_i_reg_esr_17_LC_1_11_3 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_17_LC_1_11_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_17_LC_1_11_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_17_LC_1_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31539),
            .lcout(\pid_alt.error_i_regZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87173),
            .ce(N__33462),
            .sr(N__86036));
    defparam \pid_alt.error_i_reg_esr_18_LC_1_11_4 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_18_LC_1_11_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_18_LC_1_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_18_LC_1_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31533),
            .lcout(\pid_alt.error_i_regZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87173),
            .ce(N__33462),
            .sr(N__86036));
    defparam \pid_alt.error_i_reg_esr_19_LC_1_11_5 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_19_LC_1_11_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_19_LC_1_11_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_19_LC_1_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31527),
            .lcout(\pid_alt.error_i_regZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87173),
            .ce(N__33462),
            .sr(N__86036));
    defparam \pid_alt.error_i_reg_esr_2_LC_1_11_6 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_2_LC_1_11_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_2_LC_1_11_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_i_reg_esr_2_LC_1_11_6  (
            .in0(N__31521),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_i_regZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87173),
            .ce(N__33462),
            .sr(N__86036));
    defparam \pid_alt.error_i_reg_esr_20_LC_1_11_7 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_20_LC_1_11_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_20_LC_1_11_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_20_LC_1_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31515),
            .lcout(\pid_alt.error_i_regZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87173),
            .ce(N__33462),
            .sr(N__86036));
    defparam \pid_alt.error_i_reg_esr_3_LC_1_12_0 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_3_LC_1_12_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_3_LC_1_12_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_3_LC_1_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31506),
            .lcout(\pid_alt.error_i_regZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87187),
            .ce(N__33463),
            .sr(N__86035));
    defparam \pid_alt.error_i_reg_esr_4_LC_1_12_1 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_4_LC_1_12_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_4_LC_1_12_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_4_LC_1_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31497),
            .lcout(\pid_alt.error_i_regZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87187),
            .ce(N__33463),
            .sr(N__86035));
    defparam \pid_alt.error_i_reg_esr_5_LC_1_12_2 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_5_LC_1_12_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_5_LC_1_12_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_5_LC_1_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31491),
            .lcout(\pid_alt.error_i_regZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87187),
            .ce(N__33463),
            .sr(N__86035));
    defparam \pid_alt.error_i_reg_esr_10_LC_1_12_3 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_10_LC_1_12_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_10_LC_1_12_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_10_LC_1_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31485),
            .lcout(\pid_alt.error_i_regZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87187),
            .ce(N__33463),
            .sr(N__86035));
    defparam \pid_alt.error_i_reg_esr_0_LC_1_12_6 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_0_LC_1_12_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_0_LC_1_12_6 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \pid_alt.error_i_reg_esr_0_LC_1_12_6  (
            .in0(_gnd_net_),
            .in1(N__31647),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_i_regZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87187),
            .ce(N__33463),
            .sr(N__86035));
    defparam \pid_alt.error_p_reg_esr_0_LC_1_12_7 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_0_LC_1_12_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_0_LC_1_12_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_0_LC_1_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31638),
            .lcout(\pid_alt.error_p_regZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87187),
            .ce(N__33463),
            .sr(N__86035));
    defparam \pid_alt.error_i_reg_esr_1_LC_1_13_5 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_1_LC_1_13_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_1_LC_1_13_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_1_LC_1_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31620),
            .lcout(\pid_alt.error_i_regZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87204),
            .ce(N__33464),
            .sr(N__86034));
    defparam \pid_alt.error_d_reg_esr_0_LC_1_13_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_0_LC_1_13_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_0_LC_1_13_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_0_LC_1_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31608),
            .lcout(\pid_alt.error_d_regZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87204),
            .ce(N__33464),
            .sr(N__86034));
    defparam \pid_front.error_p_reg_esr_11_LC_1_14_0 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_11_LC_1_14_0 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_11_LC_1_14_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_p_reg_esr_11_LC_1_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31593),
            .lcout(\pid_front.error_p_regZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87221),
            .ce(N__86318),
            .sr(N__86033));
    defparam \pid_front.error_p_reg_esr_12_LC_1_14_1 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_12_LC_1_14_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_12_LC_1_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_p_reg_esr_12_LC_1_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31584),
            .lcout(\pid_front.error_p_regZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87221),
            .ce(N__86318),
            .sr(N__86033));
    defparam \pid_front.error_p_reg_esr_13_LC_1_14_2 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_13_LC_1_14_2 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_13_LC_1_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_p_reg_esr_13_LC_1_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31575),
            .lcout(\pid_front.error_p_regZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87221),
            .ce(N__86318),
            .sr(N__86033));
    defparam \pid_front.error_p_reg_esr_14_LC_1_14_3 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_14_LC_1_14_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_14_LC_1_14_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_front.error_p_reg_esr_14_LC_1_14_3  (
            .in0(N__31563),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_p_regZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87221),
            .ce(N__86318),
            .sr(N__86033));
    defparam \pid_front.error_p_reg_esr_15_LC_1_14_4 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_15_LC_1_14_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_15_LC_1_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_p_reg_esr_15_LC_1_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31554),
            .lcout(\pid_front.error_p_regZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87221),
            .ce(N__86318),
            .sr(N__86033));
    defparam \pid_front.error_p_reg_esr_16_LC_1_14_5 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_16_LC_1_14_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_16_LC_1_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_p_reg_esr_16_LC_1_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31719),
            .lcout(\pid_front.error_p_regZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87221),
            .ce(N__86318),
            .sr(N__86033));
    defparam \pid_front.error_p_reg_esr_7_LC_1_14_6 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_7_LC_1_14_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_7_LC_1_14_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_front.error_p_reg_esr_7_LC_1_14_6  (
            .in0(N__31710),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_p_regZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87221),
            .ce(N__86318),
            .sr(N__86033));
    defparam \pid_front.error_p_reg_esr_18_LC_1_14_7 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_18_LC_1_14_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_18_LC_1_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_p_reg_esr_18_LC_1_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31701),
            .lcout(\pid_front.error_p_regZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87221),
            .ce(N__86318),
            .sr(N__86033));
    defparam \pid_front.error_p_reg_esr_19_LC_1_15_0 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_19_LC_1_15_0 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_19_LC_1_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_p_reg_esr_19_LC_1_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31692),
            .lcout(\pid_front.error_p_regZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87236),
            .ce(N__86317),
            .sr(N__86032));
    defparam \pid_front.error_p_reg_esr_2_LC_1_15_1 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_2_LC_1_15_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_2_LC_1_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_p_reg_esr_2_LC_1_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31683),
            .lcout(\pid_front.error_p_regZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87236),
            .ce(N__86317),
            .sr(N__86032));
    defparam \pid_front.error_p_reg_esr_20_LC_1_15_2 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_20_LC_1_15_2 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_20_LC_1_15_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_p_reg_esr_20_LC_1_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31677),
            .lcout(\pid_front.error_p_regZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87236),
            .ce(N__86317),
            .sr(N__86032));
    defparam \pid_front.error_p_reg_esr_21_LC_1_15_3 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_21_LC_1_15_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_21_LC_1_15_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_p_reg_esr_21_LC_1_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31668),
            .lcout(\pid_front.error_p_regZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87236),
            .ce(N__86317),
            .sr(N__86032));
    defparam \pid_front.error_p_reg_esr_8_LC_1_15_4 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_8_LC_1_15_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_8_LC_1_15_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_p_reg_esr_8_LC_1_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31659),
            .lcout(\pid_front.error_p_regZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87236),
            .ce(N__86317),
            .sr(N__86032));
    defparam \pid_front.error_p_reg_esr_4_LC_1_15_5 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_4_LC_1_15_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_4_LC_1_15_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_p_reg_esr_4_LC_1_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31653),
            .lcout(\pid_front.error_p_regZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87236),
            .ce(N__86317),
            .sr(N__86032));
    defparam \pid_front.error_p_reg_esr_5_LC_1_15_6 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_5_LC_1_15_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_5_LC_1_15_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_p_reg_esr_5_LC_1_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31773),
            .lcout(\pid_front.error_p_regZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87236),
            .ce(N__86317),
            .sr(N__86032));
    defparam \pid_front.error_p_reg_esr_6_LC_1_15_7 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_6_LC_1_15_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_6_LC_1_15_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_p_reg_esr_6_LC_1_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31767),
            .lcout(\pid_front.error_p_regZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87236),
            .ce(N__86317),
            .sr(N__86032));
    defparam \pid_alt.error_d_reg_prev_esr_10_LC_1_16_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_10_LC_1_16_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_10_LC_1_16_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_10_LC_1_16_0  (
            .in0(N__31734),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87247),
            .ce(N__51493),
            .sr(N__79636));
    defparam \pid_alt.error_d_reg_prev_esr_RNIGDHM_0_11_LC_1_16_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIGDHM_0_11_LC_1_16_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIGDHM_0_11_LC_1_16_1 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIGDHM_0_11_LC_1_16_1  (
            .in0(N__31892),
            .in1(N__31853),
            .in2(_gnd_net_),
            .in3(N__31843),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIGDHM_0Z0Z_11 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNIGDHM_0Z0Z_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI1FP62_10_LC_1_16_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI1FP62_10_LC_1_16_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI1FP62_10_LC_1_16_2 .LUT_INIT=16'b1111101010100000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI1FP62_10_LC_1_16_2  (
            .in0(N__33362),
            .in1(_gnd_net_),
            .in2(N__31761),
            .in3(N__31758),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI1FP62Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIDAHM_10_LC_1_16_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIDAHM_10_LC_1_16_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIDAHM_10_LC_1_16_3 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIDAHM_10_LC_1_16_3  (
            .in0(N__31914),
            .in1(N__31743),
            .in2(_gnd_net_),
            .in3(N__31733),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIDAHMZ0Z_10 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNIDAHMZ0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNITPKD4_10_LC_1_16_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNITPKD4_10_LC_1_16_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNITPKD4_10_LC_1_16_4 .LUT_INIT=16'b1001011010010110;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNITPKD4_10_LC_1_16_4  (
            .in0(N__33361),
            .in1(N__31752),
            .in2(N__31746),
            .in3(N__34905),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNITPKD4Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIDAHM_0_10_LC_1_16_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIDAHM_0_10_LC_1_16_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIDAHM_0_10_LC_1_16_5 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIDAHM_0_10_LC_1_16_5  (
            .in0(N__31913),
            .in1(N__31742),
            .in2(_gnd_net_),
            .in3(N__31732),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIDAHM_0Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_11_LC_1_16_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_11_LC_1_16_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_11_LC_1_16_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_11_LC_1_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31845),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87247),
            .ce(N__51493),
            .sr(N__79636));
    defparam \pid_alt.error_d_reg_prev_esr_RNIGDHM_11_LC_1_16_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIGDHM_11_LC_1_16_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIGDHM_11_LC_1_16_7 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIGDHM_11_LC_1_16_7  (
            .in0(N__31893),
            .in1(N__31854),
            .in2(_gnd_net_),
            .in3(N__31844),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIGDHMZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI0J511_2_LC_1_17_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI0J511_2_LC_1_17_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI0J511_2_LC_1_17_0 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI0J511_2_LC_1_17_0  (
            .in0(N__32654),
            .in1(N__32541),
            .in2(_gnd_net_),
            .in3(N__32563),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI0J511Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_4_LC_1_18_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_4_LC_1_18_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_4_LC_1_18_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_4_LC_1_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32477),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87258),
            .ce(N__51487),
            .sr(N__79653));
    defparam \pid_alt.error_d_reg_prev_esr_18_LC_1_19_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_18_LC_1_19_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_18_LC_1_19_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_18_LC_1_19_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31797),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87262),
            .ce(N__51484),
            .sr(N__79662));
    defparam \pid_alt.error_d_reg_prev_esr_RNI86IM_0_19_LC_1_19_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI86IM_0_19_LC_1_19_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI86IM_0_19_LC_1_19_1 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI86IM_0_19_LC_1_19_1  (
            .in0(N__34820),
            .in1(N__34695),
            .in2(_gnd_net_),
            .in3(N__34721),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI86IM_0Z0Z_19 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNI86IM_0Z0Z_19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIOTT02_18_LC_1_19_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIOTT02_18_LC_1_19_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIOTT02_18_LC_1_19_2 .LUT_INIT=16'b1111101010100000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIOTT02_18_LC_1_19_2  (
            .in0(N__31824),
            .in1(_gnd_net_),
            .in2(N__31827),
            .in3(N__33578),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIOTT02Z0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI53IM_18_LC_1_19_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI53IM_18_LC_1_19_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI53IM_18_LC_1_19_3 .LUT_INIT=16'b1010111100001010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI53IM_18_LC_1_19_3  (
            .in0(N__31796),
            .in1(_gnd_net_),
            .in2(N__31809),
            .in3(N__32025),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI53IMZ0Z_18 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNI53IMZ0Z_18_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI8IQ14_18_LC_1_19_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI8IQ14_18_LC_1_19_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI8IQ14_18_LC_1_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI8IQ14_18_LC_1_19_4  (
            .in0(N__34610),
            .in1(N__31818),
            .in2(N__31812),
            .in3(N__33577),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI8IQ14Z0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIGKS02_17_LC_1_19_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIGKS02_17_LC_1_19_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIGKS02_17_LC_1_19_5 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIGKS02_17_LC_1_19_5  (
            .in0(N__31977),
            .in1(N__31881),
            .in2(_gnd_net_),
            .in3(N__33341),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIGKS02Z0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI53IM_0_18_LC_1_19_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI53IM_0_18_LC_1_19_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI53IM_0_18_LC_1_19_6 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI53IM_0_18_LC_1_19_6  (
            .in0(N__32024),
            .in1(N__31805),
            .in2(_gnd_net_),
            .in3(N__31795),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI53IM_0Z0Z_18 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNI53IM_0Z0Z_18_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIOVN14_17_LC_1_19_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIOVN14_17_LC_1_19_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIOVN14_17_LC_1_19_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIOVN14_17_LC_1_19_7  (
            .in0(N__31976),
            .in1(N__34877),
            .in2(N__31875),
            .in3(N__33340),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIOVN14Z0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_8_LC_1_20_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_8_LC_1_20_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_8_LC_1_20_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_8_LC_1_20_0  (
            .in0(N__32718),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87266),
            .ce(N__51481),
            .sr(N__79669));
    defparam \pid_alt.error_d_reg_prev_esr_RNII5611_8_LC_1_20_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNII5611_8_LC_1_20_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNII5611_8_LC_1_20_1 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNII5611_8_LC_1_20_1  (
            .in0(N__33540),
            .in1(N__32687),
            .in2(_gnd_net_),
            .in3(N__32717),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNII5611Z0Z_8 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNII5611Z0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIG75T2_8_LC_1_20_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIG75T2_8_LC_1_20_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIG75T2_8_LC_1_20_2 .LUT_INIT=16'b1111110011000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIG75T2_8_LC_1_20_2  (
            .in0(_gnd_net_),
            .in1(N__33035),
            .in2(N__31872),
            .in3(N__31869),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIG75T2Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIL8611_0_9_LC_1_20_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIL8611_0_9_LC_1_20_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIL8611_0_9_LC_1_20_3 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIL8611_0_9_LC_1_20_3  (
            .in0(N__35018),
            .in1(N__34997),
            .in2(_gnd_net_),
            .in3(N__34981),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIL8611_0Z0Z_9 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNIL8611_0Z0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIN49Q5_8_LC_1_20_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIN49Q5_8_LC_1_20_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIN49Q5_8_LC_1_20_4 .LUT_INIT=16'b1001011010010110;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIN49Q5_8_LC_1_20_4  (
            .in0(N__31863),
            .in1(N__33034),
            .in2(N__31857),
            .in3(N__34497),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIN49Q5Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_9_LC_1_20_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_9_LC_1_20_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_9_LC_1_20_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_9_LC_1_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34982),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87266),
            .ce(N__51481),
            .sr(N__79669));
    defparam \pid_alt.error_i_acumm_prereg_esr_9_LC_1_20_6 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_9_LC_1_20_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_9_LC_1_20_6 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_9_LC_1_20_6  (
            .in0(_gnd_net_),
            .in1(N__33036),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87266),
            .ce(N__51481),
            .sr(N__79669));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIPNRC1_11_LC_1_20_7 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIPNRC1_11_LC_1_20_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIPNRC1_11_LC_1_20_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNIPNRC1_11_LC_1_20_7  (
            .in0(N__39398),
            .in1(N__39504),
            .in2(N__39052),
            .in3(N__39605),
            .lcout(\pid_alt.m21_e_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_p_reg_esr_2_LC_1_21_1 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_2_LC_1_21_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_2_LC_1_21_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_2_LC_1_21_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31986),
            .lcout(\pid_alt.error_p_regZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87270),
            .ce(N__33465),
            .sr(N__86030));
    defparam \pid_alt.error_d_reg_prev_esr_RNI20IM_17_LC_1_21_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI20IM_17_LC_1_21_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI20IM_17_LC_1_21_3 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI20IM_17_LC_1_21_3  (
            .in0(N__33375),
            .in1(N__33285),
            .in2(_gnd_net_),
            .in3(N__33316),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI20IMZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_p_reg_esr_17_LC_1_21_4 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_17_LC_1_21_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_17_LC_1_21_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_17_LC_1_21_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31965),
            .lcout(\pid_alt.error_p_regZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87270),
            .ce(N__33465),
            .sr(N__86030));
    defparam \pid_alt.error_d_reg_prev_esr_RNI6P511_4_LC_1_21_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI6P511_4_LC_1_21_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI6P511_4_LC_1_21_6 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI6P511_4_LC_1_21_6  (
            .in0(N__32513),
            .in1(N__32498),
            .in2(_gnd_net_),
            .in3(N__32476),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI6P511Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_p_reg_esr_4_LC_1_21_7 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_4_LC_1_21_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_4_LC_1_21_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_4_LC_1_21_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31953),
            .lcout(\pid_alt.error_p_regZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87270),
            .ce(N__33465),
            .sr(N__86030));
    defparam \pid_alt.error_p_reg_esr_20_LC_1_22_1 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_20_LC_1_22_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_20_LC_1_22_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_20_LC_1_22_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31944),
            .lcout(\pid_alt.error_p_regZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87275),
            .ce(N__33466),
            .sr(N__86029));
    defparam \pid_alt.error_p_reg_esr_12_LC_1_22_3 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_12_LC_1_22_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_12_LC_1_22_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_12_LC_1_22_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31932),
            .lcout(\pid_alt.error_p_regZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87275),
            .ce(N__33466),
            .sr(N__86029));
    defparam \pid_alt.error_p_reg_esr_10_LC_1_22_4 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_10_LC_1_22_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_10_LC_1_22_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_10_LC_1_22_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31923),
            .lcout(\pid_alt.error_p_regZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87275),
            .ce(N__33466),
            .sr(N__86029));
    defparam \pid_alt.error_p_reg_esr_11_LC_1_22_5 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_11_LC_1_22_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_11_LC_1_22_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_11_LC_1_22_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31902),
            .lcout(\pid_alt.error_p_regZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87275),
            .ce(N__33466),
            .sr(N__86029));
    defparam \pid_alt.error_p_reg_esr_15_LC_1_22_6 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_15_LC_1_22_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_15_LC_1_22_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_15_LC_1_22_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32070),
            .lcout(\pid_alt.error_p_regZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87275),
            .ce(N__33466),
            .sr(N__86029));
    defparam \pid_alt.error_p_reg_esr_9_LC_1_22_7 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_9_LC_1_22_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_9_LC_1_22_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_9_LC_1_22_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32061),
            .lcout(\pid_alt.error_p_regZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87275),
            .ce(N__33466),
            .sr(N__86029));
    defparam \pid_alt.error_p_reg_esr_13_LC_1_23_0 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_13_LC_1_23_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_13_LC_1_23_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_13_LC_1_23_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32052),
            .lcout(\pid_alt.error_p_regZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87278),
            .ce(N__33468),
            .sr(N__86027));
    defparam \pid_alt.error_p_reg_esr_14_LC_1_23_1 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_14_LC_1_23_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_14_LC_1_23_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_14_LC_1_23_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32043),
            .lcout(\pid_alt.error_p_regZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87278),
            .ce(N__33468),
            .sr(N__86027));
    defparam \pid_alt.error_p_reg_esr_18_LC_1_23_2 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_18_LC_1_23_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_18_LC_1_23_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_18_LC_1_23_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32034),
            .lcout(\pid_alt.error_p_regZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87278),
            .ce(N__33468),
            .sr(N__86027));
    defparam \pid_alt.error_p_reg_esr_5_LC_1_23_3 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_5_LC_1_23_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_5_LC_1_23_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_p_reg_esr_5_LC_1_23_3  (
            .in0(N__32013),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_p_regZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87278),
            .ce(N__33468),
            .sr(N__86027));
    defparam \pid_alt.error_p_reg_esr_6_LC_1_23_4 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_6_LC_1_23_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_6_LC_1_23_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_6_LC_1_23_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32007),
            .lcout(\pid_alt.error_p_regZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87278),
            .ce(N__33468),
            .sr(N__86027));
    defparam \pid_alt.error_p_reg_esr_7_LC_1_23_5 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_7_LC_1_23_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_7_LC_1_23_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_7_LC_1_23_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32001),
            .lcout(\pid_alt.error_p_regZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87278),
            .ce(N__33468),
            .sr(N__86027));
    defparam \pid_alt.error_p_reg_esr_19_LC_1_23_6 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_19_LC_1_23_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_19_LC_1_23_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_19_LC_1_23_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31995),
            .lcout(\pid_alt.error_p_regZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87278),
            .ce(N__33468),
            .sr(N__86027));
    defparam \pid_alt.error_p_reg_esr_16_LC_1_23_7 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_16_LC_1_23_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_16_LC_1_23_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_16_LC_1_23_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32178),
            .lcout(\pid_alt.error_p_regZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87278),
            .ce(N__33468),
            .sr(N__86027));
    defparam \pid_alt.error_d_reg_esr_12_LC_2_5_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_12_LC_2_5_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_12_LC_2_5_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_12_LC_2_5_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32169),
            .lcout(\pid_alt.error_d_regZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87071),
            .ce(N__33455),
            .sr(N__86042));
    defparam \Commands_frame_decoder.source_alt_kd_1_LC_2_7_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kd_1_LC_2_7_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kd_1_LC_2_7_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_kd_1_LC_2_7_1  (
            .in0(_gnd_net_),
            .in1(N__84182),
            .in2(_gnd_net_),
            .in3(N__86186),
            .lcout(alt_kd_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87099),
            .ce(N__33404),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kd_4_LC_2_7_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kd_4_LC_2_7_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kd_4_LC_2_7_2 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Commands_frame_decoder.source_alt_kd_4_LC_2_7_2  (
            .in0(N__86188),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85009),
            .lcout(alt_kd_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87099),
            .ce(N__33404),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kd_3_LC_2_7_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kd_3_LC_2_7_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kd_3_LC_2_7_3 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_kd_3_LC_2_7_3  (
            .in0(_gnd_net_),
            .in1(N__84001),
            .in2(_gnd_net_),
            .in3(N__86187),
            .lcout(alt_kd_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87099),
            .ce(N__33404),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kd_5_LC_2_7_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kd_5_LC_2_7_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kd_5_LC_2_7_5 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_kd_5_LC_2_7_5  (
            .in0(_gnd_net_),
            .in1(N__85177),
            .in2(_gnd_net_),
            .in3(N__86189),
            .lcout(alt_kd_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87099),
            .ce(N__33404),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kd_6_LC_2_7_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kd_6_LC_2_7_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kd_6_LC_2_7_7 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_kd_6_LC_2_7_7  (
            .in0(_gnd_net_),
            .in1(N__73628),
            .in2(_gnd_net_),
            .in3(N__86190),
            .lcout(alt_kd_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87099),
            .ce(N__33404),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kd_2_LC_2_8_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kd_2_LC_2_8_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kd_2_LC_2_8_5 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_kd_2_LC_2_8_5  (
            .in0(_gnd_net_),
            .in1(N__77548),
            .in2(_gnd_net_),
            .in3(N__86183),
            .lcout(alt_kd_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87114),
            .ce(N__33403),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kd_7_LC_2_8_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kd_7_LC_2_8_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kd_7_LC_2_8_6 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Commands_frame_decoder.source_alt_kd_7_LC_2_8_6  (
            .in0(N__86184),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85379),
            .lcout(alt_kd_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87114),
            .ce(N__33403),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.WDT_0_LC_2_9_0 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_0_LC_2_9_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_0_LC_2_9_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_0_LC_2_9_0  (
            .in0(_gnd_net_),
            .in1(N__32226),
            .in2(N__33660),
            .in3(N__33659),
            .lcout(\Commands_frame_decoder.WDTZ0Z_0 ),
            .ltout(),
            .carryin(bfn_2_9_0_),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_0 ),
            .clk(N__87130),
            .ce(),
            .sr(N__34032));
    defparam \Commands_frame_decoder.WDT_1_LC_2_9_1 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_1_LC_2_9_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_1_LC_2_9_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_1_LC_2_9_1  (
            .in0(_gnd_net_),
            .in1(N__32220),
            .in2(_gnd_net_),
            .in3(N__32214),
            .lcout(\Commands_frame_decoder.WDTZ0Z_1 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_0 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_1 ),
            .clk(N__87130),
            .ce(),
            .sr(N__34032));
    defparam \Commands_frame_decoder.WDT_2_LC_2_9_2 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_2_LC_2_9_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_2_LC_2_9_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_2_LC_2_9_2  (
            .in0(_gnd_net_),
            .in1(N__32211),
            .in2(_gnd_net_),
            .in3(N__32205),
            .lcout(\Commands_frame_decoder.WDTZ0Z_2 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_1 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_2 ),
            .clk(N__87130),
            .ce(),
            .sr(N__34032));
    defparam \Commands_frame_decoder.WDT_3_LC_2_9_3 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_3_LC_2_9_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_3_LC_2_9_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_3_LC_2_9_3  (
            .in0(_gnd_net_),
            .in1(N__32202),
            .in2(_gnd_net_),
            .in3(N__32196),
            .lcout(\Commands_frame_decoder.WDTZ0Z_3 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_2 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_3 ),
            .clk(N__87130),
            .ce(),
            .sr(N__34032));
    defparam \Commands_frame_decoder.WDT_4_LC_2_9_4 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_4_LC_2_9_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_4_LC_2_9_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_4_LC_2_9_4  (
            .in0(_gnd_net_),
            .in1(N__33747),
            .in2(_gnd_net_),
            .in3(N__32193),
            .lcout(\Commands_frame_decoder.WDTZ0Z_4 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_3 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_4 ),
            .clk(N__87130),
            .ce(),
            .sr(N__34032));
    defparam \Commands_frame_decoder.WDT_5_LC_2_9_5 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_5_LC_2_9_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_5_LC_2_9_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_5_LC_2_9_5  (
            .in0(_gnd_net_),
            .in1(N__33789),
            .in2(_gnd_net_),
            .in3(N__32190),
            .lcout(\Commands_frame_decoder.WDTZ0Z_5 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_4 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_5 ),
            .clk(N__87130),
            .ce(),
            .sr(N__34032));
    defparam \Commands_frame_decoder.WDT_6_LC_2_9_6 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_6_LC_2_9_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_6_LC_2_9_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_6_LC_2_9_6  (
            .in0(_gnd_net_),
            .in1(N__33807),
            .in2(_gnd_net_),
            .in3(N__32187),
            .lcout(\Commands_frame_decoder.WDTZ0Z_6 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_5 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_6 ),
            .clk(N__87130),
            .ce(),
            .sr(N__34032));
    defparam \Commands_frame_decoder.WDT_7_LC_2_9_7 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_7_LC_2_9_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_7_LC_2_9_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_7_LC_2_9_7  (
            .in0(_gnd_net_),
            .in1(N__33769),
            .in2(_gnd_net_),
            .in3(N__32184),
            .lcout(\Commands_frame_decoder.WDTZ0Z_7 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_6 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_7 ),
            .clk(N__87130),
            .ce(),
            .sr(N__34032));
    defparam \Commands_frame_decoder.WDT_8_LC_2_10_0 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_8_LC_2_10_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_8_LC_2_10_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_8_LC_2_10_0  (
            .in0(_gnd_net_),
            .in1(N__33627),
            .in2(_gnd_net_),
            .in3(N__32181),
            .lcout(\Commands_frame_decoder.WDTZ0Z_8 ),
            .ltout(),
            .carryin(bfn_2_10_0_),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_8 ),
            .clk(N__87147),
            .ce(),
            .sr(N__34025));
    defparam \Commands_frame_decoder.WDT_9_LC_2_10_1 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_9_LC_2_10_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_9_LC_2_10_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_9_LC_2_10_1  (
            .in0(_gnd_net_),
            .in1(N__33609),
            .in2(_gnd_net_),
            .in3(N__32265),
            .lcout(\Commands_frame_decoder.WDTZ0Z_9 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_8 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_9 ),
            .clk(N__87147),
            .ce(),
            .sr(N__34025));
    defparam \Commands_frame_decoder.WDT_10_LC_2_10_2 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_10_LC_2_10_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_10_LC_2_10_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_10_LC_2_10_2  (
            .in0(_gnd_net_),
            .in1(N__33891),
            .in2(_gnd_net_),
            .in3(N__32262),
            .lcout(\Commands_frame_decoder.WDTZ0Z_10 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_9 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_10 ),
            .clk(N__87147),
            .ce(),
            .sr(N__34025));
    defparam \Commands_frame_decoder.WDT_11_LC_2_10_3 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_11_LC_2_10_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_11_LC_2_10_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_11_LC_2_10_3  (
            .in0(_gnd_net_),
            .in1(N__33828),
            .in2(_gnd_net_),
            .in3(N__32259),
            .lcout(\Commands_frame_decoder.WDTZ0Z_11 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_10 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_11 ),
            .clk(N__87147),
            .ce(),
            .sr(N__34025));
    defparam \Commands_frame_decoder.WDT_12_LC_2_10_4 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_12_LC_2_10_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_12_LC_2_10_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_12_LC_2_10_4  (
            .in0(_gnd_net_),
            .in1(N__33851),
            .in2(_gnd_net_),
            .in3(N__32256),
            .lcout(\Commands_frame_decoder.WDTZ0Z_12 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_11 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_12 ),
            .clk(N__87147),
            .ce(),
            .sr(N__34025));
    defparam \Commands_frame_decoder.WDT_13_LC_2_10_5 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_13_LC_2_10_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_13_LC_2_10_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_13_LC_2_10_5  (
            .in0(_gnd_net_),
            .in1(N__33873),
            .in2(_gnd_net_),
            .in3(N__32253),
            .lcout(\Commands_frame_decoder.WDTZ0Z_13 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_12 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_13 ),
            .clk(N__87147),
            .ce(),
            .sr(N__34025));
    defparam \Commands_frame_decoder.WDT_14_LC_2_10_6 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_14_LC_2_10_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_14_LC_2_10_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_14_LC_2_10_6  (
            .in0(_gnd_net_),
            .in1(N__34163),
            .in2(_gnd_net_),
            .in3(N__32250),
            .lcout(\Commands_frame_decoder.WDTZ0Z_14 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_13 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_14 ),
            .clk(N__87147),
            .ce(),
            .sr(N__34025));
    defparam \Commands_frame_decoder.WDT_15_LC_2_10_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.WDT_15_LC_2_10_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_15_LC_2_10_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \Commands_frame_decoder.WDT_15_LC_2_10_7  (
            .in0(_gnd_net_),
            .in1(N__34133),
            .in2(_gnd_net_),
            .in3(N__32247),
            .lcout(\Commands_frame_decoder.WDTZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87147),
            .ce(),
            .sr(N__34025));
    defparam \Commands_frame_decoder.source_alt_ki_0_LC_2_11_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_ki_0_LC_2_11_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_ki_0_LC_2_11_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_ki_0_LC_2_11_0  (
            .in0(_gnd_net_),
            .in1(N__83795),
            .in2(_gnd_net_),
            .in3(N__86175),
            .lcout(alt_ki_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87163),
            .ce(N__33705),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_ki_1_LC_2_11_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_ki_1_LC_2_11_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_ki_1_LC_2_11_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Commands_frame_decoder.source_alt_ki_1_LC_2_11_1  (
            .in0(N__86176),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84156),
            .lcout(alt_ki_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87163),
            .ce(N__33705),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_ki_2_LC_2_11_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_ki_2_LC_2_11_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_ki_2_LC_2_11_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_ki_2_LC_2_11_2  (
            .in0(_gnd_net_),
            .in1(N__77546),
            .in2(_gnd_net_),
            .in3(N__86177),
            .lcout(alt_ki_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87163),
            .ce(N__33705),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_ki_3_LC_2_11_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_ki_3_LC_2_11_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_ki_3_LC_2_11_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Commands_frame_decoder.source_alt_ki_3_LC_2_11_3  (
            .in0(N__86178),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__83980),
            .lcout(alt_ki_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87163),
            .ce(N__33705),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_ki_4_LC_2_11_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_ki_4_LC_2_11_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_ki_4_LC_2_11_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_ki_4_LC_2_11_4  (
            .in0(_gnd_net_),
            .in1(N__84960),
            .in2(_gnd_net_),
            .in3(N__86179),
            .lcout(alt_ki_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87163),
            .ce(N__33705),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_ki_5_LC_2_11_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_ki_5_LC_2_11_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_ki_5_LC_2_11_5 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Commands_frame_decoder.source_alt_ki_5_LC_2_11_5  (
            .in0(N__86180),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85168),
            .lcout(alt_ki_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87163),
            .ce(N__33705),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_ki_6_LC_2_11_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_ki_6_LC_2_11_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_ki_6_LC_2_11_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_ki_6_LC_2_11_6  (
            .in0(_gnd_net_),
            .in1(N__73605),
            .in2(_gnd_net_),
            .in3(N__86181),
            .lcout(alt_ki_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87163),
            .ce(N__33705),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_ki_7_LC_2_11_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_ki_7_LC_2_11_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_ki_7_LC_2_11_7 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Commands_frame_decoder.source_alt_ki_7_LC_2_11_7  (
            .in0(N__86182),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85356),
            .lcout(alt_ki_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87163),
            .ce(N__33705),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNO_1_1_LC_2_12_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNO_1_1_LC_2_12_0 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNO_1_1_LC_2_12_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Commands_frame_decoder.state_RNO_1_1_LC_2_12_0  (
            .in0(_gnd_net_),
            .in1(N__85357),
            .in2(_gnd_net_),
            .in3(N__83769),
            .lcout(),
            .ltout(\Commands_frame_decoder.state_ns_0_a3_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNO_0_1_LC_2_12_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNO_0_1_LC_2_12_1 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNO_0_1_LC_2_12_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Commands_frame_decoder.state_RNO_0_1_LC_2_12_1  (
            .in0(N__33965),
            .in1(N__85132),
            .in2(N__32271),
            .in3(N__77510),
            .lcout(\Commands_frame_decoder.state_ns_0_a3_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_ns_i_a2_2_1_0_LC_2_12_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_ns_i_a2_2_1_0_LC_2_12_2 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_ns_i_a2_2_1_0_LC_2_12_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \Commands_frame_decoder.state_ns_i_a2_2_1_0_LC_2_12_2  (
            .in0(N__73563),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__83945),
            .lcout(),
            .ltout(\Commands_frame_decoder.state_ns_i_a2_2_1Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_ns_i_a2_2_0_LC_2_12_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_ns_i_a2_2_0_LC_2_12_3 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_ns_i_a2_2_0_LC_2_12_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Commands_frame_decoder.state_ns_i_a2_2_0_LC_2_12_3  (
            .in0(N__84124),
            .in1(N__38398),
            .in2(N__32268),
            .in3(N__84936),
            .lcout(\Commands_frame_decoder.N_410 ),
            .ltout(\Commands_frame_decoder.N_410_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNO_1_0_LC_2_12_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNO_1_0_LC_2_12_4 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNO_1_0_LC_2_12_4 .LUT_INIT=16'b1111000010000000;
    LogicCell40 \Commands_frame_decoder.state_RNO_1_0_LC_2_12_4  (
            .in0(N__36012),
            .in1(N__33999),
            .in2(N__32391),
            .in3(N__34184),
            .lcout(\Commands_frame_decoder.N_371 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_xy_kp_4_LC_2_13_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_kp_4_LC_2_13_0 .SEQ_MODE=4'b1001;
    defparam \Commands_frame_decoder.source_xy_kp_4_LC_2_13_0 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \Commands_frame_decoder.source_xy_kp_4_LC_2_13_0  (
            .in0(N__38443),
            .in1(N__32371),
            .in2(N__34059),
            .in3(N__84987),
            .lcout(xy_kp_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87191),
            .ce(),
            .sr(N__79607));
    defparam \Commands_frame_decoder.state_RNIRSI31_11_LC_2_13_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIRSI31_11_LC_2_13_1 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIRSI31_11_LC_2_13_1 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \Commands_frame_decoder.state_RNIRSI31_11_LC_2_13_1  (
            .in0(N__34096),
            .in1(N__38442),
            .in2(_gnd_net_),
            .in3(N__79960),
            .lcout(\Commands_frame_decoder.state_RNIRSI31Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNIGK1J_4_LC_2_13_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIGK1J_4_LC_2_13_3 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIGK1J_4_LC_2_13_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Commands_frame_decoder.state_RNIGK1J_4_LC_2_13_3  (
            .in0(_gnd_net_),
            .in1(N__38313),
            .in2(_gnd_net_),
            .in3(N__38439),
            .lcout(\Commands_frame_decoder.source_CH3data_1_sqmuxa ),
            .ltout(\Commands_frame_decoder.source_CH3data_1_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_5_LC_2_13_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_5_LC_2_13_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_5_LC_2_13_4 .LUT_INIT=16'b1111101011110000;
    LogicCell40 \Commands_frame_decoder.state_5_LC_2_13_4  (
            .in0(N__32346),
            .in1(_gnd_net_),
            .in2(N__32349),
            .in3(N__39291),
            .lcout(\Commands_frame_decoder.stateZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87191),
            .ce(),
            .sr(N__79607));
    defparam \Commands_frame_decoder.state_RNIHL1J_5_LC_2_13_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIHL1J_5_LC_2_13_5 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIHL1J_5_LC_2_13_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Commands_frame_decoder.state_RNIHL1J_5_LC_2_13_5  (
            .in0(_gnd_net_),
            .in1(N__32345),
            .in2(_gnd_net_),
            .in3(N__38440),
            .lcout(\Commands_frame_decoder.source_CH4data_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNILP1J_9_LC_2_13_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNILP1J_9_LC_2_13_7 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNILP1J_9_LC_2_13_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Commands_frame_decoder.state_RNILP1J_9_LC_2_13_7  (
            .in0(_gnd_net_),
            .in1(N__34070),
            .in2(_gnd_net_),
            .in3(N__38441),
            .lcout(\Commands_frame_decoder.source_offset4data_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNICV511_6_LC_2_14_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNICV511_6_LC_2_14_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNICV511_6_LC_2_14_0 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNICV511_6_LC_2_14_0  (
            .in0(N__35979),
            .in1(N__35951),
            .in2(_gnd_net_),
            .in3(N__35935),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNICV511Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_p_reg_esr_RNIOI4P_0_LC_2_14_1 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_RNIOI4P_0_LC_2_14_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_p_reg_esr_RNIOI4P_0_LC_2_14_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \pid_alt.error_p_reg_esr_RNIOI4P_0_LC_2_14_1  (
            .in0(_gnd_net_),
            .in1(N__32411),
            .in2(_gnd_net_),
            .in3(N__32425),
            .lcout(\pid_alt.error_p_reg_esr_RNIOI4PZ0Z_0 ),
            .ltout(\pid_alt.error_p_reg_esr_RNIOI4PZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIFPN33_1_LC_2_14_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIFPN33_1_LC_2_14_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIFPN33_1_LC_2_14_2 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIFPN33_1_LC_2_14_2  (
            .in0(N__36871),
            .in1(_gnd_net_),
            .in2(N__32436),
            .in3(N__32576),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIFPN33Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_6_LC_2_14_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_6_LC_2_14_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_6_LC_2_14_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_6_LC_2_14_3  (
            .in0(N__35936),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87208),
            .ce(N__51495),
            .sr(N__79613));
    defparam \pid_alt.error_d_reg_prev_esr_0_LC_2_14_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_0_LC_2_14_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_0_LC_2_14_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_0_LC_2_14_4  (
            .in0(N__32427),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87208),
            .ce(N__51495),
            .sr(N__79613));
    defparam \pid_alt.error_d_reg_prev_esr_RNI2Q08_0_LC_2_14_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI2Q08_0_LC_2_14_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI2Q08_0_LC_2_14_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI2Q08_0_LC_2_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32433),
            .lcout(\pid_alt.error_d_reg_prev_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_p_reg_esr_RNI3SMI1_0_LC_2_14_6 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_RNI3SMI1_0_LC_2_14_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_p_reg_esr_RNI3SMI1_0_LC_2_14_6 .LUT_INIT=16'b1010010110100101;
    LogicCell40 \pid_alt.error_p_reg_esr_RNI3SMI1_0_LC_2_14_6  (
            .in0(N__32426),
            .in1(_gnd_net_),
            .in2(N__32415),
            .in3(N__34238),
            .lcout(\pid_alt.error_p_reg_esr_RNI3SMI1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIMJHM_13_LC_2_14_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIMJHM_13_LC_2_14_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIMJHM_13_LC_2_14_7 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIMJHM_13_LC_2_14_7  (
            .in0(N__38784),
            .in1(N__38760),
            .in2(_gnd_net_),
            .in3(N__38729),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIMJHMZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNITF511_1_LC_2_15_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNITF511_1_LC_2_15_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNITF511_1_LC_2_15_0 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNITF511_1_LC_2_15_0  (
            .in0(N__33508),
            .in1(N__32605),
            .in2(_gnd_net_),
            .in3(N__32625),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNITF511Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_1_LC_2_15_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_1_LC_2_15_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_1_LC_2_15_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_1_LC_2_15_1  (
            .in0(N__32628),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87223),
            .ce(N__51494),
            .sr(N__79621));
    defparam \pid_alt.error_d_reg_prev_esr_RNITF511_0_1_LC_2_15_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNITF511_0_1_LC_2_15_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNITF511_0_1_LC_2_15_2 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNITF511_0_1_LC_2_15_2  (
            .in0(N__33509),
            .in1(N__32606),
            .in2(_gnd_net_),
            .in3(N__32626),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNITF511_0Z0Z_1 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNITF511_0Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNII5LS3_1_LC_2_15_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNII5LS3_1_LC_2_15_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNII5LS3_1_LC_2_15_3 .LUT_INIT=16'b1110100010001000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNII5LS3_1_LC_2_15_3  (
            .in0(N__32634),
            .in1(N__32400),
            .in2(N__32394),
            .in3(N__32588),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNII5LS3Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI0J511_0_2_LC_2_15_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI0J511_0_2_LC_2_15_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI0J511_0_2_LC_2_15_4 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI0J511_0_2_LC_2_15_4  (
            .in0(N__32655),
            .in1(N__32537),
            .in2(_gnd_net_),
            .in3(N__32564),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI0J511_0Z0Z_2 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNI0J511_0Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIT2B22_1_LC_2_15_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIT2B22_1_LC_2_15_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIT2B22_1_LC_2_15_5 .LUT_INIT=16'b0100101111010010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIT2B22_1_LC_2_15_5  (
            .in0(N__32627),
            .in1(N__32607),
            .in2(N__32592),
            .in3(N__33510),
            .lcout(),
            .ltout(\pid_alt.un1_pid_prereg_16_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIF0465_1_LC_2_15_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIF0465_1_LC_2_15_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIF0465_1_LC_2_15_6 .LUT_INIT=16'b0101101011110000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIF0465_1_LC_2_15_6  (
            .in0(N__32589),
            .in1(N__35212),
            .in2(N__32580),
            .in3(N__32577),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIF0465Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_2_LC_2_15_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_2_LC_2_15_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_2_LC_2_15_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_2_LC_2_15_7  (
            .in0(N__32565),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87223),
            .ce(N__51494),
            .sr(N__79621));
    defparam \pid_alt.error_d_reg_prev_esr_RNI11TA9_3_LC_2_16_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI11TA9_3_LC_2_16_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI11TA9_3_LC_2_16_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI11TA9_3_LC_2_16_0  (
            .in0(N__32444),
            .in1(N__32526),
            .in2(N__34371),
            .in3(N__35233),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI11TA9Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI3M511_3_LC_2_16_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI3M511_3_LC_2_16_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI3M511_3_LC_2_16_1 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI3M511_3_LC_2_16_1  (
            .in0(N__33482),
            .in1(N__32753),
            .in2(_gnd_net_),
            .in3(N__32776),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI3M511Z0Z_3 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNI3M511Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNICISB3_3_LC_2_16_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNICISB3_3_LC_2_16_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNICISB3_3_LC_2_16_2 .LUT_INIT=16'b1111101010100000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNICISB3_3_LC_2_16_2  (
            .in0(N__32445),
            .in1(_gnd_net_),
            .in2(N__32520),
            .in3(N__35234),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNICISB3Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI6P511_0_4_LC_2_16_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI6P511_0_4_LC_2_16_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI6P511_0_4_LC_2_16_3 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI6P511_0_4_LC_2_16_3  (
            .in0(N__32517),
            .in1(N__32499),
            .in2(_gnd_net_),
            .in3(N__32478),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI6P511_0Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_3_LC_2_16_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_3_LC_2_16_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_3_LC_2_16_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_3_LC_2_16_4  (
            .in0(N__32778),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87238),
            .ce(N__51491),
            .sr(N__79629));
    defparam \pid_alt.error_d_reg_prev_esr_RNILE0V5_2_LC_2_16_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNILE0V5_2_LC_2_16_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNILE0V5_2_LC_2_16_5 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNILE0V5_2_LC_2_16_5  (
            .in0(N__32745),
            .in1(N__32739),
            .in2(_gnd_net_),
            .in3(N__32727),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNILE0V5Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI3M511_0_3_LC_2_16_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI3M511_0_3_LC_2_16_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI3M511_0_3_LC_2_16_6 .LUT_INIT=16'b0101101010100101;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI3M511_0_3_LC_2_16_6  (
            .in0(N__32777),
            .in1(_gnd_net_),
            .in2(N__32757),
            .in3(N__33483),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI3M511_0Z0Z_3 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNI3M511_0Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNILDG87_2_LC_2_16_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNILDG87_2_LC_2_16_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNILDG87_2_LC_2_16_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNILDG87_2_LC_2_16_7  (
            .in0(N__35413),
            .in1(N__32738),
            .in2(N__32730),
            .in3(N__32726),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNILDG87Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_7_LC_2_17_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_7_LC_2_17_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_7_LC_2_17_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_7_LC_2_17_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32916),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87249),
            .ce(N__51488),
            .sr(N__79637));
    defparam \pid_alt.error_d_reg_prev_esr_RNII5611_0_8_LC_2_17_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNII5611_0_8_LC_2_17_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNII5611_0_8_LC_2_17_1 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNII5611_0_8_LC_2_17_1  (
            .in0(N__32711),
            .in1(N__33536),
            .in2(_gnd_net_),
            .in3(N__32691),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNII5611_0Z0Z_8 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNII5611_0Z0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI7T3T2_7_LC_2_17_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI7T3T2_7_LC_2_17_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI7T3T2_7_LC_2_17_2 .LUT_INIT=16'b1111110011000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI7T3T2_7_LC_2_17_2  (
            .in0(_gnd_net_),
            .in1(N__32670),
            .in2(N__32673),
            .in3(N__37172),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI7T3T2Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIF2611_7_LC_2_17_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIF2611_7_LC_2_17_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIF2611_7_LC_2_17_3 .LUT_INIT=16'b1010111100001010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIF2611_7_LC_2_17_3  (
            .in0(N__32915),
            .in1(_gnd_net_),
            .in2(N__32928),
            .in3(N__32943),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIF2611Z0Z_7 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNIF2611Z0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI5G6Q5_7_LC_2_17_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI5G6Q5_7_LC_2_17_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI5G6Q5_7_LC_2_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI5G6Q5_7_LC_2_17_4  (
            .in0(N__34319),
            .in1(N__32664),
            .in2(N__32658),
            .in3(N__37171),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI5G6Q5Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIUI2T2_6_LC_2_17_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIUI2T2_6_LC_2_17_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIUI2T2_6_LC_2_17_5 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIUI2T2_6_LC_2_17_5  (
            .in0(N__32889),
            .in1(N__32895),
            .in2(_gnd_net_),
            .in3(N__34511),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIUI2T2Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIF2611_0_7_LC_2_17_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIF2611_0_7_LC_2_17_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIF2611_0_7_LC_2_17_6 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIF2611_0_7_LC_2_17_6  (
            .in0(N__32942),
            .in1(N__32924),
            .in2(_gnd_net_),
            .in3(N__32914),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIF2611_0Z0Z_7 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNIF2611_0Z0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIJR3Q5_6_LC_2_17_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIJR3Q5_6_LC_2_17_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIJR3Q5_6_LC_2_17_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIJR3Q5_6_LC_2_17_7  (
            .in0(N__32888),
            .in1(N__35997),
            .in2(N__32874),
            .in3(N__34510),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIJR3Q5Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_esr_RNIB9IP_0_LC_2_18_0 .C_ON=1'b1;
    defparam \pid_alt.error_i_acumm_esr_RNIB9IP_0_LC_2_18_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_esr_RNIB9IP_0_LC_2_18_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \pid_alt.error_i_acumm_esr_RNIB9IP_0_LC_2_18_0  (
            .in0(_gnd_net_),
            .in1(N__37311),
            .in2(N__36839),
            .in3(_gnd_net_),
            .lcout(\pid_alt.un1_pid_prereg_0 ),
            .ltout(),
            .carryin(bfn_2_18_0_),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_esr_RNIQMD91_1_LC_2_18_1 .C_ON=1'b1;
    defparam \pid_alt.error_i_acumm_esr_RNIQMD91_1_LC_2_18_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_esr_RNIQMD91_1_LC_2_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_i_acumm_esr_RNIQMD91_1_LC_2_18_1  (
            .in0(_gnd_net_),
            .in1(N__37368),
            .in2(N__32871),
            .in3(N__32856),
            .lcout(\pid_alt.error_i_acumm_esr_RNIQMD91Z0Z_1 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_0 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_esr_RNITQE91_2_LC_2_18_2 .C_ON=1'b1;
    defparam \pid_alt.error_i_acumm_esr_RNITQE91_2_LC_2_18_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_esr_RNITQE91_2_LC_2_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_i_acumm_esr_RNITQE91_2_LC_2_18_2  (
            .in0(_gnd_net_),
            .in1(N__37341),
            .in2(N__32853),
            .in3(N__32838),
            .lcout(\pid_alt.error_i_acumm_esr_RNITQE91Z0Z_2 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_1 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_esr_RNI0VF91_3_LC_2_18_3 .C_ON=1'b1;
    defparam \pid_alt.error_i_acumm_esr_RNI0VF91_3_LC_2_18_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_esr_RNI0VF91_3_LC_2_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_i_acumm_esr_RNI0VF91_3_LC_2_18_3  (
            .in0(_gnd_net_),
            .in1(N__37218),
            .in2(N__32835),
            .in3(N__32820),
            .lcout(\pid_alt.error_i_acumm_esr_RNI0VF91Z0Z_3 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_2 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_esr_RNI33H91_4_LC_2_18_4 .C_ON=1'b1;
    defparam \pid_alt.error_i_acumm_esr_RNI33H91_4_LC_2_18_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_esr_RNI33H91_4_LC_2_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_i_acumm_esr_RNI33H91_4_LC_2_18_4  (
            .in0(_gnd_net_),
            .in1(N__37293),
            .in2(N__32817),
            .in3(N__32802),
            .lcout(\pid_alt.error_i_acumm_esr_RNI33H91Z0Z_4 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_3 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_reg_esr_RNIT8KA1_5_LC_2_18_5 .C_ON=1'b1;
    defparam \pid_alt.error_i_reg_esr_RNIT8KA1_5_LC_2_18_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_reg_esr_RNIT8KA1_5_LC_2_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_i_reg_esr_RNIT8KA1_5_LC_2_18_5  (
            .in0(_gnd_net_),
            .in1(N__48405),
            .in2(N__32799),
            .in3(N__32781),
            .lcout(\pid_alt.error_i_reg_esr_RNIT8KA1Z0Z_5 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_4 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_5_c_RNI0DLQ_LC_2_18_6 .C_ON=1'b1;
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_5_c_RNI0DLQ_LC_2_18_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_5_c_RNI0DLQ_LC_2_18_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_5_c_RNI0DLQ_LC_2_18_6  (
            .in0(_gnd_net_),
            .in1(N__39576),
            .in2(N__33120),
            .in3(N__33102),
            .lcout(\pid_alt.un1_error_i_acumm_prereg_cry_5_c_RNI0DLQ ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_5 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_6_c_RNI3HMQ_LC_2_18_7 .C_ON=1'b1;
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_6_c_RNI3HMQ_LC_2_18_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_6_c_RNI3HMQ_LC_2_18_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_6_c_RNI3HMQ_LC_2_18_7  (
            .in0(_gnd_net_),
            .in1(N__39522),
            .in2(N__33099),
            .in3(N__33078),
            .lcout(\pid_alt.un1_error_i_acumm_prereg_cry_6_c_RNI3HMQ ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_6 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_7_c_RNI6LNQ_LC_2_19_0 .C_ON=1'b1;
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_7_c_RNI6LNQ_LC_2_19_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_7_c_RNI6LNQ_LC_2_19_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_7_c_RNI6LNQ_LC_2_19_0  (
            .in0(_gnd_net_),
            .in1(N__39480),
            .in2(N__33075),
            .in3(N__33057),
            .lcout(\pid_alt.un1_error_i_acumm_prereg_cry_7_c_RNI6LNQ ),
            .ltout(),
            .carryin(bfn_2_19_0_),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_8_c_RNI9POQ_LC_2_19_1 .C_ON=1'b1;
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_8_c_RNI9POQ_LC_2_19_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_8_c_RNI9POQ_LC_2_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_8_c_RNI9POQ_LC_2_19_1  (
            .in0(_gnd_net_),
            .in1(N__39387),
            .in2(N__33054),
            .in3(N__33024),
            .lcout(\pid_alt.un1_error_i_acumm_prereg_cry_8_c_RNI9POQ ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_8 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_9_c_RNIQN3F_LC_2_19_2 .C_ON=1'b1;
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_9_c_RNIQN3F_LC_2_19_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_9_c_RNIQN3F_LC_2_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_9_c_RNIQN3F_LC_2_19_2  (
            .in0(_gnd_net_),
            .in1(N__39078),
            .in2(N__33021),
            .in3(N__33006),
            .lcout(\pid_alt.un1_error_i_acumm_prereg_cry_9_c_RNIQN3F ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_9 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_reg_esr_RNI4NMP_11_LC_2_19_3 .C_ON=1'b1;
    defparam \pid_alt.error_i_reg_esr_RNI4NMP_11_LC_2_19_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_reg_esr_RNI4NMP_11_LC_2_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_i_reg_esr_RNI4NMP_11_LC_2_19_3  (
            .in0(_gnd_net_),
            .in1(N__39624),
            .in2(N__33003),
            .in3(N__32985),
            .lcout(\pid_alt.error_i_reg_esr_RNI4NMPZ0Z_11 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_10 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_reg_esr_RNI7RNP_12_LC_2_19_4 .C_ON=1'b1;
    defparam \pid_alt.error_i_reg_esr_RNI7RNP_12_LC_2_19_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_reg_esr_RNI7RNP_12_LC_2_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_i_reg_esr_RNI7RNP_12_LC_2_19_4  (
            .in0(_gnd_net_),
            .in1(N__39330),
            .in2(N__32982),
            .in3(N__32964),
            .lcout(\pid_alt.error_i_reg_esr_RNI7RNPZ0Z_12 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_11 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_esr_RNIJ6LM_13_LC_2_19_5 .C_ON=1'b1;
    defparam \pid_alt.error_i_acumm_esr_RNIJ6LM_13_LC_2_19_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_esr_RNIJ6LM_13_LC_2_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_i_acumm_esr_RNIJ6LM_13_LC_2_19_5  (
            .in0(_gnd_net_),
            .in1(N__49401),
            .in2(N__32961),
            .in3(N__32946),
            .lcout(\pid_alt.error_i_acumm_esr_RNIJ6LMZ0Z_13 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_12 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_reg_esr_RNI15KJ_14_LC_2_19_6 .C_ON=1'b1;
    defparam \pid_alt.error_i_reg_esr_RNI15KJ_14_LC_2_19_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_reg_esr_RNI15KJ_14_LC_2_19_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_i_reg_esr_RNI15KJ_14_LC_2_19_6  (
            .in0(_gnd_net_),
            .in1(N__33249),
            .in2(_gnd_net_),
            .in3(N__33234),
            .lcout(\pid_alt.error_i_reg_esr_RNI15KJZ0Z_14 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_13 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_reg_esr_RNI38LJ_15_LC_2_19_7 .C_ON=1'b1;
    defparam \pid_alt.error_i_reg_esr_RNI38LJ_15_LC_2_19_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_reg_esr_RNI38LJ_15_LC_2_19_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_i_reg_esr_RNI38LJ_15_LC_2_19_7  (
            .in0(_gnd_net_),
            .in1(N__33231),
            .in2(_gnd_net_),
            .in3(N__33216),
            .lcout(\pid_alt.error_i_reg_esr_RNI38LJZ0Z_15 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_14 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_reg_esr_RNI5BMJ_16_LC_2_20_0 .C_ON=1'b1;
    defparam \pid_alt.error_i_reg_esr_RNI5BMJ_16_LC_2_20_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_reg_esr_RNI5BMJ_16_LC_2_20_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_i_reg_esr_RNI5BMJ_16_LC_2_20_0  (
            .in0(_gnd_net_),
            .in1(N__33213),
            .in2(_gnd_net_),
            .in3(N__33198),
            .lcout(\pid_alt.error_i_reg_esr_RNI5BMJZ0Z_16 ),
            .ltout(),
            .carryin(bfn_2_20_0_),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_reg_esr_RNI7ENJ_17_LC_2_20_1 .C_ON=1'b1;
    defparam \pid_alt.error_i_reg_esr_RNI7ENJ_17_LC_2_20_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_reg_esr_RNI7ENJ_17_LC_2_20_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_i_reg_esr_RNI7ENJ_17_LC_2_20_1  (
            .in0(_gnd_net_),
            .in1(N__33195),
            .in2(_gnd_net_),
            .in3(N__33180),
            .lcout(\pid_alt.error_i_reg_esr_RNI7ENJZ0Z_17 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_16 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_reg_esr_RNI9HOJ_18_LC_2_20_2 .C_ON=1'b1;
    defparam \pid_alt.error_i_reg_esr_RNI9HOJ_18_LC_2_20_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_reg_esr_RNI9HOJ_18_LC_2_20_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_i_reg_esr_RNI9HOJ_18_LC_2_20_2  (
            .in0(_gnd_net_),
            .in1(N__33177),
            .in2(_gnd_net_),
            .in3(N__33162),
            .lcout(\pid_alt.error_i_reg_esr_RNI9HOJZ0Z_18 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_17 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_reg_esr_RNIBKPJ_19_LC_2_20_3 .C_ON=1'b1;
    defparam \pid_alt.error_i_reg_esr_RNIBKPJ_19_LC_2_20_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_reg_esr_RNIBKPJ_19_LC_2_20_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_i_reg_esr_RNIBKPJ_19_LC_2_20_3  (
            .in0(_gnd_net_),
            .in1(N__33159),
            .in2(_gnd_net_),
            .in3(N__33144),
            .lcout(\pid_alt.error_i_reg_esr_RNIBKPJZ0Z_19 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_18 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_19_c_RNI4FRJ_LC_2_20_4 .C_ON=1'b1;
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_19_c_RNI4FRJ_LC_2_20_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_19_c_RNI4FRJ_LC_2_20_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_19_c_RNI4FRJ_LC_2_20_4  (
            .in0(_gnd_net_),
            .in1(N__33137),
            .in2(_gnd_net_),
            .in3(N__33141),
            .lcout(\pid_alt.un1_error_i_acumm_prereg_cry_19_c_RNI4FRJ ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_19 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_20_c_RNISVKK_LC_2_20_5 .C_ON=1'b0;
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_20_c_RNISVKK_LC_2_20_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_20_c_RNISVKK_LC_2_20_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_20_c_RNISVKK_LC_2_20_5  (
            .in0(N__33138),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33123),
            .lcout(\pid_alt.un1_error_i_acumm_prereg_cry_20_c_RNISVKK ),
            .ltout(\pid_alt.un1_error_i_acumm_prereg_cry_20_c_RNISVKK_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNO_0_24_LC_2_20_6 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNO_0_24_LC_2_20_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNO_0_24_LC_2_20_6 .LUT_INIT=16'b1111111001111111;
    LogicCell40 \pid_alt.pid_prereg_esr_RNO_0_24_LC_2_20_6  (
            .in0(N__35150),
            .in1(N__35103),
            .in2(N__33378),
            .in3(N__35180),
            .lcout(\pid_alt.un1_pid_prereg_0_axb_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI20IM_0_17_LC_2_20_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI20IM_0_17_LC_2_20_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI20IM_0_17_LC_2_20_7 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI20IM_0_17_LC_2_20_7  (
            .in0(N__33374),
            .in1(N__33284),
            .in2(_gnd_net_),
            .in3(N__33327),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI20IM_0Z0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_11_LC_2_21_0 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_11_LC_2_21_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_11_LC_2_21_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_11_LC_2_21_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33363),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87268),
            .ce(N__51479),
            .sr(N__79670));
    defparam \pid_alt.error_i_acumm_prereg_esr_17_LC_2_21_1 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_17_LC_2_21_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_17_LC_2_21_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_17_LC_2_21_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35370),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87268),
            .ce(N__51479),
            .sr(N__79670));
    defparam \pid_alt.error_i_acumm_prereg_esr_21_LC_2_21_2 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_21_LC_2_21_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_21_LC_2_21_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_21_LC_2_21_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35058),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87268),
            .ce(N__51479),
            .sr(N__79670));
    defparam \pid_alt.error_i_acumm_prereg_esr_18_LC_2_21_3 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_18_LC_2_21_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_18_LC_2_21_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_18_LC_2_21_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33342),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87268),
            .ce(N__51479),
            .sr(N__79670));
    defparam \pid_alt.error_i_acumm_prereg_esr_20_LC_2_21_5 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_20_LC_2_21_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_20_LC_2_21_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_20_LC_2_21_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34755),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87268),
            .ce(N__51479),
            .sr(N__79670));
    defparam \pid_alt.error_d_reg_prev_esr_17_LC_2_21_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_17_LC_2_21_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_17_LC_2_21_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_17_LC_2_21_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33323),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87268),
            .ce(N__51479),
            .sr(N__79670));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIC8F4_16_LC_2_22_0 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIC8F4_16_LC_2_22_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIC8F4_16_LC_2_22_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNIC8F4_16_LC_2_22_0  (
            .in0(N__33273),
            .in1(N__33564),
            .in2(N__33267),
            .in3(N__33588),
            .lcout(),
            .ltout(\pid_alt.m7_e_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIRRP7_14_LC_2_22_1 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIRRP7_14_LC_2_22_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIRRP7_14_LC_2_22_1 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNIRRP7_14_LC_2_22_1  (
            .in0(N__33258),
            .in1(N__35430),
            .in2(N__33252),
            .in3(N__33558),
            .lcout(\pid_alt.N_545 ),
            .ltout(\pid_alt.N_545_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI175B_12_LC_2_22_2 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI175B_12_LC_2_22_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI175B_12_LC_2_22_2 .LUT_INIT=16'b1101110011111100;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNI175B_12_LC_2_22_2  (
            .in0(N__49439),
            .in1(N__49464),
            .in2(N__33591),
            .in3(N__39369),
            .lcout(\pid_alt.N_158 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_16_LC_2_22_3 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_16_LC_2_22_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_16_LC_2_22_3 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_16_LC_2_22_3  (
            .in0(_gnd_net_),
            .in1(N__35265),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87273),
            .ce(N__51476),
            .sr(N__79676));
    defparam \pid_alt.error_i_acumm_prereg_esr_19_LC_2_22_5 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_19_LC_2_22_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_19_LC_2_22_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_19_LC_2_22_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33582),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87273),
            .ce(N__51476),
            .sr(N__79676));
    defparam \pid_alt.error_i_acumm_prereg_esr_14_LC_2_22_7 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_14_LC_2_22_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_14_LC_2_22_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_14_LC_2_22_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36370),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87273),
            .ce(N__51476),
            .sr(N__79676));
    defparam \pid_alt.error_p_reg_esr_8_LC_2_23_2 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_8_LC_2_23_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_8_LC_2_23_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_8_LC_2_23_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33552),
            .lcout(\pid_alt.error_p_regZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87277),
            .ce(N__33467),
            .sr(N__86026));
    defparam \pid_alt.error_p_reg_esr_1_LC_2_23_4 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_1_LC_2_23_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_1_LC_2_23_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_1_LC_2_23_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33519),
            .lcout(\pid_alt.error_p_regZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87277),
            .ce(N__33467),
            .sr(N__86026));
    defparam \pid_alt.error_p_reg_esr_3_LC_2_23_7 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_3_LC_2_23_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_3_LC_2_23_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_3_LC_2_23_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33492),
            .lcout(\pid_alt.error_p_regZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87277),
            .ce(N__33467),
            .sr(N__86026));
    defparam \Commands_frame_decoder.source_alt_kd_0_LC_3_6_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kd_0_LC_3_6_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kd_0_LC_3_6_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_kd_0_LC_3_6_1  (
            .in0(_gnd_net_),
            .in1(N__83797),
            .in2(_gnd_net_),
            .in3(N__86185),
            .lcout(alt_kd_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87072),
            .ce(N__33408),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.WDT_RNIRGQ51_11_LC_3_9_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.WDT_RNIRGQ51_11_LC_3_9_0 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.WDT_RNIRGQ51_11_LC_3_9_0 .LUT_INIT=16'b0101010101110111;
    LogicCell40 \Commands_frame_decoder.WDT_RNIRGQ51_11_LC_3_9_0  (
            .in0(N__33870),
            .in1(N__33846),
            .in2(_gnd_net_),
            .in3(N__33825),
            .lcout(\Commands_frame_decoder.state_0_sqmuxacf0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.preinit_RNIR9JL1_LC_3_9_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.preinit_RNIR9JL1_LC_3_9_1 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.preinit_RNIR9JL1_LC_3_9_1 .LUT_INIT=16'b0000010100000111;
    LogicCell40 \Commands_frame_decoder.preinit_RNIR9JL1_LC_3_9_1  (
            .in0(N__34127),
            .in1(N__34157),
            .in2(N__33645),
            .in3(N__33871),
            .lcout(\Commands_frame_decoder.state_0_sqmuxacf1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.WDT_RNIET8A1_0_4_LC_3_9_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.WDT_RNIET8A1_0_4_LC_3_9_2 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.WDT_RNIET8A1_0_4_LC_3_9_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \Commands_frame_decoder.WDT_RNIET8A1_0_4_LC_3_9_2  (
            .in0(N__33805),
            .in1(N__33787),
            .in2(N__33770),
            .in3(N__33745),
            .lcout(),
            .ltout(\Commands_frame_decoder.WDT8lto9_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.WDT_RNII01C2_8_LC_3_9_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.WDT_RNII01C2_8_LC_3_9_3 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.WDT_RNII01C2_8_LC_3_9_3 .LUT_INIT=16'b1010101010001010;
    LogicCell40 \Commands_frame_decoder.WDT_RNII01C2_8_LC_3_9_3  (
            .in0(N__33890),
            .in1(N__33608),
            .in2(N__33687),
            .in3(N__33626),
            .lcout(\Commands_frame_decoder.WDT8lt12_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.preinit_RNIC9QE2_LC_3_9_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.preinit_RNIC9QE2_LC_3_9_4 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.preinit_RNIC9QE2_LC_3_9_4 .LUT_INIT=16'b0000000001110011;
    LogicCell40 \Commands_frame_decoder.preinit_RNIC9QE2_LC_3_9_4  (
            .in0(N__34158),
            .in1(N__34128),
            .in2(N__33684),
            .in3(N__33642),
            .lcout(),
            .ltout(\Commands_frame_decoder.state_0_sqmuxacf0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.WDT_RNIPJEG6_8_LC_3_9_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.WDT_RNIPJEG6_8_LC_3_9_5 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.WDT_RNIPJEG6_8_LC_3_9_5 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \Commands_frame_decoder.WDT_RNIPJEG6_8_LC_3_9_5  (
            .in0(_gnd_net_),
            .in1(N__33675),
            .in2(N__33669),
            .in3(N__33666),
            .lcout(\Commands_frame_decoder.state_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.preinit_LC_3_9_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.preinit_LC_3_9_6 .SEQ_MODE=4'b1001;
    defparam \Commands_frame_decoder.preinit_LC_3_9_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Commands_frame_decoder.preinit_LC_3_9_6  (
            .in0(_gnd_net_),
            .in1(N__38465),
            .in2(_gnd_net_),
            .in3(N__33644),
            .lcout(\Commands_frame_decoder.preinitZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87115),
            .ce(),
            .sr(N__79580));
    defparam \Commands_frame_decoder.source_data_valid_LC_3_9_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_data_valid_LC_3_9_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_data_valid_LC_3_9_7 .LUT_INIT=16'b1111101011001010;
    LogicCell40 \Commands_frame_decoder.source_data_valid_LC_3_9_7  (
            .in0(N__33643),
            .in1(N__41344),
            .in2(N__38469),
            .in3(N__33696),
            .lcout(debug_CH3_20A_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87115),
            .ce(),
            .sr(N__79580));
    defparam \Commands_frame_decoder.WDT_RNITK4L_8_LC_3_10_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.WDT_RNITK4L_8_LC_3_10_0 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.WDT_RNITK4L_8_LC_3_10_0 .LUT_INIT=16'b0001000100010001;
    LogicCell40 \Commands_frame_decoder.WDT_RNITK4L_8_LC_3_10_0  (
            .in0(N__33625),
            .in1(N__33607),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\Commands_frame_decoder.WDT_RNITK4LZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.WDT_RNI2VDI1_10_LC_3_10_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.WDT_RNI2VDI1_10_LC_3_10_1 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.WDT_RNI2VDI1_10_LC_3_10_1 .LUT_INIT=16'b0000000111111111;
    LogicCell40 \Commands_frame_decoder.WDT_RNI2VDI1_10_LC_3_10_1  (
            .in0(N__33827),
            .in1(N__33889),
            .in2(N__33852),
            .in3(N__33872),
            .lcout(\Commands_frame_decoder.WDT_RNI2VDI1Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.WDT_RNIHV6P_11_LC_3_10_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.WDT_RNIHV6P_11_LC_3_10_2 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.WDT_RNIHV6P_11_LC_3_10_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \Commands_frame_decoder.WDT_RNIHV6P_11_LC_3_10_2  (
            .in0(_gnd_net_),
            .in1(N__33847),
            .in2(_gnd_net_),
            .in3(N__33826),
            .lcout(\Commands_frame_decoder.WDT_RNIHV6PZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.WDT_RNIET8A1_4_LC_3_10_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.WDT_RNIET8A1_4_LC_3_10_3 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.WDT_RNIET8A1_4_LC_3_10_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \Commands_frame_decoder.WDT_RNIET8A1_4_LC_3_10_3  (
            .in0(N__33806),
            .in1(N__33788),
            .in2(N__33771),
            .in3(N__33746),
            .lcout(),
            .ltout(\Commands_frame_decoder.WDT_RNIET8A1Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.WDT_RNIUG2B4_4_LC_3_10_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.WDT_RNIUG2B4_4_LC_3_10_4 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.WDT_RNIUG2B4_4_LC_3_10_4 .LUT_INIT=16'b0001010101010101;
    LogicCell40 \Commands_frame_decoder.WDT_RNIUG2B4_4_LC_3_10_4  (
            .in0(N__33729),
            .in1(N__33723),
            .in2(N__33717),
            .in3(N__33714),
            .lcout(\Commands_frame_decoder.WDT8lt14_0 ),
            .ltout(\Commands_frame_decoder.WDT8lt14_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.WDT_RNIPRJG5_15_LC_3_10_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.WDT_RNIPRJG5_15_LC_3_10_5 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.WDT_RNIPRJG5_15_LC_3_10_5 .LUT_INIT=16'b0100010001000000;
    LogicCell40 \Commands_frame_decoder.WDT_RNIPRJG5_15_LC_3_10_5  (
            .in0(N__38401),
            .in1(N__34129),
            .in2(N__33708),
            .in3(N__34159),
            .lcout(\Commands_frame_decoder.N_365_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNIQRI31_10_LC_3_10_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIQRI31_10_LC_3_10_6 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIQRI31_10_LC_3_10_6 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \Commands_frame_decoder.state_RNIQRI31_10_LC_3_10_6  (
            .in0(N__39239),
            .in1(N__38402),
            .in2(_gnd_net_),
            .in3(N__79967),
            .lcout(\Commands_frame_decoder.state_RNIQRI31Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNITVPE1_1_LC_3_11_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNITVPE1_1_LC_3_11_0 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNITVPE1_1_LC_3_11_0 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \Commands_frame_decoder.state_RNITVPE1_1_LC_3_11_0  (
            .in0(N__83723),
            .in1(N__33942),
            .in2(N__85378),
            .in3(N__35685),
            .lcout(\Commands_frame_decoder.N_406 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.count_0_LC_3_11_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.count_0_LC_3_11_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.count_0_LC_3_11_2 .LUT_INIT=16'b0000000001111000;
    LogicCell40 \Commands_frame_decoder.count_0_LC_3_11_2  (
            .in0(N__33911),
            .in1(N__38462),
            .in2(N__34014),
            .in3(N__79932),
            .lcout(\Commands_frame_decoder.countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87148),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_data_valid_RNO_0_LC_3_11_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_data_valid_RNO_0_LC_3_11_3 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.source_data_valid_RNO_0_LC_3_11_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Commands_frame_decoder.source_data_valid_RNO_0_LC_3_11_3  (
            .in0(_gnd_net_),
            .in1(N__34009),
            .in2(_gnd_net_),
            .in3(N__33910),
            .lcout(\Commands_frame_decoder.count_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.un1_state57_i_LC_3_11_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.un1_state57_i_LC_3_11_4 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.un1_state57_i_LC_3_11_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \Commands_frame_decoder.un1_state57_i_LC_3_11_4  (
            .in0(_gnd_net_),
            .in1(N__38460),
            .in2(_gnd_net_),
            .in3(N__79931),
            .lcout(\Commands_frame_decoder.un1_state57_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_4_LC_3_11_5 .C_ON=1'b0;
    defparam \uart_pc.data_4_LC_3_11_5 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_4_LC_3_11_5 .LUT_INIT=16'b0101000101000000;
    LogicCell40 \uart_pc.data_4_LC_3_11_5  (
            .in0(N__35757),
            .in1(N__38160),
            .in2(N__38037),
            .in3(N__84983),
            .lcout(uart_pc_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87148),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNIG48S_7_LC_3_11_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIG48S_7_LC_3_11_6 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIG48S_7_LC_3_11_6 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \Commands_frame_decoder.state_RNIG48S_7_LC_3_11_6  (
            .in0(N__34058),
            .in1(N__38461),
            .in2(_gnd_net_),
            .in3(N__79930),
            .lcout(\Commands_frame_decoder.state_RNIG48SZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.count_RNIA5DM6_0_LC_3_11_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.count_RNIA5DM6_0_LC_3_11_7 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.count_RNIA5DM6_0_LC_3_11_7 .LUT_INIT=16'b0000000001110000;
    LogicCell40 \Commands_frame_decoder.count_RNIA5DM6_0_LC_3_11_7  (
            .in0(N__38459),
            .in1(N__34010),
            .in2(N__33915),
            .in3(N__33980),
            .lcout(\Commands_frame_decoder.N_372 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNI6QPK_1_LC_3_12_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNI6QPK_1_LC_3_12_0 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNI6QPK_1_LC_3_12_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \Commands_frame_decoder.state_RNI6QPK_1_LC_3_12_0  (
            .in0(_gnd_net_),
            .in1(N__33909),
            .in2(_gnd_net_),
            .in3(N__33939),
            .lcout(\Commands_frame_decoder.N_370_2 ),
            .ltout(\Commands_frame_decoder.N_370_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNO_0_0_LC_3_12_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNO_0_0_LC_3_12_1 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNO_0_0_LC_3_12_1 .LUT_INIT=16'b0011001100100011;
    LogicCell40 \Commands_frame_decoder.state_RNO_0_0_LC_3_12_1  (
            .in0(N__33966),
            .in1(N__33993),
            .in2(N__33987),
            .in3(N__33984),
            .lcout(),
            .ltout(\Commands_frame_decoder.state_ns_i_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_0_LC_3_12_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_0_LC_3_12_2 .SEQ_MODE=4'b1001;
    defparam \Commands_frame_decoder.state_0_LC_3_12_2 .LUT_INIT=16'b0001000001010000;
    LogicCell40 \Commands_frame_decoder.state_0_LC_3_12_2  (
            .in0(N__33923),
            .in1(N__39298),
            .in2(N__33969),
            .in3(N__33940),
            .lcout(\Commands_frame_decoder.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87164),
            .ce(),
            .sr(N__79598));
    defparam \Commands_frame_decoder.state_1_LC_3_12_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_1_LC_3_12_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_1_LC_3_12_3 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \Commands_frame_decoder.state_1_LC_3_12_3  (
            .in0(N__33941),
            .in1(N__34196),
            .in2(N__33954),
            .in3(N__39289),
            .lcout(\Commands_frame_decoder.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87164),
            .ce(),
            .sr(N__79598));
    defparam \Commands_frame_decoder.state_14_LC_3_12_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_14_LC_3_12_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_14_LC_3_12_4 .LUT_INIT=16'b1111101010101010;
    LogicCell40 \Commands_frame_decoder.state_14_LC_3_12_4  (
            .in0(N__33924),
            .in1(_gnd_net_),
            .in2(N__34215),
            .in3(N__38400),
            .lcout(\Commands_frame_decoder.stateZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87164),
            .ce(),
            .sr(N__79598));
    defparam \Commands_frame_decoder.state_13_LC_3_12_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_13_LC_3_12_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_13_LC_3_12_5 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \Commands_frame_decoder.state_13_LC_3_12_5  (
            .in0(N__34214),
            .in1(N__39896),
            .in2(_gnd_net_),
            .in3(N__39288),
            .lcout(\Commands_frame_decoder.stateZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87164),
            .ce(),
            .sr(N__79598));
    defparam \Commands_frame_decoder.state_RNITUI31_13_LC_3_12_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNITUI31_13_LC_3_12_6 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNITUI31_13_LC_3_12_6 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \Commands_frame_decoder.state_RNITUI31_13_LC_3_12_6  (
            .in0(N__34210),
            .in1(N__38399),
            .in2(_gnd_net_),
            .in3(N__79924),
            .lcout(\Commands_frame_decoder.state_RNITUI31Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_2_LC_3_12_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_2_LC_3_12_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_2_LC_3_12_7 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \Commands_frame_decoder.state_2_LC_3_12_7  (
            .in0(N__38534),
            .in1(N__34197),
            .in2(N__34188),
            .in3(N__39290),
            .lcout(\Commands_frame_decoder.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87164),
            .ce(),
            .sr(N__79598));
    defparam \Commands_frame_decoder.state_12_LC_3_13_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_12_LC_3_13_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_12_LC_3_13_0 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \Commands_frame_decoder.state_12_LC_3_13_0  (
            .in0(N__38231),
            .in1(N__38448),
            .in2(N__34101),
            .in3(N__39283),
            .lcout(\Commands_frame_decoder.stateZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87178),
            .ce(),
            .sr(N__79603));
    defparam \Commands_frame_decoder.WDT_RNIPRJG5_0_15_LC_3_13_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.WDT_RNIPRJG5_0_15_LC_3_13_1 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.WDT_RNIPRJG5_0_15_LC_3_13_1 .LUT_INIT=16'b0000000100001111;
    LogicCell40 \Commands_frame_decoder.WDT_RNIPRJG5_0_15_LC_3_13_1  (
            .in0(N__34173),
            .in1(N__34164),
            .in2(N__38463),
            .in3(N__34134),
            .lcout(\Commands_frame_decoder.N_403 ),
            .ltout(\Commands_frame_decoder.N_403_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_11_LC_3_13_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_11_LC_3_13_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_11_LC_3_13_2 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \Commands_frame_decoder.state_11_LC_3_13_2  (
            .in0(N__34100),
            .in1(N__39240),
            .in2(N__34104),
            .in3(N__38447),
            .lcout(\Commands_frame_decoder.stateZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87178),
            .ce(),
            .sr(N__79603));
    defparam \Commands_frame_decoder.state_8_LC_3_13_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_8_LC_3_13_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_8_LC_3_13_4 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \Commands_frame_decoder.state_8_LC_3_13_4  (
            .in0(N__34056),
            .in1(N__38450),
            .in2(N__34083),
            .in3(N__39286),
            .lcout(\Commands_frame_decoder.stateZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87178),
            .ce(),
            .sr(N__79603));
    defparam \Commands_frame_decoder.state_9_LC_3_13_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_9_LC_3_13_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_9_LC_3_13_5 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \Commands_frame_decoder.state_9_LC_3_13_5  (
            .in0(N__39287),
            .in1(N__34079),
            .in2(N__38464),
            .in3(N__34071),
            .lcout(\Commands_frame_decoder.stateZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87178),
            .ce(),
            .sr(N__79603));
    defparam \Commands_frame_decoder.state_7_LC_3_13_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_7_LC_3_13_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_7_LC_3_13_6 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \Commands_frame_decoder.state_7_LC_3_13_6  (
            .in0(N__34057),
            .in1(N__38449),
            .in2(N__38213),
            .in3(N__39285),
            .lcout(\Commands_frame_decoder.stateZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87178),
            .ce(),
            .sr(N__79603));
    defparam \Commands_frame_decoder.state_6_LC_3_13_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_6_LC_3_13_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_6_LC_3_13_7 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \Commands_frame_decoder.state_6_LC_3_13_7  (
            .in0(N__39284),
            .in1(N__38209),
            .in2(_gnd_net_),
            .in3(N__35679),
            .lcout(\Commands_frame_decoder.stateZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87178),
            .ce(),
            .sr(N__79603));
    defparam \pid_alt.pid_prereg_esr_RNIBRUM_15_LC_3_14_0 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNIBRUM_15_LC_3_14_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNIBRUM_15_LC_3_14_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_alt.pid_prereg_esr_RNIBRUM_15_LC_3_14_0  (
            .in0(N__34437),
            .in1(N__34539),
            .in2(N__34572),
            .in3(N__34641),
            .lcout(),
            .ltout(\pid_alt.source_pid_1_sqmuxa_0_a2_2_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNIT4CP1_14_LC_3_14_1 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNIT4CP1_14_LC_3_14_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNIT4CP1_14_LC_3_14_1 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \pid_alt.pid_prereg_esr_RNIT4CP1_14_LC_3_14_1  (
            .in0(N__34425),
            .in1(N__34449),
            .in2(N__34290),
            .in3(N__34281),
            .lcout(\pid_alt.N_539 ),
            .ltout(\pid_alt.N_539_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.source_pid_1_esr_RNO_0_4_LC_3_14_2 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_esr_RNO_0_4_LC_3_14_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.source_pid_1_esr_RNO_0_4_LC_3_14_2 .LUT_INIT=16'b0000000011101010;
    LogicCell40 \pid_alt.source_pid_1_esr_RNO_0_4_LC_3_14_2  (
            .in0(N__37623),
            .in1(N__35640),
            .in2(N__34287),
            .in3(N__35568),
            .lcout(),
            .ltout(\pid_alt.source_pid_9_0_0_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.source_pid_1_esr_4_LC_3_14_3 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_esr_4_LC_3_14_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_esr_4_LC_3_14_3 .LUT_INIT=16'b0000101100001111;
    LogicCell40 \pid_alt.source_pid_1_esr_4_LC_3_14_3  (
            .in0(N__35569),
            .in1(N__35594),
            .in2(N__34284),
            .in3(N__37694),
            .lcout(throttle_order_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87192),
            .ce(N__35529),
            .sr(N__37818));
    defparam \pid_alt.pid_prereg_esr_RNICSUM_17_LC_3_14_4 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNICSUM_17_LC_3_14_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNICSUM_17_LC_3_14_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_alt.pid_prereg_esr_RNICSUM_17_LC_3_14_4  (
            .in0(N__34584),
            .in1(N__34596),
            .in2(N__34557),
            .in3(N__34413),
            .lcout(\pid_alt.source_pid_1_sqmuxa_0_a2_2_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.source_pid_1_esr_5_LC_3_14_5 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_esr_5_LC_3_14_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_esr_5_LC_3_14_5 .LUT_INIT=16'b1110000010100000;
    LogicCell40 \pid_alt.source_pid_1_esr_5_LC_3_14_5  (
            .in0(N__37624),
            .in1(N__37693),
            .in2(N__35661),
            .in3(N__35595),
            .lcout(throttle_order_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87192),
            .ce(N__35529),
            .sr(N__37818));
    defparam \pid_alt.un1_pid_prereg_un1_pid_prereg_0_cry_0_c_THRU_CRY_0_LC_3_15_0 .C_ON=1'b1;
    defparam \pid_alt.un1_pid_prereg_un1_pid_prereg_0_cry_0_c_THRU_CRY_0_LC_3_15_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un1_pid_prereg_un1_pid_prereg_0_cry_0_c_THRU_CRY_0_LC_3_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_alt.un1_pid_prereg_un1_pid_prereg_0_cry_0_c_THRU_CRY_0_LC_3_15_0  (
            .in0(_gnd_net_),
            .in1(N__34265),
            .in2(N__34275),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_3_15_0_),
            .carryout(\pid_alt.un1_pid_prereg_un1_pid_prereg_0_cry_0_c_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_0_LC_3_15_1 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_0_LC_3_15_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_0_LC_3_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_0_LC_3_15_1  (
            .in0(_gnd_net_),
            .in1(N__34251),
            .in2(N__34245),
            .in3(N__34218),
            .lcout(\pid_alt.pid_preregZ0Z_0 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_un1_pid_prereg_0_cry_0_c_THRU_CO ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_0 ),
            .clk(N__87209),
            .ce(N__51492),
            .sr(N__79614));
    defparam \pid_alt.pid_prereg_esr_1_LC_3_15_2 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_1_LC_3_15_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_1_LC_3_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_1_LC_3_15_2  (
            .in0(_gnd_net_),
            .in1(N__36872),
            .in2(N__34401),
            .in3(N__34392),
            .lcout(\pid_alt.pid_preregZ0Z_1 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_0 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_1 ),
            .clk(N__87209),
            .ce(N__51492),
            .sr(N__79614));
    defparam \pid_alt.pid_prereg_esr_2_LC_3_15_3 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_2_LC_3_15_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_2_LC_3_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_2_LC_3_15_3  (
            .in0(_gnd_net_),
            .in1(N__34389),
            .in2(N__35214),
            .in3(N__34383),
            .lcout(\pid_alt.pid_preregZ0Z_2 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_1 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_2 ),
            .clk(N__87209),
            .ce(N__51492),
            .sr(N__79614));
    defparam \pid_alt.pid_prereg_esr_3_LC_3_15_4 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_3_LC_3_15_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_3_LC_3_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_3_LC_3_15_4  (
            .in0(_gnd_net_),
            .in1(N__34380),
            .in2(N__35424),
            .in3(N__34374),
            .lcout(\pid_alt.pid_preregZ0Z_3 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_2 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_3 ),
            .clk(N__87209),
            .ce(N__51492),
            .sr(N__79614));
    defparam \pid_alt.pid_prereg_esr_4_LC_3_15_5 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_4_LC_3_15_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_4_LC_3_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_4_LC_3_15_5  (
            .in0(_gnd_net_),
            .in1(N__34367),
            .in2(N__34356),
            .in3(N__34347),
            .lcout(\pid_alt.pid_preregZ0Z_4 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_3 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_4 ),
            .clk(N__87209),
            .ce(N__51492),
            .sr(N__79614));
    defparam \pid_alt.pid_prereg_esr_5_LC_3_15_6 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_5_LC_3_15_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_5_LC_3_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_5_LC_3_15_6  (
            .in0(_gnd_net_),
            .in1(N__36209),
            .in2(N__36177),
            .in3(N__34344),
            .lcout(\pid_alt.pid_preregZ0Z_5 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_4 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_5 ),
            .clk(N__87209),
            .ce(N__51492),
            .sr(N__79614));
    defparam \pid_alt.pid_prereg_esr_6_LC_3_15_7 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_6_LC_3_15_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_6_LC_3_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_6_LC_3_15_7  (
            .in0(_gnd_net_),
            .in1(N__35859),
            .in2(N__35853),
            .in3(N__34341),
            .lcout(\pid_alt.pid_preregZ0Z_6 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_5 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_6 ),
            .clk(N__87209),
            .ce(N__51492),
            .sr(N__79614));
    defparam \pid_alt.pid_prereg_esr_7_LC_3_16_0 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_7_LC_3_16_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_7_LC_3_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_7_LC_3_16_0  (
            .in0(_gnd_net_),
            .in1(N__35990),
            .in2(N__34338),
            .in3(N__34329),
            .lcout(\pid_alt.pid_preregZ0Z_7 ),
            .ltout(),
            .carryin(bfn_3_16_0_),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_7 ),
            .clk(N__87224),
            .ce(N__51489),
            .sr(N__79622));
    defparam \pid_alt.pid_prereg_esr_8_LC_3_16_1 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_8_LC_3_16_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_8_LC_3_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_8_LC_3_16_1  (
            .in0(_gnd_net_),
            .in1(N__34326),
            .in2(N__34320),
            .in3(N__34305),
            .lcout(\pid_alt.pid_preregZ0Z_8 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_7 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_8 ),
            .clk(N__87224),
            .ce(N__51489),
            .sr(N__79622));
    defparam \pid_alt.pid_prereg_esr_9_LC_3_16_2 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_9_LC_3_16_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_9_LC_3_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_9_LC_3_16_2  (
            .in0(_gnd_net_),
            .in1(N__34302),
            .in2(N__34496),
            .in3(N__34473),
            .lcout(\pid_alt.pid_preregZ0Z_9 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_8 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_9 ),
            .clk(N__87224),
            .ce(N__51489),
            .sr(N__79622));
    defparam \pid_alt.pid_prereg_esr_10_LC_3_16_3 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_10_LC_3_16_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_10_LC_3_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_10_LC_3_16_3  (
            .in0(_gnd_net_),
            .in1(N__34935),
            .in2(N__34962),
            .in3(N__34470),
            .lcout(\pid_alt.pid_preregZ0Z_10 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_9 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_10 ),
            .clk(N__87224),
            .ce(N__51489),
            .sr(N__79622));
    defparam \pid_alt.pid_prereg_esr_11_LC_3_16_4 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_11_LC_3_16_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_11_LC_3_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_11_LC_3_16_4  (
            .in0(_gnd_net_),
            .in1(N__34467),
            .in2(N__34901),
            .in3(N__34458),
            .lcout(\pid_alt.pid_preregZ0Z_11 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_10 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_11 ),
            .clk(N__87224),
            .ce(N__51489),
            .sr(N__79622));
    defparam \pid_alt.pid_prereg_esr_12_LC_3_16_5 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_12_LC_3_16_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_12_LC_3_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_12_LC_3_16_5  (
            .in0(_gnd_net_),
            .in1(N__38544),
            .in2(N__38606),
            .in3(N__34455),
            .lcout(\pid_alt.pid_preregZ0Z_12 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_11 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_12 ),
            .clk(N__87224),
            .ce(N__51489),
            .sr(N__79622));
    defparam \pid_alt.pid_prereg_esr_13_LC_3_16_6 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_13_LC_3_16_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_13_LC_3_16_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_13_LC_3_16_6  (
            .in0(_gnd_net_),
            .in1(N__38844),
            .in2(N__38682),
            .in3(N__34452),
            .lcout(\pid_alt.pid_preregZ0Z_13 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_12 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_13 ),
            .clk(N__87224),
            .ce(N__51489),
            .sr(N__79622));
    defparam \pid_alt.pid_prereg_esr_14_LC_3_16_7 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_14_LC_3_16_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_14_LC_3_16_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_14_LC_3_16_7  (
            .in0(_gnd_net_),
            .in1(N__36072),
            .in2(N__38802),
            .in3(N__34440),
            .lcout(\pid_alt.pid_preregZ0Z_14 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_13 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_14 ),
            .clk(N__87224),
            .ce(N__51489),
            .sr(N__79622));
    defparam \pid_alt.pid_prereg_esr_15_LC_3_17_0 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_15_LC_3_17_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_15_LC_3_17_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_15_LC_3_17_0  (
            .in0(_gnd_net_),
            .in1(N__36168),
            .in2(N__36347),
            .in3(N__34428),
            .lcout(\pid_alt.pid_preregZ0Z_15 ),
            .ltout(),
            .carryin(bfn_3_17_0_),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_15 ),
            .clk(N__87239),
            .ce(N__51485),
            .sr(N__79630));
    defparam \pid_alt.pid_prereg_esr_16_LC_3_17_1 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_16_LC_3_17_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_16_LC_3_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_16_LC_3_17_1  (
            .in0(_gnd_net_),
            .in1(N__35247),
            .in2(N__36119),
            .in3(N__34416),
            .lcout(\pid_alt.pid_preregZ0Z_16 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_15 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_16 ),
            .clk(N__87239),
            .ce(N__51485),
            .sr(N__79630));
    defparam \pid_alt.pid_prereg_esr_17_LC_3_17_2 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_17_LC_3_17_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_17_LC_3_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_17_LC_3_17_2  (
            .in0(_gnd_net_),
            .in1(N__35343),
            .in2(N__35355),
            .in3(N__34404),
            .lcout(\pid_alt.pid_preregZ0Z_17 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_16 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_17 ),
            .clk(N__87239),
            .ce(N__51485),
            .sr(N__79630));
    defparam \pid_alt.pid_prereg_esr_18_LC_3_17_3 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_18_LC_3_17_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_18_LC_3_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_18_LC_3_17_3  (
            .in0(_gnd_net_),
            .in1(N__34653),
            .in2(N__34878),
            .in3(N__34632),
            .lcout(\pid_alt.pid_preregZ0Z_18 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_17 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_18 ),
            .clk(N__87239),
            .ce(N__51485),
            .sr(N__79630));
    defparam \pid_alt.pid_prereg_esr_19_LC_3_17_4 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_19_LC_3_17_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_19_LC_3_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_19_LC_3_17_4  (
            .in0(_gnd_net_),
            .in1(N__34629),
            .in2(N__34617),
            .in3(N__34587),
            .lcout(\pid_alt.pid_preregZ0Z_19 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_18 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_19 ),
            .clk(N__87239),
            .ce(N__51485),
            .sr(N__79630));
    defparam \pid_alt.pid_prereg_esr_20_LC_3_17_5 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_20_LC_3_17_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_20_LC_3_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_20_LC_3_17_5  (
            .in0(_gnd_net_),
            .in1(N__34779),
            .in2(N__34803),
            .in3(N__34575),
            .lcout(\pid_alt.pid_preregZ0Z_20 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_19 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_20 ),
            .clk(N__87239),
            .ce(N__51485),
            .sr(N__79630));
    defparam \pid_alt.pid_prereg_esr_21_LC_3_17_6 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_21_LC_3_17_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_21_LC_3_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_21_LC_3_17_6  (
            .in0(_gnd_net_),
            .in1(N__34836),
            .in2(N__34740),
            .in3(N__34560),
            .lcout(\pid_alt.pid_preregZ0Z_21 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_20 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_21 ),
            .clk(N__87239),
            .ce(N__51485),
            .sr(N__79630));
    defparam \pid_alt.pid_prereg_esr_22_LC_3_17_7 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_22_LC_3_17_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_22_LC_3_17_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_22_LC_3_17_7  (
            .in0(_gnd_net_),
            .in1(N__34667),
            .in2(N__34680),
            .in3(N__34542),
            .lcout(\pid_alt.pid_preregZ0Z_22 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_21 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_22 ),
            .clk(N__87239),
            .ce(N__51485),
            .sr(N__79630));
    defparam \pid_alt.pid_prereg_esr_23_LC_3_18_0 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_23_LC_3_18_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_23_LC_3_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_23_LC_3_18_0  (
            .in0(_gnd_net_),
            .in1(N__34668),
            .in2(N__35034),
            .in3(N__34530),
            .lcout(\pid_alt.pid_preregZ0Z_23 ),
            .ltout(),
            .carryin(bfn_3_18_0_),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_23 ),
            .clk(N__87250),
            .ce(N__51482),
            .sr(N__79638));
    defparam \pid_alt.pid_prereg_esr_24_LC_3_18_1 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_24_LC_3_18_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_24_LC_3_18_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_alt.pid_prereg_esr_24_LC_3_18_1  (
            .in0(_gnd_net_),
            .in1(N__34527),
            .in2(_gnd_net_),
            .in3(N__34515),
            .lcout(\pid_alt.pid_preregZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87250),
            .ce(N__51482),
            .sr(N__79638));
    defparam \pid_alt.error_i_acumm_prereg_esr_7_LC_3_18_7 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_7_LC_3_18_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_7_LC_3_18_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_7_LC_3_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34512),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87250),
            .ce(N__51482),
            .sr(N__79638));
    defparam \pid_alt.error_d_reg_prev_esr_RNICG9B1_0_20_LC_3_19_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNICG9B1_0_20_LC_3_19_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNICG9B1_0_20_LC_3_19_0 .LUT_INIT=16'b0001100011100111;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNICG9B1_0_20_LC_3_19_0  (
            .in0(N__35140),
            .in1(N__35093),
            .in2(N__35181),
            .in3(N__35054),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNICG9B1_0Z0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI86IM_19_LC_3_19_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI86IM_19_LC_3_19_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI86IM_19_LC_3_19_1 .LUT_INIT=16'b1000100011101110;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI86IM_19_LC_3_19_1  (
            .in0(N__34727),
            .in1(N__34827),
            .in2(_gnd_net_),
            .in3(N__34694),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI86IMZ0Z_19 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNI86IMZ0Z_19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIK3024_19_LC_3_19_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIK3024_19_LC_3_19_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIK3024_19_LC_3_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIK3024_19_LC_3_19_2  (
            .in0(N__34802),
            .in1(N__34770),
            .in2(N__34782),
            .in3(N__34753),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIK3024Z0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIGGKM_20_LC_3_19_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIGGKM_20_LC_3_19_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIGGKM_20_LC_3_19_3 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIGGKM_20_LC_3_19_3  (
            .in0(N__35092),
            .in1(N__35173),
            .in2(_gnd_net_),
            .in3(N__35139),
            .lcout(\pid_alt.un1_pid_prereg_236_1 ),
            .ltout(\pid_alt.un1_pid_prereg_236_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIS5212_19_LC_3_19_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIS5212_19_LC_3_19_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIS5212_19_LC_3_19_4 .LUT_INIT=16'b1111110011000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIS5212_19_LC_3_19_4  (
            .in0(_gnd_net_),
            .in1(N__34764),
            .in2(N__34758),
            .in3(N__34754),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIS5212Z0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_20_LC_3_19_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_20_LC_3_19_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_20_LC_3_19_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_20_LC_3_19_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35151),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87255),
            .ce(N__51480),
            .sr(N__79646));
    defparam \pid_alt.error_d_reg_prev_esr_19_LC_3_19_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_19_LC_3_19_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_19_LC_3_19_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_19_LC_3_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34728),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87255),
            .ce(N__51480),
            .sr(N__79646));
    defparam \pid_alt.error_d_reg_prev_esr_RNICG9B1_1_20_LC_3_19_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNICG9B1_1_20_LC_3_19_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNICG9B1_1_20_LC_3_19_7 .LUT_INIT=16'b0110010101011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNICG9B1_1_20_LC_3_19_7  (
            .in0(N__35055),
            .in1(N__35177),
            .in2(N__35104),
            .in3(N__35141),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNICG9B1_1Z0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNICG9B1_20_LC_3_20_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNICG9B1_20_LC_3_20_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNICG9B1_20_LC_3_20_0 .LUT_INIT=16'b1111110101000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNICG9B1_20_LC_3_20_0  (
            .in0(N__35178),
            .in1(N__35142),
            .in2(N__35105),
            .in3(N__35056),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNICG9B1Z0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNICG9B1_2_20_LC_3_20_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNICG9B1_2_20_LC_3_20_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNICG9B1_2_20_LC_3_20_2 .LUT_INIT=16'b0100001010111101;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNICG9B1_2_20_LC_3_20_2  (
            .in0(N__35179),
            .in1(N__35143),
            .in2(N__35106),
            .in3(N__35057),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNICG9B1_2Z0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIL8611_9_LC_3_20_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIL8611_9_LC_3_20_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIL8611_9_LC_3_20_4 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIL8611_9_LC_3_20_4  (
            .in0(N__35022),
            .in1(N__35001),
            .in2(_gnd_net_),
            .in3(N__34986),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIL8611Z0Z_9 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNIL8611Z0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNICI045_9_LC_3_20_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNICI045_9_LC_3_20_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNICI045_9_LC_3_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNICI045_9_LC_3_20_5  (
            .in0(N__34958),
            .in1(N__34919),
            .in2(N__34938),
            .in3(N__37144),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNICI045Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI57T82_7_LC_3_20_6 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI57T82_7_LC_3_20_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI57T82_7_LC_3_20_6 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNI57T82_7_LC_3_20_6  (
            .in0(N__37247),
            .in1(N__48448),
            .in2(N__39556),
            .in3(N__36879),
            .lcout(\pid_alt.m21_e_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNISAR62_9_LC_3_20_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNISAR62_9_LC_3_20_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNISAR62_9_LC_3_20_7 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNISAR62_9_LC_3_20_7  (
            .in0(N__34926),
            .in1(N__34920),
            .in2(_gnd_net_),
            .in3(N__37145),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNISAR62Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_16_LC_3_21_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_16_LC_3_21_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_16_LC_3_21_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_16_LC_3_21_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35301),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87264),
            .ce(N__51477),
            .sr(N__79663));
    defparam \pid_alt.error_d_reg_prev_esr_RNI8BR02_16_LC_3_21_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI8BR02_16_LC_3_21_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI8BR02_16_LC_3_21_2 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI8BR02_16_LC_3_21_2  (
            .in0(N__34851),
            .in1(N__34845),
            .in2(_gnd_net_),
            .in3(N__35369),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI8BR02Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIVSHM_16_LC_3_21_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIVSHM_16_LC_3_21_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIVSHM_16_LC_3_21_3 .LUT_INIT=16'b1010111100001010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIVSHM_16_LC_3_21_3  (
            .in0(N__35300),
            .in1(_gnd_net_),
            .in2(N__35313),
            .in3(N__35328),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIVSHMZ0Z_16 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNIVSHMZ0Z_16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI8DL14_16_LC_3_21_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI8DL14_16_LC_3_21_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI8DL14_16_LC_3_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI8DL14_16_LC_3_21_4  (
            .in0(N__35342),
            .in1(N__34844),
            .in2(N__35373),
            .in3(N__35368),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI8DL14Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI02Q02_15_LC_3_21_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI02Q02_15_LC_3_21_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI02Q02_15_LC_3_21_5 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI02Q02_15_LC_3_21_5  (
            .in0(N__35274),
            .in1(N__51576),
            .in2(_gnd_net_),
            .in3(N__35261),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI02Q02Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIVSHM_0_16_LC_3_21_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIVSHM_0_16_LC_3_21_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIVSHM_0_16_LC_3_21_6 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIVSHM_0_16_LC_3_21_6  (
            .in0(N__35327),
            .in1(N__35309),
            .in2(_gnd_net_),
            .in3(N__35299),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIVSHM_0Z0Z_16 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNIVSHM_0Z0Z_16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIOQI14_15_LC_3_21_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIOQI14_15_LC_3_21_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIOQI14_15_LC_3_21_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIOQI14_15_LC_3_21_7  (
            .in0(N__36129),
            .in1(N__51575),
            .in2(N__35268),
            .in3(N__35260),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIOQI14Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_13_LC_3_22_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_13_LC_3_22_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_13_LC_3_22_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_13_LC_3_22_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38736),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87269),
            .ce(N__51474),
            .sr(N__79671));
    defparam \pid_alt.error_i_acumm_prereg_esr_6_LC_3_22_3 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_6_LC_3_22_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_6_LC_3_22_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_6_LC_3_22_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35886),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87269),
            .ce(N__51474),
            .sr(N__79671));
    defparam \pid_alt.error_i_acumm_prereg_esr_4_LC_3_22_4 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_4_LC_3_22_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_4_LC_3_22_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_4_LC_3_22_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35238),
            .lcout(\pid_alt.error_i_acumm7lto4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87269),
            .ce(N__51474),
            .sr(N__79671));
    defparam \pid_alt.error_i_acumm_prereg_esr_13_LC_3_22_5 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_13_LC_3_22_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_13_LC_3_22_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_13_LC_3_22_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38827),
            .lcout(\pid_alt.error_i_acumm7lto13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87269),
            .ce(N__51474),
            .sr(N__79671));
    defparam \pid_alt.error_i_acumm_prereg_esr_2_LC_3_22_6 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_2_LC_3_22_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_2_LC_3_22_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_2_LC_3_22_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35213),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87269),
            .ce(N__51474),
            .sr(N__79671));
    defparam \pid_alt.error_i_acumm_prereg_esr_15_LC_3_22_7 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_15_LC_3_22_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_15_LC_3_22_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_15_LC_3_22_7  (
            .in0(N__36151),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87269),
            .ce(N__51474),
            .sr(N__79671));
    defparam \pid_alt.error_i_acumm_prereg_esr_3_LC_3_23_1 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_3_LC_3_23_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_3_LC_3_23_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_3_LC_3_23_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35420),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87274),
            .ce(N__51473),
            .sr(N__79677));
    defparam \pid_alt.source_pid_1_esr_13_LC_4_9_5 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_esr_13_LC_4_9_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_esr_13_LC_4_9_5 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \pid_alt.source_pid_1_esr_13_LC_4_9_5  (
            .in0(N__37717),
            .in1(N__37631),
            .in2(_gnd_net_),
            .in3(N__37775),
            .lcout(throttle_order_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87100),
            .ce(N__35525),
            .sr(N__37813));
    defparam \pid_alt.source_pid_1_esr_12_LC_4_9_6 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_esr_12_LC_4_9_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_esr_12_LC_4_9_6 .LUT_INIT=16'b1111010000000000;
    LogicCell40 \pid_alt.source_pid_1_esr_12_LC_4_9_6  (
            .in0(N__37774),
            .in1(N__37718),
            .in2(N__37642),
            .in3(N__37548),
            .lcout(throttle_order_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87100),
            .ce(N__35525),
            .sr(N__37813));
    defparam \pid_alt.pid_prereg_esr_RNI3A6GE_13_LC_4_10_0 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNI3A6GE_13_LC_4_10_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNI3A6GE_13_LC_4_10_0 .LUT_INIT=16'b0010000011111111;
    LogicCell40 \pid_alt.pid_prereg_esr_RNI3A6GE_13_LC_4_10_0  (
            .in0(N__37713),
            .in1(N__37759),
            .in2(N__35610),
            .in3(N__35616),
            .lcout(\pid_alt.un1_reset_0_i ),
            .ltout(\pid_alt.un1_reset_0_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.state_RNIOVDUE_1_LC_4_10_1 .C_ON=1'b0;
    defparam \pid_alt.state_RNIOVDUE_1_LC_4_10_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.state_RNIOVDUE_1_LC_4_10_1 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \pid_alt.state_RNIOVDUE_1_LC_4_10_1  (
            .in0(N__65399),
            .in1(_gnd_net_),
            .in2(N__35388),
            .in3(_gnd_net_),
            .lcout(\pid_alt.N_72_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNIP29I1_4_LC_4_10_2 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNIP29I1_4_LC_4_10_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNIP29I1_4_LC_4_10_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \pid_alt.pid_prereg_esr_RNIP29I1_4_LC_4_10_2  (
            .in0(N__35578),
            .in1(N__65397),
            .in2(N__37770),
            .in3(N__35641),
            .lcout(\pid_alt.source_pid_1_sqmuxa_0_a2_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNIIM6H1_6_LC_4_10_3 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNIIM6H1_6_LC_4_10_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNIIM6H1_6_LC_4_10_3 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \pid_alt.pid_prereg_esr_RNIIM6H1_6_LC_4_10_3  (
            .in0(N__37901),
            .in1(N__37931),
            .in2(N__37873),
            .in3(N__37961),
            .lcout(),
            .ltout(\pid_alt.source_pid_1_sqmuxa_0_o2_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNIFQKS1_10_LC_4_10_4 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNIFQKS1_10_LC_4_10_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNIFQKS1_10_LC_4_10_4 .LUT_INIT=16'b1111001111111111;
    LogicCell40 \pid_alt.pid_prereg_esr_RNIFQKS1_10_LC_4_10_4  (
            .in0(_gnd_net_),
            .in1(N__37458),
            .in2(N__35385),
            .in3(N__37493),
            .lcout(\pid_alt.N_51 ),
            .ltout(\pid_alt.N_51_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNIVVFP6_4_LC_4_10_5 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNIVVFP6_4_LC_4_10_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNIVVFP6_4_LC_4_10_5 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \pid_alt.pid_prereg_esr_RNIVVFP6_4_LC_4_10_5  (
            .in0(N__35693),
            .in1(N__37712),
            .in2(N__35382),
            .in3(N__35379),
            .lcout(),
            .ltout(\pid_alt.N_57_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNI4AMM7_24_LC_4_10_6 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNI4AMM7_24_LC_4_10_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNI4AMM7_24_LC_4_10_6 .LUT_INIT=16'b0000000000000111;
    LogicCell40 \pid_alt.pid_prereg_esr_RNI4AMM7_24_LC_4_10_6  (
            .in0(N__37630),
            .in1(N__65398),
            .in2(N__35619),
            .in3(N__65987),
            .lcout(\pid_alt.un1_reset_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNIHMCQ4_4_LC_4_10_7 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNIHMCQ4_4_LC_4_10_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNIHMCQ4_4_LC_4_10_7 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \pid_alt.pid_prereg_esr_RNIHMCQ4_4_LC_4_10_7  (
            .in0(N__35642),
            .in1(N__37467),
            .in2(N__35697),
            .in3(N__35579),
            .lcout(\pid_alt.source_pid_1_sqmuxa_0_a2_1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNIG2382_12_LC_4_11_1 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNIG2382_12_LC_4_11_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNIG2382_12_LC_4_11_1 .LUT_INIT=16'b0011001110111011;
    LogicCell40 \pid_alt.pid_prereg_esr_RNIG2382_12_LC_4_11_1  (
            .in0(N__35601),
            .in1(N__37760),
            .in2(_gnd_net_),
            .in3(N__37546),
            .lcout(\pid_alt.N_52 ),
            .ltout(\pid_alt.N_52_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNI3BD63_4_LC_4_11_2 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNI3BD63_4_LC_4_11_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNI3BD63_4_LC_4_11_2 .LUT_INIT=16'b1111010111110000;
    LogicCell40 \pid_alt.pid_prereg_esr_RNI3BD63_4_LC_4_11_2  (
            .in0(N__35580),
            .in1(_gnd_net_),
            .in2(N__35550),
            .in3(N__35643),
            .lcout(\pid_alt.N_54 ),
            .ltout(\pid_alt.N_54_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.source_pid_1_esr_0_LC_4_11_3 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_esr_0_LC_4_11_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_esr_0_LC_4_11_3 .LUT_INIT=16'b1100100010001000;
    LogicCell40 \pid_alt.source_pid_1_esr_0_LC_4_11_3  (
            .in0(N__37618),
            .in1(N__35445),
            .in2(N__35547),
            .in3(N__37710),
            .lcout(throttle_order_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87131),
            .ce(N__35524),
            .sr(N__37812));
    defparam \pid_alt.source_pid_1_esr_1_LC_4_11_4 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_esr_1_LC_4_11_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_esr_1_LC_4_11_4 .LUT_INIT=16'b1110000011000000;
    LogicCell40 \pid_alt.source_pid_1_esr_1_LC_4_11_4  (
            .in0(N__37708),
            .in1(N__37619),
            .in2(N__35481),
            .in3(N__35539),
            .lcout(throttle_order_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87131),
            .ce(N__35524),
            .sr(N__37812));
    defparam \pid_alt.source_pid_1_esr_2_LC_4_11_5 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_esr_2_LC_4_11_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_esr_2_LC_4_11_5 .LUT_INIT=16'b1010100010001000;
    LogicCell40 \pid_alt.source_pid_1_esr_2_LC_4_11_5  (
            .in0(N__35496),
            .in1(N__37638),
            .in2(N__35544),
            .in3(N__37711),
            .lcout(throttle_order_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87131),
            .ce(N__35524),
            .sr(N__37812));
    defparam \pid_alt.source_pid_1_esr_3_LC_4_11_6 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_esr_3_LC_4_11_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_esr_3_LC_4_11_6 .LUT_INIT=16'b1111100000000000;
    LogicCell40 \pid_alt.source_pid_1_esr_3_LC_4_11_6  (
            .in0(N__37709),
            .in1(N__35543),
            .in2(N__37646),
            .in3(N__35462),
            .lcout(throttle_order_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87131),
            .ce(N__35524),
            .sr(N__37812));
    defparam \pid_alt.pid_prereg_esr_RNIQT5H1_0_LC_4_11_7 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNIQT5H1_0_LC_4_11_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNIQT5H1_0_LC_4_11_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_alt.pid_prereg_esr_RNIQT5H1_0_LC_4_11_7  (
            .in0(N__35495),
            .in1(N__35477),
            .in2(N__35463),
            .in3(N__35444),
            .lcout(\pid_alt.source_pid_1_sqmuxa_0_a2_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_5_LC_4_12_0 .C_ON=1'b0;
    defparam \uart_pc.data_5_LC_4_12_0 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_5_LC_4_12_0 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \uart_pc.data_5_LC_4_12_0  (
            .in0(N__35780),
            .in1(N__35756),
            .in2(N__73590),
            .in3(N__37980),
            .lcout(uart_pc_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87149),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_2_LC_4_12_1 .C_ON=1'b0;
    defparam \uart_pc.data_2_LC_4_12_1 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_2_LC_4_12_1 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \uart_pc.data_2_LC_4_12_1  (
            .in0(N__35754),
            .in1(N__35778),
            .in2(N__77527),
            .in3(N__38078),
            .lcout(uart_pc_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87149),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_3_LC_4_12_2 .C_ON=1'b0;
    defparam \uart_pc.data_3_LC_4_12_2 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_3_LC_4_12_2 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \uart_pc.data_3_LC_4_12_2  (
            .in0(N__35779),
            .in1(N__35755),
            .in2(N__38058),
            .in3(N__83938),
            .lcout(uart_pc_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87149),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_ns_0_a3_0_1_2_LC_4_12_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_ns_0_a3_0_1_2_LC_4_12_3 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_ns_0_a3_0_1_2_LC_4_12_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \Commands_frame_decoder.state_ns_0_a3_0_1_2_LC_4_12_3  (
            .in0(_gnd_net_),
            .in1(N__85097),
            .in2(_gnd_net_),
            .in3(N__77459),
            .lcout(\Commands_frame_decoder.state_ns_0_a3_0_1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_0_LC_4_12_5 .C_ON=1'b0;
    defparam \uart_pc.data_0_LC_4_12_5 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_0_LC_4_12_5 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \uart_pc.data_0_LC_4_12_5  (
            .in0(N__35751),
            .in1(N__35773),
            .in2(N__38127),
            .in3(N__83755),
            .lcout(uart_pc_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87149),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_1_4_LC_4_12_6 .C_ON=1'b0;
    defparam \uart_pc.data_1_4_LC_4_12_6 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_1_4_LC_4_12_6 .LUT_INIT=16'b0000101011001010;
    LogicCell40 \uart_pc.data_1_4_LC_4_12_6  (
            .in0(N__85098),
            .in1(N__38007),
            .in2(N__35781),
            .in3(N__35752),
            .lcout(uart_pc_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87149),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_1_LC_4_12_7 .C_ON=1'b0;
    defparam \uart_pc.data_1_LC_4_12_7 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_1_LC_4_12_7 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \uart_pc.data_1_LC_4_12_7  (
            .in0(N__35753),
            .in1(N__35777),
            .in2(N__38103),
            .in3(N__84123),
            .lcout(uart_pc_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87149),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNIE28S_5_LC_4_13_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIE28S_5_LC_4_13_0 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIE28S_5_LC_4_13_0 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \Commands_frame_decoder.state_RNIE28S_5_LC_4_13_0  (
            .in0(N__79946),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35678),
            .lcout(\Commands_frame_decoder.source_CH4data_1_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNIIM0I_5_LC_4_13_1 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNIIM0I_5_LC_4_13_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNIIM0I_5_LC_4_13_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \pid_alt.pid_prereg_esr_RNIIM0I_5_LC_4_13_1  (
            .in0(_gnd_net_),
            .in1(N__37536),
            .in2(_gnd_net_),
            .in3(N__35660),
            .lcout(\pid_alt.N_154 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNILR1B2_2_LC_4_13_2 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_RNILR1B2_2_LC_4_13_2 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNILR1B2_2_LC_4_13_2 .LUT_INIT=16'b1011101110101010;
    LogicCell40 \uart_pc.timer_Count_RNILR1B2_2_LC_4_13_2  (
            .in0(N__79945),
            .in1(N__40205),
            .in2(_gnd_net_),
            .in3(N__38151),
            .lcout(\uart_pc.timer_Count_RNILR1B2Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNIMQ8T1_2_LC_4_13_3 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_RNIMQ8T1_2_LC_4_13_3 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNIMQ8T1_2_LC_4_13_3 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \uart_pc.timer_Count_RNIMQ8T1_2_LC_4_13_3  (
            .in0(N__38152),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79947),
            .lcout(\uart_pc.timer_Count_RNIMQ8T1Z0Z_2 ),
            .ltout(\uart_pc.timer_Count_RNIMQ8T1Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_6_LC_4_13_4 .C_ON=1'b0;
    defparam \uart_pc.data_6_LC_4_13_4 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_6_LC_4_13_4 .LUT_INIT=16'b0010111100100000;
    LogicCell40 \uart_pc.data_6_LC_4_13_4  (
            .in0(N__38256),
            .in1(N__35750),
            .in2(N__35721),
            .in3(N__85308),
            .lcout(uart_pc_data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87165),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNIF38S_6_LC_4_13_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIF38S_6_LC_4_13_7 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIF38S_6_LC_4_13_7 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \Commands_frame_decoder.state_RNIF38S_6_LC_4_13_7  (
            .in0(N__38202),
            .in1(N__38374),
            .in2(_gnd_net_),
            .in3(N__79944),
            .lcout(\Commands_frame_decoder.state_RNIF38SZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_CH1data_3_LC_4_14_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH1data_3_LC_4_14_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH1data_3_LC_4_14_0 .LUT_INIT=16'b0010111100100000;
    LogicCell40 \Commands_frame_decoder.source_CH1data_3_LC_4_14_0  (
            .in0(N__83947),
            .in1(N__35711),
            .in2(N__38511),
            .in3(N__36557),
            .lcout(alt_command_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87179),
            .ce(),
            .sr(N__79604));
    defparam \Commands_frame_decoder.source_CH1data_1_LC_4_14_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH1data_1_LC_4_14_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH1data_1_LC_4_14_1 .LUT_INIT=16'b0100111101000000;
    LogicCell40 \Commands_frame_decoder.source_CH1data_1_LC_4_14_1  (
            .in0(N__35707),
            .in1(N__84132),
            .in2(N__38510),
            .in3(N__36692),
            .lcout(alt_command_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87179),
            .ce(),
            .sr(N__79604));
    defparam \Commands_frame_decoder.source_CH1data8lto7_2_LC_4_14_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH1data8lto7_2_LC_4_14_2 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.source_CH1data8lto7_2_LC_4_14_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \Commands_frame_decoder.source_CH1data8lto7_2_LC_4_14_2  (
            .in0(N__85288),
            .in1(N__73579),
            .in2(N__85029),
            .in3(N__85131),
            .lcout(),
            .ltout(\Commands_frame_decoder.source_CH1data8lto7Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_CH1data8lto7_LC_4_14_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH1data8lto7_LC_4_14_3 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.source_CH1data8lto7_LC_4_14_3 .LUT_INIT=16'b0001000011110000;
    LogicCell40 \Commands_frame_decoder.source_CH1data8lto7_LC_4_14_3  (
            .in0(N__77499),
            .in1(N__84131),
            .in2(N__35718),
            .in3(N__83946),
            .lcout(\Commands_frame_decoder.source_CH1data8 ),
            .ltout(\Commands_frame_decoder.source_CH1data8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_CH1data_0_LC_4_14_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH1data_0_LC_4_14_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH1data_0_LC_4_14_4 .LUT_INIT=16'b0011101100001000;
    LogicCell40 \Commands_frame_decoder.source_CH1data_0_LC_4_14_4  (
            .in0(N__83757),
            .in1(N__38502),
            .in2(N__35715),
            .in3(N__36755),
            .lcout(alt_command_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87179),
            .ce(),
            .sr(N__79604));
    defparam \Commands_frame_decoder.source_CH1data_2_LC_4_14_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH1data_2_LC_4_14_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH1data_2_LC_4_14_5 .LUT_INIT=16'b0011101100001000;
    LogicCell40 \Commands_frame_decoder.source_CH1data_2_LC_4_14_5  (
            .in0(N__77500),
            .in1(N__38506),
            .in2(N__35712),
            .in3(N__36626),
            .lcout(alt_command_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87179),
            .ce(),
            .sr(N__79604));
    defparam \Commands_frame_decoder.state_RNO_2_0_LC_4_14_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNO_2_0_LC_4_14_6 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNO_2_0_LC_4_14_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Commands_frame_decoder.state_RNO_2_0_LC_4_14_6  (
            .in0(N__83756),
            .in1(N__85130),
            .in2(N__85321),
            .in3(N__77498),
            .lcout(\Commands_frame_decoder.state_ns_i_a2_0_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_5_LC_4_15_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_5_LC_4_15_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_5_LC_4_15_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_5_LC_4_15_0  (
            .in0(N__35838),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87193),
            .ce(N__51490),
            .sr(N__79608));
    defparam \pid_alt.error_d_reg_prev_esr_RNI9S511_5_LC_4_15_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI9S511_5_LC_4_15_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI9S511_5_LC_4_15_1 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI9S511_5_LC_4_15_1  (
            .in0(N__35804),
            .in1(N__35813),
            .in2(_gnd_net_),
            .in3(N__35836),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI9S511Z0Z_5 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNI9S511Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIL81T2_5_LC_4_15_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIL81T2_5_LC_4_15_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIL81T2_5_LC_4_15_2 .LUT_INIT=16'b1111110011000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIL81T2_5_LC_4_15_2  (
            .in0(_gnd_net_),
            .in1(N__35901),
            .in2(N__36000),
            .in3(N__35885),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIL81T2Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNICV511_0_6_LC_4_15_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNICV511_0_6_LC_4_15_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNICV511_0_6_LC_4_15_3 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNICV511_0_6_LC_4_15_3  (
            .in0(N__35978),
            .in1(N__35955),
            .in2(_gnd_net_),
            .in3(N__35937),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNICV511_0Z0Z_6 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNICV511_0Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI171A6_5_LC_4_15_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI171A6_5_LC_4_15_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI171A6_5_LC_4_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI171A6_5_LC_4_15_4  (
            .in0(N__35852),
            .in1(N__35895),
            .in2(N__35889),
            .in3(N__35884),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI171A6Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNICUVC3_4_LC_4_15_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNICUVC3_4_LC_4_15_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNICUVC3_4_LC_4_15_5 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNICUVC3_4_LC_4_15_5  (
            .in0(N__35787),
            .in1(N__36198),
            .in2(_gnd_net_),
            .in3(N__37202),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNICUVC3Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI9S511_0_5_LC_4_15_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI9S511_0_5_LC_4_15_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI9S511_0_5_LC_4_15_6 .LUT_INIT=16'b0101101010100101;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI9S511_0_5_LC_4_15_6  (
            .in0(N__35837),
            .in1(_gnd_net_),
            .in2(N__35817),
            .in3(N__35805),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI9S511_0Z0Z_5 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNI9S511_0Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIOGSO6_4_LC_4_15_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIOGSO6_4_LC_4_15_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIOGSO6_4_LC_4_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIOGSO6_4_LC_4_15_7  (
            .in0(N__36216),
            .in1(N__36197),
            .in2(N__36180),
            .in3(N__37201),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIOGSO6Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI88G14_14_LC_4_16_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI88G14_14_LC_4_16_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI88G14_14_LC_4_16_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI88G14_14_LC_4_16_0  (
            .in0(N__36101),
            .in1(N__36162),
            .in2(N__36348),
            .in3(N__36152),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI88G14Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIPMHM_14_LC_4_16_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIPMHM_14_LC_4_16_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIPMHM_14_LC_4_16_1 .LUT_INIT=16'b1010111100001010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIPMHM_14_LC_4_16_1  (
            .in0(N__36065),
            .in1(_gnd_net_),
            .in2(N__36045),
            .in3(N__36093),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIPMHMZ0Z_14 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNIPMHMZ0Z_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIOOO02_14_LC_4_16_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIOOO02_14_LC_4_16_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIOOO02_14_LC_4_16_2 .LUT_INIT=16'b1111101010100000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIOOO02_14_LC_4_16_2  (
            .in0(N__36102),
            .in1(_gnd_net_),
            .in2(N__36156),
            .in3(N__36153),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIOOO02Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNISPHM_0_15_LC_4_16_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNISPHM_0_15_LC_4_16_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNISPHM_0_15_LC_4_16_3 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNISPHM_0_15_LC_4_16_3  (
            .in0(N__51605),
            .in1(N__51516),
            .in2(_gnd_net_),
            .in3(N__51553),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNISPHM_0Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIPMHM_0_14_LC_4_16_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIPMHM_0_14_LC_4_16_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIPMHM_0_14_LC_4_16_4 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIPMHM_0_14_LC_4_16_4  (
            .in0(N__36092),
            .in1(N__36041),
            .in2(_gnd_net_),
            .in3(N__36064),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIPMHM_0Z0Z_14 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNIPMHM_0Z0Z_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNICQF44_13_LC_4_16_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNICQF44_13_LC_4_16_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNICQF44_13_LC_4_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNICQF44_13_LC_4_16_5  (
            .in0(N__38798),
            .in1(N__36026),
            .in2(N__36075),
            .in3(N__36371),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNICQF44Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_14_LC_4_16_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_14_LC_4_16_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_14_LC_4_16_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_14_LC_4_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36066),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87210),
            .ce(N__51486),
            .sr(N__79615));
    defparam \pid_alt.error_d_reg_prev_esr_RNIGFN02_13_LC_4_16_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIGFN02_13_LC_4_16_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIGFN02_13_LC_4_16_7 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIGFN02_13_LC_4_16_7  (
            .in0(N__36033),
            .in1(N__36027),
            .in2(_gnd_net_),
            .in3(N__36372),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIGFN02Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_axb_1_LC_4_17_2 .C_ON=1'b0;
    defparam \pid_alt.error_axb_1_LC_4_17_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_axb_1_LC_4_17_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_alt.error_axb_1_LC_4_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38874),
            .lcout(\pid_alt.error_axbZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNIVT8S_2_LC_4_17_3 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_RNIVT8S_2_LC_4_17_3 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNIVT8S_2_LC_4_17_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uart_pc.timer_Count_RNIVT8S_2_LC_4_17_3  (
            .in0(_gnd_net_),
            .in1(N__40322),
            .in2(_gnd_net_),
            .in3(N__40443),
            .lcout(\uart_pc.N_126_li ),
            .ltout(\uart_pc.N_126_li_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_RNIMQ8T1_4_LC_4_17_4 .C_ON=1'b0;
    defparam \uart_pc.state_RNIMQ8T1_4_LC_4_17_4 .SEQ_MODE=4'b0000;
    defparam \uart_pc.state_RNIMQ8T1_4_LC_4_17_4 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \uart_pc.state_RNIMQ8T1_4_LC_4_17_4  (
            .in0(N__40551),
            .in1(N__40386),
            .in2(N__36330),
            .in3(N__79942),
            .lcout(\uart_pc.N_143 ),
            .ltout(\uart_pc.N_143_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_1_LC_4_17_5 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_1_LC_4_17_5 .SEQ_MODE=4'b1000;
    defparam \uart_pc.timer_Count_1_LC_4_17_5 .LUT_INIT=16'b0101010000000000;
    LogicCell40 \uart_pc.timer_Count_1_LC_4_17_5  (
            .in0(N__79943),
            .in1(N__41919),
            .in2(N__36327),
            .in3(N__36324),
            .lcout(\uart_pc.timer_CountZ1Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87225),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_0_c_inv_LC_4_17_6 .C_ON=1'b0;
    defparam \pid_alt.error_cry_0_c_inv_LC_4_17_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_0_c_inv_LC_4_17_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_alt.error_cry_0_c_inv_LC_4_17_6  (
            .in0(N__36318),
            .in1(N__56484),
            .in2(_gnd_net_),
            .in3(N__38890),
            .lcout(\pid_alt.drone_altitude_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNO_0_1_LC_4_17_7 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_RNO_0_1_LC_4_17_7 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNO_0_1_LC_4_17_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart_pc.timer_Count_RNO_0_1_LC_4_17_7  (
            .in0(_gnd_net_),
            .in1(N__41877),
            .in2(_gnd_net_),
            .in3(N__40085),
            .lcout(\uart_pc.timer_Count_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_0_c_LC_4_18_0 .C_ON=1'b1;
    defparam \pid_alt.error_cry_0_c_LC_4_18_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_0_c_LC_4_18_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_alt.error_cry_0_c_LC_4_18_0  (
            .in0(_gnd_net_),
            .in1(N__36317),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_18_0_),
            .carryout(\pid_alt.error_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_0_c_RNI1N2F_LC_4_18_1 .C_ON=1'b1;
    defparam \pid_alt.error_cry_0_c_RNI1N2F_LC_4_18_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_0_c_RNI1N2F_LC_4_18_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_cry_0_c_RNI1N2F_LC_4_18_1  (
            .in0(_gnd_net_),
            .in1(N__36306),
            .in2(_gnd_net_),
            .in3(N__36258),
            .lcout(\pid_alt.error_1 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_0 ),
            .carryout(\pid_alt.error_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_1_c_RNI3Q3F_LC_4_18_2 .C_ON=1'b1;
    defparam \pid_alt.error_cry_1_c_RNI3Q3F_LC_4_18_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_1_c_RNI3Q3F_LC_4_18_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_cry_1_c_RNI3Q3F_LC_4_18_2  (
            .in0(_gnd_net_),
            .in1(N__54165),
            .in2(_gnd_net_),
            .in3(N__36810),
            .lcout(\pid_alt.error_2 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_1 ),
            .carryout(\pid_alt.error_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_2_c_RNI5T4F_LC_4_18_3 .C_ON=1'b1;
    defparam \pid_alt.error_cry_2_c_RNI5T4F_LC_4_18_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_2_c_RNI5T4F_LC_4_18_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_cry_2_c_RNI5T4F_LC_4_18_3  (
            .in0(_gnd_net_),
            .in1(N__54147),
            .in2(_gnd_net_),
            .in3(N__36762),
            .lcout(\pid_alt.error_3 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_2 ),
            .carryout(\pid_alt.error_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_3_c_RNIKE1T_LC_4_18_4 .C_ON=1'b1;
    defparam \pid_alt.error_cry_3_c_RNIKE1T_LC_4_18_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_3_c_RNIKE1T_LC_4_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_cry_3_c_RNIKE1T_LC_4_18_4  (
            .in0(_gnd_net_),
            .in1(N__38862),
            .in2(N__36759),
            .in3(N__36702),
            .lcout(\pid_alt.error_4 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_3 ),
            .carryout(\pid_alt.error_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_4_c_RNINI2T_LC_4_18_5 .C_ON=1'b1;
    defparam \pid_alt.error_cry_4_c_RNINI2T_LC_4_18_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_4_c_RNINI2T_LC_4_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_cry_4_c_RNINI2T_LC_4_18_5  (
            .in0(_gnd_net_),
            .in1(N__38850),
            .in2(N__36699),
            .in3(N__36633),
            .lcout(\pid_alt.error_5 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_4 ),
            .carryout(\pid_alt.error_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_5_c_RNIQM3T_LC_4_18_6 .C_ON=1'b1;
    defparam \pid_alt.error_cry_5_c_RNIQM3T_LC_4_18_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_5_c_RNIQM3T_LC_4_18_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_cry_5_c_RNIQM3T_LC_4_18_6  (
            .in0(_gnd_net_),
            .in1(N__39024),
            .in2(N__36630),
            .in3(N__36567),
            .lcout(\pid_alt.error_6 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_5 ),
            .carryout(\pid_alt.error_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_6_c_RNITQ4T_LC_4_18_7 .C_ON=1'b1;
    defparam \pid_alt.error_cry_6_c_RNITQ4T_LC_4_18_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_6_c_RNITQ4T_LC_4_18_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_cry_6_c_RNITQ4T_LC_4_18_7  (
            .in0(_gnd_net_),
            .in1(N__39012),
            .in2(N__36564),
            .in3(N__36501),
            .lcout(\pid_alt.error_7 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_6 ),
            .carryout(\pid_alt.error_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_7_c_RNI9LEM_LC_4_19_0 .C_ON=1'b1;
    defparam \pid_alt.error_cry_7_c_RNI9LEM_LC_4_19_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_7_c_RNI9LEM_LC_4_19_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_cry_7_c_RNI9LEM_LC_4_19_0  (
            .in0(_gnd_net_),
            .in1(N__39006),
            .in2(N__39141),
            .in3(N__36465),
            .lcout(\pid_alt.error_8 ),
            .ltout(),
            .carryin(bfn_4_19_0_),
            .carryout(\pid_alt.error_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_8_c_RNICPFM_LC_4_19_1 .C_ON=1'b1;
    defparam \pid_alt.error_cry_8_c_RNICPFM_LC_4_19_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_8_c_RNICPFM_LC_4_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_cry_8_c_RNICPFM_LC_4_19_1  (
            .in0(_gnd_net_),
            .in1(N__39000),
            .in2(N__39132),
            .in3(N__36420),
            .lcout(\pid_alt.error_9 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_8 ),
            .carryout(\pid_alt.error_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_9_c_RNIMMUJ_LC_4_19_2 .C_ON=1'b1;
    defparam \pid_alt.error_cry_9_c_RNIMMUJ_LC_4_19_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_9_c_RNIMMUJ_LC_4_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_cry_9_c_RNIMMUJ_LC_4_19_2  (
            .in0(_gnd_net_),
            .in1(N__39147),
            .in2(N__39123),
            .in3(N__36375),
            .lcout(\pid_alt.error_10 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_9 ),
            .carryout(\pid_alt.error_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_10_c_RNI0SDO_LC_4_19_3 .C_ON=1'b1;
    defparam \pid_alt.error_cry_10_c_RNI0SDO_LC_4_19_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_10_c_RNI0SDO_LC_4_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_cry_10_c_RNI0SDO_LC_4_19_3  (
            .in0(_gnd_net_),
            .in1(N__54315),
            .in2(N__39114),
            .in3(N__37065),
            .lcout(\pid_alt.error_11 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_10 ),
            .carryout(\pid_alt.error_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_11_c_RNI5JAH_LC_4_19_4 .C_ON=1'b1;
    defparam \pid_alt.error_cry_11_c_RNI5JAH_LC_4_19_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_11_c_RNI5JAH_LC_4_19_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pid_alt.error_cry_11_c_RNI5JAH_LC_4_19_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__40629),
            .in3(N__37017),
            .lcout(\pid_alt.error_12 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_11 ),
            .carryout(\pid_alt.error_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_12_c_RNI7MBH_LC_4_19_5 .C_ON=1'b1;
    defparam \pid_alt.error_cry_12_c_RNI7MBH_LC_4_19_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_12_c_RNI7MBH_LC_4_19_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_cry_12_c_RNI7MBH_LC_4_19_5  (
            .in0(_gnd_net_),
            .in1(N__40614),
            .in2(_gnd_net_),
            .in3(N__36969),
            .lcout(\pid_alt.error_13 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_12 ),
            .carryout(\pid_alt.error_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_13_c_RNI9PCH_LC_4_19_6 .C_ON=1'b1;
    defparam \pid_alt.error_cry_13_c_RNI9PCH_LC_4_19_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_13_c_RNI9PCH_LC_4_19_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_cry_13_c_RNI9PCH_LC_4_19_6  (
            .in0(_gnd_net_),
            .in1(N__40602),
            .in2(_gnd_net_),
            .in3(N__36927),
            .lcout(\pid_alt.error_14 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_13 ),
            .carryout(\pid_alt.error_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_14_c_RNIBSDH_LC_4_19_7 .C_ON=1'b0;
    defparam \pid_alt.error_cry_14_c_RNIBSDH_LC_4_19_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_14_c_RNIBSDH_LC_4_19_7 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \pid_alt.error_cry_14_c_RNIBSDH_LC_4_19_7  (
            .in0(N__40665),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36924),
            .lcout(\pid_alt.error_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI935T_0_LC_4_20_1 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI935T_0_LC_4_20_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI935T_0_LC_4_20_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNI935T_0_LC_4_20_1  (
            .in0(_gnd_net_),
            .in1(N__37382),
            .in2(_gnd_net_),
            .in3(N__37322),
            .lcout(\pid_alt.m21_e_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_1_LC_4_20_2 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_1_LC_4_20_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_1_LC_4_20_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_1_LC_4_20_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36873),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87256),
            .ce(N__51478),
            .sr(N__79647));
    defparam \pid_alt.error_i_acumm_prereg_esr_0_LC_4_20_3 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_0_LC_4_20_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_0_LC_4_20_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_0_LC_4_20_3  (
            .in0(N__37310),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36840),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87256),
            .ce(N__51478),
            .sr(N__79647));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNILF5T_6_LC_4_20_4 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNILF5T_6_LC_4_20_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNILF5T_6_LC_4_20_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNILF5T_6_LC_4_20_4  (
            .in0(_gnd_net_),
            .in1(N__39557),
            .in2(_gnd_net_),
            .in3(N__39604),
            .lcout(\pid_alt.m35_e_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_5_LC_4_20_7 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_5_LC_4_20_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_5_LC_4_20_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_5_LC_4_20_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37203),
            .lcout(\pid_alt.error_i_acumm7lto5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87256),
            .ce(N__51478),
            .sr(N__79647));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI4CCV_10_LC_4_21_0 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI4CCV_10_LC_4_21_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI4CCV_10_LC_4_21_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNI4CCV_10_LC_4_21_0  (
            .in0(N__39095),
            .in1(N__39410),
            .in2(N__39059),
            .in3(N__39499),
            .lcout(\pid_alt.m35_e_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_8_LC_4_21_1 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_8_LC_4_21_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_8_LC_4_21_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_8_LC_4_21_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37176),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87260),
            .ce(N__51475),
            .sr(N__79654));
    defparam \pid_alt.error_i_acumm_prereg_esr_10_LC_4_21_2 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_10_LC_4_21_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_10_LC_4_21_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_10_LC_4_21_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37152),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87260),
            .ce(N__51475),
            .sr(N__79654));
    defparam \pid_alt.error_i_acumm_prereg_esr_12_LC_4_21_3 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_12_LC_4_21_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_12_LC_4_21_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_12_LC_4_21_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38571),
            .lcout(\pid_alt.error_i_acumm7lto12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87260),
            .ce(N__51475),
            .sr(N__79654));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNICP62_10_LC_4_21_4 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNICP62_10_LC_4_21_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNICP62_10_LC_4_21_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNICP62_10_LC_4_21_4  (
            .in0(_gnd_net_),
            .in1(N__39094),
            .in2(_gnd_net_),
            .in3(N__39361),
            .lcout(),
            .ltout(\pid_alt.m21_e_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIIO7C2_2_LC_4_21_5 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIIO7C2_2_LC_4_21_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIIO7C2_2_LC_4_21_5 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNIIO7C2_2_LC_4_21_5  (
            .in0(N__37280),
            .in1(N__37352),
            .in2(N__37131),
            .in3(N__37128),
            .lcout(),
            .ltout(\pid_alt.m21_e_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIO7B05_21_LC_4_21_6 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIO7B05_21_LC_4_21_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIO7B05_21_LC_4_21_6 .LUT_INIT=16'b1110101000101010;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNIO7B05_21_LC_4_21_6  (
            .in0(N__49474),
            .in1(N__37116),
            .in2(N__37110),
            .in3(N__39341),
            .lcout(),
            .ltout(\pid_alt.N_111_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.state_RNIAAPN5_1_LC_4_21_7 .C_ON=1'b0;
    defparam \pid_alt.state_RNIAAPN5_1_LC_4_21_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.state_RNIAAPN5_1_LC_4_21_7 .LUT_INIT=16'b1111111111000000;
    LogicCell40 \pid_alt.state_RNIAAPN5_1_LC_4_21_7  (
            .in0(_gnd_net_),
            .in1(N__65457),
            .in2(N__37107),
            .in3(N__66004),
            .lcout(\pid_alt.un1_reset_1_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIAP1A_13_LC_4_22_0 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIAP1A_13_LC_4_22_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIAP1A_13_LC_4_22_0 .LUT_INIT=16'b1011101110101010;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNIAP1A_13_LC_4_22_0  (
            .in0(N__49478),
            .in1(N__49438),
            .in2(_gnd_net_),
            .in3(N__49415),
            .lcout(\pid_alt.N_9_0 ),
            .ltout(\pid_alt.N_9_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI4SOH2_10_LC_4_22_1 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI4SOH2_10_LC_4_22_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI4SOH2_10_LC_4_22_1 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNI4SOH2_10_LC_4_22_1  (
            .in0(N__37404),
            .in1(N__37398),
            .in2(N__37389),
            .in3(N__39431),
            .lcout(\pid_alt.N_62_mux ),
            .ltout(\pid_alt.N_62_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_esr_1_LC_4_22_2 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_esr_1_LC_4_22_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_esr_1_LC_4_22_2 .LUT_INIT=16'b1100010010000000;
    LogicCell40 \pid_alt.error_i_acumm_esr_1_LC_4_22_2  (
            .in0(N__37241),
            .in1(N__37386),
            .in2(N__37371),
            .in3(N__37258),
            .lcout(\pid_alt.error_i_acummZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87265),
            .ce(N__49376),
            .sr(N__49341));
    defparam \pid_alt.error_i_acumm_esr_2_LC_4_22_3 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_esr_2_LC_4_22_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_esr_2_LC_4_22_3 .LUT_INIT=16'b1000100011000000;
    LogicCell40 \pid_alt.error_i_acumm_esr_2_LC_4_22_3  (
            .in0(N__48426),
            .in1(N__37356),
            .in2(N__37265),
            .in3(N__37242),
            .lcout(\pid_alt.error_i_acummZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87265),
            .ce(N__49376),
            .sr(N__49341));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIEPGB3_5_LC_4_22_4 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIEPGB3_5_LC_4_22_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIEPGB3_5_LC_4_22_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNIEPGB3_5_LC_4_22_4  (
            .in0(N__39432),
            .in1(N__48457),
            .in2(_gnd_net_),
            .in3(N__48424),
            .lcout(\pid_alt.N_159 ),
            .ltout(\pid_alt.N_159_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_esr_0_LC_4_22_5 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_esr_0_LC_4_22_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_esr_0_LC_4_22_5 .LUT_INIT=16'b1011100000000000;
    LogicCell40 \pid_alt.error_i_acumm_esr_0_LC_4_22_5  (
            .in0(N__48425),
            .in1(N__37240),
            .in2(N__37329),
            .in3(N__37326),
            .lcout(\pid_alt.error_i_acummZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87265),
            .ce(N__49376),
            .sr(N__49341));
    defparam \pid_alt.error_i_acumm_esr_4_LC_4_22_6 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_esr_4_LC_4_22_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_esr_4_LC_4_22_6 .LUT_INIT=16'b1111000111111101;
    LogicCell40 \pid_alt.error_i_acumm_esr_4_LC_4_22_6  (
            .in0(N__39433),
            .in1(N__48458),
            .in2(N__37248),
            .in3(N__48428),
            .lcout(\pid_alt.error_i_acummZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87265),
            .ce(N__49376),
            .sr(N__49341));
    defparam \pid_alt.error_i_acumm_esr_3_LC_4_22_7 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_esr_3_LC_4_22_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_esr_3_LC_4_22_7 .LUT_INIT=16'b1000100011000000;
    LogicCell40 \pid_alt.error_i_acumm_esr_3_LC_4_22_7  (
            .in0(N__48427),
            .in1(N__37281),
            .in2(N__37266),
            .in3(N__37243),
            .lcout(\pid_alt.error_i_acummZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87265),
            .ce(N__49376),
            .sr(N__49341));
    defparam \uart_drone_sync.aux_2__0__0_LC_5_5_2 .C_ON=1'b0;
    defparam \uart_drone_sync.aux_2__0__0_LC_5_5_2 .SEQ_MODE=4'b1000;
    defparam \uart_drone_sync.aux_2__0__0_LC_5_5_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone_sync.aux_2__0__0_LC_5_5_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37434),
            .lcout(\uart_drone_sync.aux_2__0__0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87045),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone_sync.aux_1__0__0_LC_5_5_3 .C_ON=1'b0;
    defparam \uart_drone_sync.aux_1__0__0_LC_5_5_3 .SEQ_MODE=4'b1000;
    defparam \uart_drone_sync.aux_1__0__0_LC_5_5_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone_sync.aux_1__0__0_LC_5_5_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41067),
            .lcout(\uart_drone_sync.aux_1__0__0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87045),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone_sync.aux_3__0__0_LC_5_6_0 .C_ON=1'b0;
    defparam \uart_drone_sync.aux_3__0__0_LC_5_6_0 .SEQ_MODE=4'b1000;
    defparam \uart_drone_sync.aux_3__0__0_LC_5_6_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone_sync.aux_3__0__0_LC_5_6_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37428),
            .lcout(\uart_drone_sync.aux_3__0__0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87053),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone_sync.Q_0__0_LC_5_6_1 .C_ON=1'b0;
    defparam \uart_drone_sync.Q_0__0_LC_5_6_1 .SEQ_MODE=4'b1000;
    defparam \uart_drone_sync.Q_0__0_LC_5_6_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone_sync.Q_0__0_LC_5_6_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37422),
            .lcout(debug_CH0_16A_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87053),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc_sync.Q_0__0_LC_5_6_6 .C_ON=1'b0;
    defparam \uart_pc_sync.Q_0__0_LC_5_6_6 .SEQ_MODE=4'b1000;
    defparam \uart_pc_sync.Q_0__0_LC_5_6_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_pc_sync.Q_0__0_LC_5_6_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39726),
            .lcout(debug_CH2_18A_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87053),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_2_LC_5_8_4 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_2_LC_5_8_4 .SEQ_MODE=4'b1000;
    defparam \uart_drone.timer_Count_2_LC_5_8_4 .LUT_INIT=16'b0000000010101000;
    LogicCell40 \uart_drone.timer_Count_2_LC_5_8_4  (
            .in0(N__37416),
            .in1(N__39811),
            .in2(N__39776),
            .in3(N__79995),
            .lcout(\uart_drone.timer_CountZ1Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87073),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_4_LC_5_8_6 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_4_LC_5_8_6 .SEQ_MODE=4'b1000;
    defparam \uart_drone.timer_Count_4_LC_5_8_6 .LUT_INIT=16'b0000000010101000;
    LogicCell40 \uart_drone.timer_Count_4_LC_5_8_6  (
            .in0(N__37782),
            .in1(N__39812),
            .in2(N__39777),
            .in3(N__79996),
            .lcout(\uart_drone.timer_CountZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87073),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_RNI5A9J_1_LC_5_9_0 .C_ON=1'b1;
    defparam \uart_drone.timer_Count_RNI5A9J_1_LC_5_9_0 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNI5A9J_1_LC_5_9_0 .LUT_INIT=16'b0001000100010001;
    LogicCell40 \uart_drone.timer_Count_RNI5A9J_1_LC_5_9_0  (
            .in0(N__39868),
            .in1(N__37508),
            .in2(N__39873),
            .in3(_gnd_net_),
            .lcout(\uart_drone.un1_state_2_0_a3_0 ),
            .ltout(),
            .carryin(bfn_5_9_0_),
            .carryout(\uart_drone.un4_timer_Count_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_RNO_0_2_LC_5_9_1 .C_ON=1'b1;
    defparam \uart_drone.timer_Count_RNO_0_2_LC_5_9_1 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNO_0_2_LC_5_9_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_drone.timer_Count_RNO_0_2_LC_5_9_1  (
            .in0(_gnd_net_),
            .in1(N__39835),
            .in2(_gnd_net_),
            .in3(N__37410),
            .lcout(\uart_drone.timer_Count_RNO_0_0_2 ),
            .ltout(),
            .carryin(\uart_drone.un4_timer_Count_1_cry_1 ),
            .carryout(\uart_drone.un4_timer_Count_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_RNO_0_3_LC_5_9_2 .C_ON=1'b1;
    defparam \uart_drone.timer_Count_RNO_0_3_LC_5_9_2 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNO_0_3_LC_5_9_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_drone.timer_Count_RNO_0_3_LC_5_9_2  (
            .in0(_gnd_net_),
            .in1(N__50832),
            .in2(_gnd_net_),
            .in3(N__37407),
            .lcout(\uart_drone.timer_Count_RNO_0_0_3 ),
            .ltout(),
            .carryin(\uart_drone.un4_timer_Count_1_cry_2 ),
            .carryout(\uart_drone.un4_timer_Count_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_RNO_0_4_LC_5_9_3 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_RNO_0_4_LC_5_9_3 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNO_0_4_LC_5_9_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uart_drone.timer_Count_RNO_0_4_LC_5_9_3  (
            .in0(_gnd_net_),
            .in1(N__50758),
            .in2(_gnd_net_),
            .in3(N__37785),
            .lcout(\uart_drone.timer_Count_RNO_0_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNIHKIA2_12_LC_5_9_4 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNIHKIA2_12_LC_5_9_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNIHKIA2_12_LC_5_9_4 .LUT_INIT=16'b1111010011111100;
    LogicCell40 \pid_alt.pid_prereg_esr_RNIHKIA2_12_LC_5_9_4  (
            .in0(N__37776),
            .in1(N__37719),
            .in2(N__37647),
            .in3(N__37547),
            .lcout(\pid_alt.source_pid_9_0_tz_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_RNO_0_1_LC_5_9_5 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_RNO_0_1_LC_5_9_5 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNO_0_1_LC_5_9_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_drone.timer_Count_RNO_0_1_LC_5_9_5  (
            .in0(N__37509),
            .in1(N__39872),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\uart_drone.timer_Count_RNO_0_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_1_LC_5_9_6 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_1_LC_5_9_6 .SEQ_MODE=4'b1000;
    defparam \uart_drone.timer_Count_1_LC_5_9_6 .LUT_INIT=16'b0000000011100000;
    LogicCell40 \uart_drone.timer_Count_1_LC_5_9_6  (
            .in0(N__39767),
            .in1(N__39816),
            .in2(N__37512),
            .in3(N__79997),
            .lcout(\uart_drone.timer_CountZ1Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87085),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.source_pid_1_10_LC_5_10_0 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_10_LC_5_10_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_10_LC_5_10_0 .LUT_INIT=16'b1101110111110000;
    LogicCell40 \pid_alt.source_pid_1_10_LC_5_10_0  (
            .in0(N__37834),
            .in1(N__37500),
            .in2(N__44656),
            .in3(N__65407),
            .lcout(throttle_order_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87101),
            .ce(),
            .sr(N__37814));
    defparam \pid_alt.pid_prereg_esr_RNIIM6H1_0_6_LC_5_10_1 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNIIM6H1_0_6_LC_5_10_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNIIM6H1_0_6_LC_5_10_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_alt.pid_prereg_esr_RNIIM6H1_0_6_LC_5_10_1  (
            .in0(N__37907),
            .in1(N__37937),
            .in2(N__37878),
            .in3(N__37967),
            .lcout(),
            .ltout(\pid_alt.source_pid_1_sqmuxa_0_a2_1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNI4GSA2_10_LC_5_10_2 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNI4GSA2_10_LC_5_10_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNI4GSA2_10_LC_5_10_2 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \pid_alt.pid_prereg_esr_RNI4GSA2_10_LC_5_10_2  (
            .in0(N__37456),
            .in1(N__37499),
            .in2(N__37470),
            .in3(N__65400),
            .lcout(\pid_alt.source_pid_1_sqmuxa_0_a2_1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.source_pid_1_11_LC_5_10_3 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_11_LC_5_10_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_11_LC_5_10_3 .LUT_INIT=16'b1111101001110010;
    LogicCell40 \pid_alt.source_pid_1_11_LC_5_10_3  (
            .in0(N__65401),
            .in1(N__37835),
            .in2(N__41500),
            .in3(N__37457),
            .lcout(throttle_order_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87101),
            .ce(),
            .sr(N__37814));
    defparam \pid_alt.source_pid_1_6_LC_5_10_4 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_6_LC_5_10_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_6_LC_5_10_4 .LUT_INIT=16'b1010111111001100;
    LogicCell40 \pid_alt.source_pid_1_6_LC_5_10_4  (
            .in0(N__37968),
            .in1(N__41431),
            .in2(N__37842),
            .in3(N__65408),
            .lcout(throttle_order_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87101),
            .ce(),
            .sr(N__37814));
    defparam \pid_alt.source_pid_1_7_LC_5_10_5 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_7_LC_5_10_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_7_LC_5_10_5 .LUT_INIT=16'b1111101001110010;
    LogicCell40 \pid_alt.source_pid_1_7_LC_5_10_5  (
            .in0(N__65402),
            .in1(N__37839),
            .in2(N__47188),
            .in3(N__37938),
            .lcout(throttle_order_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87101),
            .ce(),
            .sr(N__37814));
    defparam \pid_alt.source_pid_1_8_LC_5_10_6 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_8_LC_5_10_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_8_LC_5_10_6 .LUT_INIT=16'b1111110001110100;
    LogicCell40 \pid_alt.source_pid_1_8_LC_5_10_6  (
            .in0(N__37840),
            .in1(N__65403),
            .in2(N__41408),
            .in3(N__37908),
            .lcout(throttle_order_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87101),
            .ce(),
            .sr(N__37814));
    defparam \pid_alt.source_pid_1_9_LC_5_10_7 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_9_LC_5_10_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_9_LC_5_10_7 .LUT_INIT=16'b1010110011111100;
    LogicCell40 \pid_alt.source_pid_1_9_LC_5_10_7  (
            .in0(N__37877),
            .in1(N__41224),
            .in2(N__65432),
            .in3(N__37841),
            .lcout(throttle_order_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87101),
            .ce(),
            .sr(N__37814));
    defparam \scaler_4.source_data_1_esr_5_LC_5_11_0 .C_ON=1'b0;
    defparam \scaler_4.source_data_1_esr_5_LC_5_11_0 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_5_LC_5_11_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \scaler_4.source_data_1_esr_5_LC_5_11_0  (
            .in0(N__42726),
            .in1(N__42674),
            .in2(_gnd_net_),
            .in3(N__42753),
            .lcout(scaler_4_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87116),
            .ce(N__42425),
            .sr(N__79581));
    defparam \uart_pc.data_Aux_RNO_0_0_LC_5_11_1 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_RNO_0_0_LC_5_11_1 .SEQ_MODE=4'b0000;
    defparam \uart_pc.data_Aux_RNO_0_0_LC_5_11_1 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \uart_pc.data_Aux_RNO_0_0_LC_5_11_1  (
            .in0(N__39948),
            .in1(N__39993),
            .in2(_gnd_net_),
            .in3(N__41583),
            .lcout(\uart_pc.data_Auxce_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_Aux_RNO_0_1_LC_5_11_2 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_RNO_0_1_LC_5_11_2 .SEQ_MODE=4'b0000;
    defparam \uart_pc.data_Aux_RNO_0_1_LC_5_11_2 .LUT_INIT=16'b0000000000001010;
    LogicCell40 \uart_pc.data_Aux_RNO_0_1_LC_5_11_2  (
            .in0(N__41584),
            .in1(_gnd_net_),
            .in2(N__40006),
            .in3(N__39949),
            .lcout(\uart_pc.data_Auxce_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_Aux_RNO_0_2_LC_5_11_3 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_RNO_0_2_LC_5_11_3 .SEQ_MODE=4'b0000;
    defparam \uart_pc.data_Aux_RNO_0_2_LC_5_11_3 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \uart_pc.data_Aux_RNO_0_2_LC_5_11_3  (
            .in0(N__39950),
            .in1(N__39997),
            .in2(_gnd_net_),
            .in3(N__41585),
            .lcout(\uart_pc.data_Auxce_0_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_Aux_RNO_0_3_LC_5_11_4 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_RNO_0_3_LC_5_11_4 .SEQ_MODE=4'b0000;
    defparam \uart_pc.data_Aux_RNO_0_3_LC_5_11_4 .LUT_INIT=16'b0000000010100000;
    LogicCell40 \uart_pc.data_Aux_RNO_0_3_LC_5_11_4  (
            .in0(N__41586),
            .in1(_gnd_net_),
            .in2(N__40007),
            .in3(N__39951),
            .lcout(\uart_pc.data_Auxce_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_Aux_RNO_0_4_LC_5_11_5 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_RNO_0_4_LC_5_11_5 .SEQ_MODE=4'b0000;
    defparam \uart_pc.data_Aux_RNO_0_4_LC_5_11_5 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \uart_pc.data_Aux_RNO_0_4_LC_5_11_5  (
            .in0(N__39952),
            .in1(N__40001),
            .in2(_gnd_net_),
            .in3(N__41587),
            .lcout(\uart_pc.data_Auxce_0_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_Aux_RNO_0_5_LC_5_11_6 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_RNO_0_5_LC_5_11_6 .SEQ_MODE=4'b0000;
    defparam \uart_pc.data_Aux_RNO_0_5_LC_5_11_6 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \uart_pc.data_Aux_RNO_0_5_LC_5_11_6  (
            .in0(N__41588),
            .in1(_gnd_net_),
            .in2(N__40008),
            .in3(N__39953),
            .lcout(\uart_pc.data_Auxce_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_Aux_RNO_0_6_LC_5_11_7 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_RNO_0_6_LC_5_11_7 .SEQ_MODE=4'b0000;
    defparam \uart_pc.data_Aux_RNO_0_6_LC_5_11_7 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \uart_pc.data_Aux_RNO_0_6_LC_5_11_7  (
            .in0(N__39954),
            .in1(N__40005),
            .in2(_gnd_net_),
            .in3(N__41589),
            .lcout(\uart_pc.data_Auxce_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_Aux_0_LC_5_12_0 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_0_LC_5_12_0 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_Aux_0_LC_5_12_0 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \uart_pc.data_Aux_0_LC_5_12_0  (
            .in0(N__38133),
            .in1(N__40212),
            .in2(N__38126),
            .in3(N__40490),
            .lcout(\uart_pc.data_AuxZ1Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87132),
            .ce(),
            .sr(N__39912));
    defparam \uart_pc.data_Aux_1_LC_5_12_1 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_1_LC_5_12_1 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_Aux_1_LC_5_12_1 .LUT_INIT=16'b1100110011100100;
    LogicCell40 \uart_pc.data_Aux_1_LC_5_12_1  (
            .in0(N__38109),
            .in1(N__38102),
            .in2(N__40239),
            .in3(N__40493),
            .lcout(\uart_pc.data_AuxZ1Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87132),
            .ce(),
            .sr(N__39912));
    defparam \uart_pc.data_Aux_2_LC_5_12_2 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_2_LC_5_12_2 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_Aux_2_LC_5_12_2 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \uart_pc.data_Aux_2_LC_5_12_2  (
            .in0(N__38085),
            .in1(N__40213),
            .in2(N__38079),
            .in3(N__40491),
            .lcout(\uart_pc.data_AuxZ1Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87132),
            .ce(),
            .sr(N__39912));
    defparam \uart_pc.data_Aux_3_LC_5_12_3 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_3_LC_5_12_3 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_Aux_3_LC_5_12_3 .LUT_INIT=16'b1101100011001100;
    LogicCell40 \uart_pc.data_Aux_3_LC_5_12_3  (
            .in0(N__40487),
            .in1(N__38054),
            .in2(N__40240),
            .in3(N__38064),
            .lcout(\uart_pc.data_AuxZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87132),
            .ce(),
            .sr(N__39912));
    defparam \uart_pc.data_Aux_4_LC_5_12_4 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_4_LC_5_12_4 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_Aux_4_LC_5_12_4 .LUT_INIT=16'b1111110100001000;
    LogicCell40 \uart_pc.data_Aux_4_LC_5_12_4  (
            .in0(N__38043),
            .in1(N__40214),
            .in2(N__40497),
            .in3(N__38030),
            .lcout(\uart_pc.data_AuxZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87132),
            .ce(),
            .sr(N__39912));
    defparam \uart_pc.data_Aux_5_LC_5_12_5 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_5_LC_5_12_5 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_Aux_5_LC_5_12_5 .LUT_INIT=16'b1101100011001100;
    LogicCell40 \uart_pc.data_Aux_5_LC_5_12_5  (
            .in0(N__40488),
            .in1(N__38006),
            .in2(N__40241),
            .in3(N__38016),
            .lcout(\uart_pc.data_AuxZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87132),
            .ce(),
            .sr(N__39912));
    defparam \uart_pc.data_Aux_6_LC_5_12_6 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_6_LC_5_12_6 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_Aux_6_LC_5_12_6 .LUT_INIT=16'b1010101011001010;
    LogicCell40 \uart_pc.data_Aux_6_LC_5_12_6  (
            .in0(N__37979),
            .in1(N__40215),
            .in2(N__37995),
            .in3(N__40492),
            .lcout(\uart_pc.data_AuxZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87132),
            .ce(),
            .sr(N__39912));
    defparam \uart_pc.data_Aux_7_LC_5_12_7 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_7_LC_5_12_7 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_Aux_7_LC_5_12_7 .LUT_INIT=16'b1101100011001100;
    LogicCell40 \uart_pc.data_Aux_7_LC_5_12_7  (
            .in0(N__40489),
            .in1(N__38255),
            .in2(N__40242),
            .in3(N__41715),
            .lcout(\uart_pc.data_AuxZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87132),
            .ce(),
            .sr(N__39912));
    defparam \uart_pc.timer_Count_RNIPD2K1_2_LC_5_13_0 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_RNIPD2K1_2_LC_5_13_0 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNIPD2K1_2_LC_5_13_0 .LUT_INIT=16'b1100110010000000;
    LogicCell40 \uart_pc.timer_Count_RNIPD2K1_2_LC_5_13_0  (
            .in0(N__40440),
            .in1(N__40521),
            .in2(N__40323),
            .in3(N__40383),
            .lcout(\uart_pc.data_rdyc_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_RNO_0_3_LC_5_13_3 .C_ON=1'b0;
    defparam \uart_pc.state_RNO_0_3_LC_5_13_3 .SEQ_MODE=4'b0000;
    defparam \uart_pc.state_RNO_0_3_LC_5_13_3 .LUT_INIT=16'b0000000001111111;
    LogicCell40 \uart_pc.state_RNO_0_3_LC_5_13_3  (
            .in0(N__40385),
            .in1(N__40442),
            .in2(N__40119),
            .in3(N__41627),
            .lcout(),
            .ltout(\uart_pc.N_145_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_3_LC_5_13_4 .C_ON=1'b0;
    defparam \uart_pc.state_3_LC_5_13_4 .SEQ_MODE=4'b1000;
    defparam \uart_pc.state_3_LC_5_13_4 .LUT_INIT=16'b0000000000001011;
    LogicCell40 \uart_pc.state_3_LC_5_13_4  (
            .in0(N__40118),
            .in1(N__38241),
            .in2(N__38244),
            .in3(N__79992),
            .lcout(\uart_pc.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87150),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNI5UFA2_3_LC_5_13_5 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_RNI5UFA2_3_LC_5_13_5 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNI5UFA2_3_LC_5_13_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uart_pc.timer_Count_RNI5UFA2_3_LC_5_13_5  (
            .in0(N__40384),
            .in1(N__40441),
            .in2(_gnd_net_),
            .in3(N__41714),
            .lcout(\uart_pc.N_144_1 ),
            .ltout(\uart_pc.N_144_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_4_LC_5_13_6 .C_ON=1'b0;
    defparam \uart_pc.state_4_LC_5_13_6 .SEQ_MODE=4'b1000;
    defparam \uart_pc.state_4_LC_5_13_6 .LUT_INIT=16'b1100110011101100;
    LogicCell40 \uart_pc.state_4_LC_5_13_6  (
            .in0(N__41628),
            .in1(N__41951),
            .in2(N__38235),
            .in3(N__79993),
            .lcout(\uart_pc.stateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87150),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNIVGCQ_12_LC_5_13_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIVGCQ_12_LC_5_13_7 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIVGCQ_12_LC_5_13_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Commands_frame_decoder.state_RNIVGCQ_12_LC_5_13_7  (
            .in0(_gnd_net_),
            .in1(N__38232),
            .in2(_gnd_net_),
            .in3(N__38368),
            .lcout(\Commands_frame_decoder.source_xy_ki_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kp_4_LC_5_14_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kp_4_LC_5_14_0 .SEQ_MODE=4'b1001;
    defparam \Commands_frame_decoder.source_alt_kp_4_LC_5_14_0 .LUT_INIT=16'b1110101000101010;
    LogicCell40 \Commands_frame_decoder.source_alt_kp_4_LC_5_14_0  (
            .in0(N__38174),
            .in1(N__38367),
            .in2(N__38217),
            .in3(N__85019),
            .lcout(alt_kp_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87166),
            .ce(),
            .sr(N__79599));
    defparam \uart_pc.data_rdy_LC_5_14_1 .C_ON=1'b0;
    defparam \uart_pc.data_rdy_LC_5_14_1 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_rdy_LC_5_14_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uart_pc.data_rdy_LC_5_14_1  (
            .in0(_gnd_net_),
            .in1(N__38153),
            .in2(_gnd_net_),
            .in3(N__40238),
            .lcout(uart_pc_data_rdy),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87166),
            .ce(),
            .sr(N__79599));
    defparam \Commands_frame_decoder.state_RNIEI1J_2_LC_5_14_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIEI1J_2_LC_5_14_2 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIEI1J_2_LC_5_14_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Commands_frame_decoder.state_RNIEI1J_2_LC_5_14_2  (
            .in0(_gnd_net_),
            .in1(N__38535),
            .in2(_gnd_net_),
            .in3(N__38366),
            .lcout(\Commands_frame_decoder.un1_sink_data_valid_2_0 ),
            .ltout(\Commands_frame_decoder.un1_sink_data_valid_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNIBV7S_2_LC_5_14_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIBV7S_2_LC_5_14_3 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIBV7S_2_LC_5_14_3 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \Commands_frame_decoder.state_RNIBV7S_2_LC_5_14_3  (
            .in0(N__79929),
            .in1(_gnd_net_),
            .in2(N__38514),
            .in3(_gnd_net_),
            .lcout(\Commands_frame_decoder.un1_sink_data_valid_2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNIC08S_3_LC_5_14_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIC08S_3_LC_5_14_4 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIC08S_3_LC_5_14_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \Commands_frame_decoder.state_RNIC08S_3_LC_5_14_4  (
            .in0(_gnd_net_),
            .in1(N__79928),
            .in2(_gnd_net_),
            .in3(N__38322),
            .lcout(\Commands_frame_decoder.source_CH2data_1_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_3_LC_5_14_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_3_LC_5_14_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_3_LC_5_14_5 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \Commands_frame_decoder.state_3_LC_5_14_5  (
            .in0(N__38478),
            .in1(N__38491),
            .in2(_gnd_net_),
            .in3(N__39307),
            .lcout(\Commands_frame_decoder.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87166),
            .ce(),
            .sr(N__79599));
    defparam \Commands_frame_decoder.state_RNIFJ1J_3_LC_5_14_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIFJ1J_3_LC_5_14_6 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIFJ1J_3_LC_5_14_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Commands_frame_decoder.state_RNIFJ1J_3_LC_5_14_6  (
            .in0(_gnd_net_),
            .in1(N__38477),
            .in2(_gnd_net_),
            .in3(N__38365),
            .lcout(\Commands_frame_decoder.source_CH2data_1_sqmuxa ),
            .ltout(\Commands_frame_decoder.source_CH2data_1_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_4_LC_5_14_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_4_LC_5_14_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_4_LC_5_14_7 .LUT_INIT=16'b1111110011110000;
    LogicCell40 \Commands_frame_decoder.state_4_LC_5_14_7  (
            .in0(_gnd_net_),
            .in1(N__38309),
            .in2(N__38316),
            .in3(N__39308),
            .lcout(\Commands_frame_decoder.stateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87166),
            .ce(),
            .sr(N__79599));
    defparam \pid_front.error_p_reg_esr_17_LC_5_15_0 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_17_LC_5_15_0 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_17_LC_5_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_p_reg_esr_17_LC_5_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38295),
            .lcout(\pid_front.error_p_regZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87180),
            .ce(N__86288),
            .sr(N__86031));
    defparam \pid_front.error_p_reg_esr_3_LC_5_15_1 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_3_LC_5_15_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_3_LC_5_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_p_reg_esr_3_LC_5_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38280),
            .lcout(\pid_front.error_p_regZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87180),
            .ce(N__86288),
            .sr(N__86031));
    defparam \pid_front.error_p_reg_esr_9_LC_5_15_2 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_9_LC_5_15_2 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_9_LC_5_15_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_p_reg_esr_9_LC_5_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38271),
            .lcout(\pid_front.error_p_regZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87180),
            .ce(N__86288),
            .sr(N__86031));
    defparam \pid_alt.error_d_reg_prev_esr_RNI64JA4_12_LC_5_16_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI64JA4_12_LC_5_16_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI64JA4_12_LC_5_16_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI64JA4_12_LC_5_16_0  (
            .in0(N__38828),
            .in1(N__38835),
            .in2(N__38681),
            .in3(N__38690),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI64JA4Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIJGHM_12_LC_5_16_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIJGHM_12_LC_5_16_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIJGHM_12_LC_5_16_1 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIJGHM_12_LC_5_16_1  (
            .in0(N__38651),
            .in1(N__38660),
            .in2(_gnd_net_),
            .in3(N__38632),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIJGHMZ0Z_12 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNIJGHMZ0Z_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNISAO32_12_LC_5_16_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNISAO32_12_LC_5_16_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNISAO32_12_LC_5_16_2 .LUT_INIT=16'b1111101010100000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNISAO32_12_LC_5_16_2  (
            .in0(N__38829),
            .in1(_gnd_net_),
            .in2(N__38805),
            .in3(N__38691),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNISAO32Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIMJHM_0_13_LC_5_16_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIMJHM_0_13_LC_5_16_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIMJHM_0_13_LC_5_16_3 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIMJHM_0_13_LC_5_16_3  (
            .in0(N__38783),
            .in1(N__38759),
            .in2(_gnd_net_),
            .in3(N__38719),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIMJHM_0Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_12_LC_5_16_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_12_LC_5_16_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_12_LC_5_16_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_12_LC_5_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38634),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87194),
            .ce(N__51483),
            .sr(N__79609));
    defparam \pid_alt.error_d_reg_prev_esr_RNIAPQ62_11_LC_5_16_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIAPQ62_11_LC_5_16_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIAPQ62_11_LC_5_16_5 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIAPQ62_11_LC_5_16_5  (
            .in0(N__38613),
            .in1(N__38586),
            .in2(_gnd_net_),
            .in3(N__38570),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIAPQ62Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIJGHM_0_12_LC_5_16_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIJGHM_0_12_LC_5_16_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIJGHM_0_12_LC_5_16_6 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIJGHM_0_12_LC_5_16_6  (
            .in0(N__38661),
            .in1(N__38652),
            .in2(_gnd_net_),
            .in3(N__38633),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIJGHM_0Z0Z_12 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNIJGHM_0Z0Z_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIB8KD4_11_LC_5_16_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIB8KD4_11_LC_5_16_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIB8KD4_11_LC_5_16_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIB8KD4_11_LC_5_16_7  (
            .in0(N__38607),
            .in1(N__38585),
            .in2(N__38574),
            .in3(N__38569),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIB8KD4Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_0_LC_5_17_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_0_LC_5_17_0 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_0_LC_5_17_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_0_LC_5_17_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59332),
            .lcout(drone_altitude_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87211),
            .ce(N__54129),
            .sr(N__79616));
    defparam \dron_frame_decoder_1.source_Altitude_esr_1_LC_5_17_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_1_LC_5_17_1 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_1_LC_5_17_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_1_LC_5_17_1  (
            .in0(N__59204),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(drone_altitude_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87211),
            .ce(N__54129),
            .sr(N__79616));
    defparam \dron_frame_decoder_1.source_Altitude_esr_4_LC_5_17_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_4_LC_5_17_2 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_4_LC_5_17_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_4_LC_5_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58935),
            .lcout(\dron_frame_decoder_1.drone_altitude_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87211),
            .ce(N__54129),
            .sr(N__79616));
    defparam \dron_frame_decoder_1.source_Altitude_esr_5_LC_5_17_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_5_LC_5_17_3 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_5_LC_5_17_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_5_LC_5_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58834),
            .lcout(\dron_frame_decoder_1.drone_altitude_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87211),
            .ce(N__54129),
            .sr(N__79616));
    defparam \dron_frame_decoder_1.source_Altitude_esr_6_LC_5_17_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_6_LC_5_17_4 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_6_LC_5_17_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_6_LC_5_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58758),
            .lcout(\dron_frame_decoder_1.drone_altitude_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87211),
            .ce(N__54129),
            .sr(N__79616));
    defparam \dron_frame_decoder_1.source_Altitude_esr_7_LC_5_17_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_7_LC_5_17_5 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_7_LC_5_17_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_7_LC_5_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58658),
            .lcout(\dron_frame_decoder_1.drone_altitude_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87211),
            .ce(N__54129),
            .sr(N__79616));
    defparam \scaler_4.un3_source_data_un3_source_data_0_axb_7_LC_5_18_0 .C_ON=1'b0;
    defparam \scaler_4.un3_source_data_un3_source_data_0_axb_7_LC_5_18_0 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_axb_7_LC_5_18_0 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_axb_7_LC_5_18_0  (
            .in0(_gnd_net_),
            .in1(N__53897),
            .in2(_gnd_net_),
            .in3(N__53930),
            .lcout(\scaler_4.un3_source_data_0_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_CH4data_ess_7_LC_5_18_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH4data_ess_7_LC_5_18_1 .SEQ_MODE=4'b1001;
    defparam \Commands_frame_decoder.source_CH4data_ess_7_LC_5_18_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH4data_ess_7_LC_5_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85362),
            .lcout(frame_decoder_CH4data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87226),
            .ce(N__41531),
            .sr(N__79623));
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIHIDC_4_LC_5_18_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIHIDC_4_LC_5_18_2 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIHIDC_4_LC_5_18_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_RNIHIDC_4_LC_5_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38868),
            .lcout(drone_altitude_i_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIIJDC_5_LC_5_18_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIIJDC_5_LC_5_18_3 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIIJDC_5_LC_5_18_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_RNIIJDC_5_LC_5_18_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38856),
            .lcout(drone_altitude_i_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIJKDC_6_LC_5_18_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIJKDC_6_LC_5_18_4 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIJKDC_6_LC_5_18_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_RNIJKDC_6_LC_5_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39030),
            .lcout(drone_altitude_i_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIKLDC_7_LC_5_18_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIKLDC_7_LC_5_18_5 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIKLDC_7_LC_5_18_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_RNIKLDC_7_LC_5_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39018),
            .lcout(drone_altitude_i_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNILMDC_8_LC_5_18_6 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNILMDC_8_LC_5_18_6 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNILMDC_8_LC_5_18_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_RNILMDC_8_LC_5_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40656),
            .lcout(drone_altitude_i_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIMNDC_9_LC_5_18_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIMNDC_9_LC_5_18_7 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIMNDC_9_LC_5_18_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_RNIMNDC_9_LC_5_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40644),
            .lcout(drone_altitude_i_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kp_e_0_0_LC_5_19_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_0_LC_5_19_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_0_LC_5_19_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_kp_e_0_0_LC_5_19_0  (
            .in0(_gnd_net_),
            .in1(N__83787),
            .in2(_gnd_net_),
            .in3(N__86167),
            .lcout(alt_kp_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87240),
            .ce(N__39165),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kp_e_0_1_LC_5_19_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_1_LC_5_19_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_1_LC_5_19_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Commands_frame_decoder.source_alt_kp_e_0_1_LC_5_19_1  (
            .in0(N__86168),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84160),
            .lcout(alt_kp_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87240),
            .ce(N__39165),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kp_e_0_2_LC_5_19_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_2_LC_5_19_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_2_LC_5_19_2 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \Commands_frame_decoder.source_alt_kp_e_0_2_LC_5_19_2  (
            .in0(N__77570),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__86169),
            .lcout(alt_kp_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87240),
            .ce(N__39165),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kp_e_0_3_LC_5_19_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_3_LC_5_19_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_3_LC_5_19_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Commands_frame_decoder.source_alt_kp_e_0_3_LC_5_19_3  (
            .in0(N__86170),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__83984),
            .lcout(alt_kp_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87240),
            .ce(N__39165),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kp_0_e_0_4_LC_5_19_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kp_0_e_0_4_LC_5_19_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kp_0_e_0_4_LC_5_19_4 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \Commands_frame_decoder.source_alt_kp_0_e_0_4_LC_5_19_4  (
            .in0(N__85188),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__86166),
            .lcout(alt_kp_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87240),
            .ce(N__39165),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kp_e_0_5_LC_5_19_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_5_LC_5_19_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_5_LC_5_19_5 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Commands_frame_decoder.source_alt_kp_e_0_5_LC_5_19_5  (
            .in0(N__86171),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73627),
            .lcout(alt_kp_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87240),
            .ce(N__39165),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kp_e_0_6_LC_5_19_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_6_LC_5_19_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_6_LC_5_19_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_kp_e_0_6_LC_5_19_6  (
            .in0(_gnd_net_),
            .in1(N__85361),
            .in2(_gnd_net_),
            .in3(N__86172),
            .lcout(alt_kp_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87240),
            .ce(N__39165),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIUHR9_10_LC_5_19_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIUHR9_10_LC_5_19_7 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIUHR9_10_LC_5_19_7 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_RNIUHR9_10_LC_5_19_7  (
            .in0(_gnd_net_),
            .in1(N__40692),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(drone_altitude_i_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_CH1data_esr_4_LC_5_20_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH1data_esr_4_LC_5_20_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH1data_esr_4_LC_5_20_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH1data_esr_4_LC_5_20_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85039),
            .lcout(alt_command_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87251),
            .ce(N__39105),
            .sr(N__79639));
    defparam \Commands_frame_decoder.source_CH1data_esr_5_LC_5_20_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH1data_esr_5_LC_5_20_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH1data_esr_5_LC_5_20_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Commands_frame_decoder.source_CH1data_esr_5_LC_5_20_1  (
            .in0(N__85187),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(alt_command_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87251),
            .ce(N__39105),
            .sr(N__79639));
    defparam \Commands_frame_decoder.source_CH1data_esr_6_LC_5_20_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH1data_esr_6_LC_5_20_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH1data_esr_6_LC_5_20_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH1data_esr_6_LC_5_20_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73626),
            .lcout(alt_command_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87251),
            .ce(N__39105),
            .sr(N__79639));
    defparam \Commands_frame_decoder.source_CH1data_esr_7_LC_5_20_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH1data_esr_7_LC_5_20_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH1data_esr_7_LC_5_20_3 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \Commands_frame_decoder.source_CH1data_esr_7_LC_5_20_3  (
            .in0(_gnd_net_),
            .in1(N__85363),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(alt_command_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87251),
            .ce(N__39105),
            .sr(N__79639));
    defparam \pid_alt.error_i_acumm_10_LC_5_21_0 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_10_LC_5_21_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_10_LC_5_21_0 .LUT_INIT=16'b1010111111001100;
    LogicCell40 \pid_alt.error_i_acumm_10_LC_5_21_0  (
            .in0(N__39096),
            .in1(N__39074),
            .in2(N__39458),
            .in3(N__65449),
            .lcout(\pid_alt.error_i_acummZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87257),
            .ce(),
            .sr(N__49351));
    defparam \pid_alt.error_i_acumm_11_LC_5_21_1 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_11_LC_5_21_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_11_LC_5_21_1 .LUT_INIT=16'b1101111111010000;
    LogicCell40 \pid_alt.error_i_acumm_11_LC_5_21_1  (
            .in0(N__39448),
            .in1(N__39060),
            .in2(N__65454),
            .in3(N__39620),
            .lcout(\pid_alt.error_i_acummZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87257),
            .ce(),
            .sr(N__49351));
    defparam \pid_alt.error_i_acumm_6_LC_5_21_2 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_6_LC_5_21_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_6_LC_5_21_2 .LUT_INIT=16'b1100111110101010;
    LogicCell40 \pid_alt.error_i_acumm_6_LC_5_21_2  (
            .in0(N__39572),
            .in1(N__39606),
            .in2(N__39459),
            .in3(N__65450),
            .lcout(\pid_alt.error_i_acummZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87257),
            .ce(),
            .sr(N__49351));
    defparam \pid_alt.error_i_acumm_7_LC_5_21_3 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_7_LC_5_21_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_7_LC_5_21_3 .LUT_INIT=16'b1101111111010000;
    LogicCell40 \pid_alt.error_i_acumm_7_LC_5_21_3  (
            .in0(N__39449),
            .in1(N__39558),
            .in2(N__65455),
            .in3(N__39518),
            .lcout(\pid_alt.error_i_acummZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87257),
            .ce(),
            .sr(N__49351));
    defparam \pid_alt.error_i_acumm_8_LC_5_21_4 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_8_LC_5_21_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_8_LC_5_21_4 .LUT_INIT=16'b1011100011111100;
    LogicCell40 \pid_alt.error_i_acumm_8_LC_5_21_4  (
            .in0(N__39500),
            .in1(N__65439),
            .in2(N__39479),
            .in3(N__39451),
            .lcout(\pid_alt.error_i_acummZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87257),
            .ce(),
            .sr(N__49351));
    defparam \pid_alt.error_i_acumm_9_LC_5_21_5 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_9_LC_5_21_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_9_LC_5_21_5 .LUT_INIT=16'b1111110001011100;
    LogicCell40 \pid_alt.error_i_acumm_9_LC_5_21_5  (
            .in0(N__39450),
            .in1(N__39386),
            .in2(N__65456),
            .in3(N__39411),
            .lcout(\pid_alt.error_i_acummZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87257),
            .ce(),
            .sr(N__49351));
    defparam \pid_alt.state_RNIVV066_1_LC_5_21_6 .C_ON=1'b0;
    defparam \pid_alt.state_RNIVV066_1_LC_5_21_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.state_RNIVV066_1_LC_5_21_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \pid_alt.state_RNIVV066_1_LC_5_21_6  (
            .in0(_gnd_net_),
            .in1(N__65437),
            .in2(_gnd_net_),
            .in3(N__49328),
            .lcout(\pid_alt.N_72_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_12_LC_5_21_7 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_12_LC_5_21_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_12_LC_5_21_7 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \pid_alt.error_i_acumm_12_LC_5_21_7  (
            .in0(N__65438),
            .in1(N__39368),
            .in2(N__39329),
            .in3(N__39342),
            .lcout(\pid_alt.error_i_acummZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87257),
            .ce(),
            .sr(N__49351));
    defparam \Commands_frame_decoder.state_10_LC_5_22_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_10_LC_5_22_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_10_LC_5_22_1 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \Commands_frame_decoder.state_10_LC_5_22_1  (
            .in0(N__39220),
            .in1(N__40293),
            .in2(_gnd_net_),
            .in3(N__39309),
            .lcout(\Commands_frame_decoder.stateZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87261),
            .ce(),
            .sr(N__79655));
    defparam \reset_module_System.count_RNI9O1P_2_LC_7_1_0 .C_ON=1'b0;
    defparam \reset_module_System.count_RNI9O1P_2_LC_7_1_0 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNI9O1P_2_LC_7_1_0 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \reset_module_System.count_RNI9O1P_2_LC_7_1_0  (
            .in0(N__40754),
            .in1(N__40799),
            .in2(N__40824),
            .in3(N__41184),
            .lcout(\reset_module_System.reset6_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNI97FD_5_LC_7_1_2 .C_ON=1'b0;
    defparam \reset_module_System.count_RNI97FD_5_LC_7_1_2 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNI97FD_5_LC_7_1_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \reset_module_System.count_RNI97FD_5_LC_7_1_2  (
            .in0(N__40724),
            .in1(N__40739),
            .in2(N__40710),
            .in3(N__40769),
            .lcout(\reset_module_System.reset6_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_2_LC_7_1_5 .C_ON=1'b0;
    defparam \reset_module_System.count_2_LC_7_1_5 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_2_LC_7_1_5 .LUT_INIT=16'b0100110011001100;
    LogicCell40 \reset_module_System.count_2_LC_7_1_5  (
            .in0(N__40973),
            .in1(N__40809),
            .in2(N__41031),
            .in3(N__40997),
            .lcout(\reset_module_System.countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__86997),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.reset_LC_7_1_7 .C_ON=1'b0;
    defparam \reset_module_System.reset_LC_7_1_7 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.reset_LC_7_1_7 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \reset_module_System.reset_LC_7_1_7  (
            .in0(N__41026),
            .in1(N__40971),
            .in2(_gnd_net_),
            .in3(N__40996),
            .lcout(reset_system),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__86997),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNI10J41_1_LC_7_2_1 .C_ON=1'b0;
    defparam \reset_module_System.count_RNI10J41_1_LC_7_2_1 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNI10J41_1_LC_7_2_1 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \reset_module_System.count_RNI10J41_1_LC_7_2_1  (
            .in0(N__40878),
            .in1(N__40785),
            .in2(N__40842),
            .in3(N__40949),
            .lcout(\reset_module_System.reset6_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNI53692_14_LC_7_2_5 .C_ON=1'b0;
    defparam \reset_module_System.count_RNI53692_14_LC_7_2_5 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNI53692_14_LC_7_2_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \reset_module_System.count_RNI53692_14_LC_7_2_5  (
            .in0(N__40895),
            .in1(N__39675),
            .in2(N__40860),
            .in3(N__41139),
            .lcout(),
            .ltout(\reset_module_System.reset6_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNIN3HK3_12_LC_7_2_6 .C_ON=1'b0;
    defparam \reset_module_System.count_RNIN3HK3_12_LC_7_2_6 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNIN3HK3_12_LC_7_2_6 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \reset_module_System.count_RNIN3HK3_12_LC_7_2_6  (
            .in0(N__40917),
            .in1(N__41050),
            .in2(N__39669),
            .in3(N__39666),
            .lcout(\reset_module_System.reset6_19 ),
            .ltout(\reset_module_System.reset6_19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_0_LC_7_2_7 .C_ON=1'b0;
    defparam \reset_module_System.count_0_LC_7_2_7 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_0_LC_7_2_7 .LUT_INIT=16'b1101010101010101;
    LogicCell40 \reset_module_System.count_0_LC_7_2_7  (
            .in0(N__41051),
            .in1(N__41030),
            .in2(N__39660),
            .in3(N__40972),
            .lcout(\reset_module_System.countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87002),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.rudder_esr_5_LC_7_4_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_esr_5_LC_7_4_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.rudder_esr_5_LC_7_4_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.rudder_esr_5_LC_7_4_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39657),
            .lcout(\ppm_encoder_1.rudderZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87017),
            .ce(N__50146),
            .sr(N__79557));
    defparam \uart_pc_sync.aux_1__0__0_LC_7_5_0 .C_ON=1'b0;
    defparam \uart_pc_sync.aux_1__0__0_LC_7_5_0 .SEQ_MODE=4'b1000;
    defparam \uart_pc_sync.aux_1__0__0_LC_7_5_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_pc_sync.aux_1__0__0_LC_7_5_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39630),
            .lcout(\uart_pc_sync.aux_1__0_Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87024),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc_sync.aux_0__0__0_LC_7_5_7 .C_ON=1'b0;
    defparam \uart_pc_sync.aux_0__0__0_LC_7_5_7 .SEQ_MODE=4'b1000;
    defparam \uart_pc_sync.aux_0__0__0_LC_7_5_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_pc_sync.aux_0__0__0_LC_7_5_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39642),
            .lcout(\uart_pc_sync.aux_0__0_Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87024),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc_sync.aux_3__0__0_LC_7_6_0 .C_ON=1'b0;
    defparam \uart_pc_sync.aux_3__0__0_LC_7_6_0 .SEQ_MODE=4'b1000;
    defparam \uart_pc_sync.aux_3__0__0_LC_7_6_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_pc_sync.aux_3__0__0_LC_7_6_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39711),
            .lcout(\uart_pc_sync.aux_3__0_Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87034),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc_sync.aux_2__0__0_LC_7_6_6 .C_ON=1'b0;
    defparam \uart_pc_sync.aux_2__0__0_LC_7_6_6 .SEQ_MODE=4'b1000;
    defparam \uart_pc_sync.aux_2__0__0_LC_7_6_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_pc_sync.aux_2__0__0_LC_7_6_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39717),
            .lcout(\uart_pc_sync.aux_2__0_Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87034),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.rudder_esr_ctle_14_LC_7_7_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_esr_ctle_14_LC_7_7_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.rudder_esr_ctle_14_LC_7_7_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \ppm_encoder_1.rudder_esr_ctle_14_LC_7_7_6  (
            .in0(_gnd_net_),
            .in1(N__65054),
            .in2(_gnd_net_),
            .in3(N__79955),
            .lcout(\ppm_encoder_1.pid_altitude_dv_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_1_LC_7_8_3 .C_ON=1'b0;
    defparam \uart_drone.state_1_LC_7_8_3 .SEQ_MODE=4'b1000;
    defparam \uart_drone.state_1_LC_7_8_3 .LUT_INIT=16'b0101000001000000;
    LogicCell40 \uart_drone.state_1_LC_7_8_3  (
            .in0(N__79958),
            .in1(N__39693),
            .in2(N__47978),
            .in3(N__39702),
            .lcout(\uart_drone.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87054),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_RNO_0_0_LC_7_8_4 .C_ON=1'b0;
    defparam \uart_drone.state_RNO_0_0_LC_7_8_4 .SEQ_MODE=4'b0000;
    defparam \uart_drone.state_RNO_0_0_LC_7_8_4 .LUT_INIT=16'b0000000011011101;
    LogicCell40 \uart_drone.state_RNO_0_0_LC_7_8_4  (
            .in0(N__39701),
            .in1(N__47951),
            .in2(_gnd_net_),
            .in3(N__79957),
            .lcout(),
            .ltout(\uart_drone.state_srsts_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_0_LC_7_8_5 .C_ON=1'b0;
    defparam \uart_drone.state_0_LC_7_8_5 .SEQ_MODE=4'b1000;
    defparam \uart_drone.state_0_LC_7_8_5 .LUT_INIT=16'b1110111100001111;
    LogicCell40 \uart_drone.state_0_LC_7_8_5  (
            .in0(N__50770),
            .in1(N__40069),
            .in2(N__39705),
            .in3(N__44712),
            .lcout(\uart_drone.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87054),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_RNIAT1D1_4_LC_7_8_6 .C_ON=1'b0;
    defparam \uart_drone.state_RNIAT1D1_4_LC_7_8_6 .SEQ_MODE=4'b0000;
    defparam \uart_drone.state_RNIAT1D1_4_LC_7_8_6 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \uart_drone.state_RNIAT1D1_4_LC_7_8_6  (
            .in0(N__44711),
            .in1(N__50769),
            .in2(N__40071),
            .in3(N__79956),
            .lcout(\uart_drone.N_143 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_RNO_0_2_LC_7_9_2 .C_ON=1'b0;
    defparam \uart_drone.state_RNO_0_2_LC_7_9_2 .SEQ_MODE=4'b0000;
    defparam \uart_drone.state_RNO_0_2_LC_7_9_2 .LUT_INIT=16'b0000001000001110;
    LogicCell40 \uart_drone.state_RNO_0_2_LC_7_9_2  (
            .in0(N__44739),
            .in1(N__39691),
            .in2(N__80000),
            .in3(N__47950),
            .lcout(),
            .ltout(\uart_drone.state_srsts_i_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_2_LC_7_9_3 .C_ON=1'b0;
    defparam \uart_drone.state_2_LC_7_9_3 .SEQ_MODE=4'b1000;
    defparam \uart_drone.state_2_LC_7_9_3 .LUT_INIT=16'b1011000011110000;
    LogicCell40 \uart_drone.state_2_LC_7_9_3  (
            .in0(N__39692),
            .in1(N__50823),
            .in2(N__39678),
            .in3(N__50784),
            .lcout(\uart_drone.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87062),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_0_LC_7_9_4 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_0_LC_7_9_4 .SEQ_MODE=4'b1000;
    defparam \uart_drone.timer_Count_0_LC_7_9_4 .LUT_INIT=16'b0000000001010100;
    LogicCell40 \uart_drone.timer_Count_0_LC_7_9_4  (
            .in0(N__79973),
            .in1(N__39797),
            .in2(N__39774),
            .in3(N__39867),
            .lcout(\uart_drone.timer_CountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87062),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_3_LC_7_9_6 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_3_LC_7_9_6 .SEQ_MODE=4'b1000;
    defparam \uart_drone.timer_Count_3_LC_7_9_6 .LUT_INIT=16'b0101010000000000;
    LogicCell40 \uart_drone.timer_Count_3_LC_7_9_6  (
            .in0(N__79974),
            .in1(N__39798),
            .in2(N__39775),
            .in3(N__39849),
            .lcout(\uart_drone.timer_CountZ1Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87062),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_RNI9E9J_2_LC_7_10_0 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_RNI9E9J_2_LC_7_10_0 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNI9E9J_2_LC_7_10_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uart_drone.timer_Count_RNI9E9J_2_LC_7_10_0  (
            .in0(_gnd_net_),
            .in1(N__39839),
            .in2(_gnd_net_),
            .in3(N__50813),
            .lcout(\uart_drone.N_126_li ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_RNIDGR31_2_LC_7_10_1 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_RNIDGR31_2_LC_7_10_1 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNIDGR31_2_LC_7_10_1 .LUT_INIT=16'b1100110010000000;
    LogicCell40 \uart_drone.timer_Count_RNIDGR31_2_LC_7_10_1  (
            .in0(N__50812),
            .in1(N__44699),
            .in2(N__39840),
            .in3(N__50782),
            .lcout(\uart_drone.data_rdyc_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_4_LC_7_10_2 .C_ON=1'b0;
    defparam \uart_drone.state_4_LC_7_10_2 .SEQ_MODE=4'b1000;
    defparam \uart_drone.state_4_LC_7_10_2 .LUT_INIT=16'b1111111101000000;
    LogicCell40 \uart_drone.state_4_LC_7_10_2  (
            .in0(N__79969),
            .in1(N__44966),
            .in2(N__50724),
            .in3(N__39810),
            .lcout(\uart_drone.stateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87074),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_RNIUPE73_3_LC_7_10_3 .C_ON=1'b0;
    defparam \uart_pc.state_RNIUPE73_3_LC_7_10_3 .SEQ_MODE=4'b0000;
    defparam \uart_pc.state_RNIUPE73_3_LC_7_10_3 .LUT_INIT=16'b1010101000100010;
    LogicCell40 \uart_pc.state_RNIUPE73_3_LC_7_10_3  (
            .in0(N__41677),
            .in1(N__41649),
            .in2(_gnd_net_),
            .in3(N__41700),
            .lcout(\uart_pc.un1_state_7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_RNI40411_2_LC_7_10_4 .C_ON=1'b0;
    defparam \uart_drone.state_RNI40411_2_LC_7_10_4 .SEQ_MODE=4'b0000;
    defparam \uart_drone.state_RNI40411_2_LC_7_10_4 .LUT_INIT=16'b0101010011111100;
    LogicCell40 \uart_drone.state_RNI40411_2_LC_7_10_4  (
            .in0(N__50783),
            .in1(N__44965),
            .in2(N__44740),
            .in3(N__50814),
            .lcout(\uart_drone.timer_Count_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_RNO_0_0_LC_7_10_5 .C_ON=1'b0;
    defparam \uart_pc.state_RNO_0_0_LC_7_10_5 .SEQ_MODE=4'b0000;
    defparam \uart_pc.state_RNO_0_0_LC_7_10_5 .LUT_INIT=16'b0000000011011101;
    LogicCell40 \uart_pc.state_RNO_0_0_LC_7_10_5  (
            .in0(N__40031),
            .in1(N__40243),
            .in2(_gnd_net_),
            .in3(N__79968),
            .lcout(),
            .ltout(\uart_pc.state_srsts_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_0_LC_7_10_6 .C_ON=1'b0;
    defparam \uart_pc.state_0_LC_7_10_6 .SEQ_MODE=4'b1000;
    defparam \uart_pc.state_0_LC_7_10_6 .LUT_INIT=16'b1100111110001111;
    LogicCell40 \uart_pc.state_0_LC_7_10_6  (
            .in0(N__40581),
            .in1(N__40560),
            .in2(N__39729),
            .in3(N__40382),
            .lcout(\uart_pc.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87074),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_7_10_7.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_7_10_7.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_7_10_7.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_7_10_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_RNI9ADK1_4_LC_7_11_0 .C_ON=1'b0;
    defparam \uart_drone.state_RNI9ADK1_4_LC_7_11_0 .SEQ_MODE=4'b0000;
    defparam \uart_drone.state_RNI9ADK1_4_LC_7_11_0 .LUT_INIT=16'b1111111101001100;
    LogicCell40 \uart_drone.state_RNI9ADK1_4_LC_7_11_0  (
            .in0(N__40070),
            .in1(N__44972),
            .in2(N__40050),
            .in3(N__44708),
            .lcout(\uart_drone.un1_state_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_1_LC_7_11_3 .C_ON=1'b0;
    defparam \uart_pc.state_1_LC_7_11_3 .SEQ_MODE=4'b1000;
    defparam \uart_pc.state_1_LC_7_11_3 .LUT_INIT=16'b0000000011001000;
    LogicCell40 \uart_pc.state_1_LC_7_11_3  (
            .in0(N__40138),
            .in1(N__40250),
            .in2(N__40035),
            .in3(N__79952),
            .lcout(\uart_pc.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87086),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.bit_Count_RNI4U6E1_2_LC_7_11_5 .C_ON=1'b0;
    defparam \uart_pc.bit_Count_RNI4U6E1_2_LC_7_11_5 .SEQ_MODE=4'b0000;
    defparam \uart_pc.bit_Count_RNI4U6E1_2_LC_7_11_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uart_pc.bit_Count_RNI4U6E1_2_LC_7_11_5  (
            .in0(N__39928),
            .in1(N__39967),
            .in2(_gnd_net_),
            .in3(N__41555),
            .lcout(\uart_pc.N_152 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un2_source_data_0_cry_1_c_RNO_LC_7_11_6 .C_ON=1'b0;
    defparam \scaler_4.un2_source_data_0_cry_1_c_RNO_LC_7_11_6 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un2_source_data_0_cry_1_c_RNO_LC_7_11_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \scaler_4.un2_source_data_0_cry_1_c_RNO_LC_7_11_6  (
            .in0(N__42714),
            .in1(N__42675),
            .in2(_gnd_net_),
            .in3(N__42748),
            .lcout(\scaler_4.un2_source_data_0_cry_1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_RNIOU0N_4_LC_7_11_7 .C_ON=1'b0;
    defparam \uart_drone.state_RNIOU0N_4_LC_7_11_7 .SEQ_MODE=4'b0000;
    defparam \uart_drone.state_RNIOU0N_4_LC_7_11_7 .LUT_INIT=16'b1111111100000101;
    LogicCell40 \uart_drone.state_RNIOU0N_4_LC_7_11_7  (
            .in0(N__44709),
            .in1(_gnd_net_),
            .in2(N__44976),
            .in3(N__79951),
            .lcout(\uart_drone.state_RNIOU0NZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.bit_Count_1_LC_7_12_0 .C_ON=1'b0;
    defparam \uart_pc.bit_Count_1_LC_7_12_0 .SEQ_MODE=4'b1000;
    defparam \uart_pc.bit_Count_1_LC_7_12_0 .LUT_INIT=16'b0000000001101010;
    LogicCell40 \uart_pc.bit_Count_1_LC_7_12_0  (
            .in0(N__39991),
            .in1(N__41567),
            .in2(N__41679),
            .in3(N__40019),
            .lcout(\uart_pc.bit_CountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87102),
            .ce(),
            .sr(N__79588));
    defparam \uart_pc.bit_Count_2_LC_7_12_1 .C_ON=1'b0;
    defparam \uart_pc.bit_Count_2_LC_7_12_1 .SEQ_MODE=4'b1000;
    defparam \uart_pc.bit_Count_2_LC_7_12_1 .LUT_INIT=16'b0001010101000000;
    LogicCell40 \uart_pc.bit_Count_2_LC_7_12_1  (
            .in0(N__40020),
            .in1(N__39992),
            .in2(N__40263),
            .in3(N__39932),
            .lcout(\uart_pc.bit_CountZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87102),
            .ce(),
            .sr(N__79588));
    defparam \uart_pc.state_RNIEAGS_4_LC_7_12_3 .C_ON=1'b0;
    defparam \uart_pc.state_RNIEAGS_4_LC_7_12_3 .SEQ_MODE=4'b0000;
    defparam \uart_pc.state_RNIEAGS_4_LC_7_12_3 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \uart_pc.state_RNIEAGS_4_LC_7_12_3  (
            .in0(N__40559),
            .in1(N__41650),
            .in2(_gnd_net_),
            .in3(N__79927),
            .lcout(\uart_pc.state_RNIEAGSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNISTI31_12_LC_7_12_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNISTI31_12_LC_7_12_5 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNISTI31_12_LC_7_12_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \Commands_frame_decoder.state_RNISTI31_12_LC_7_12_5  (
            .in0(_gnd_net_),
            .in1(N__39897),
            .in2(_gnd_net_),
            .in3(N__79925),
            .lcout(\Commands_frame_decoder.source_xy_ki_1_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_data_valid_2_sqmuxa_i_LC_7_12_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_data_valid_2_sqmuxa_i_LC_7_12_7 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_data_valid_2_sqmuxa_i_LC_7_12_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \dron_frame_decoder_1.source_data_valid_2_sqmuxa_i_LC_7_12_7  (
            .in0(_gnd_net_),
            .in1(N__50964),
            .in2(_gnd_net_),
            .in3(N__79926),
            .lcout(\dron_frame_decoder_1.source_data_valid_2_sqmuxa_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNII68S_9_LC_7_13_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNII68S_9_LC_7_13_0 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNII68S_9_LC_7_13_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \Commands_frame_decoder.state_RNII68S_9_LC_7_13_0  (
            .in0(_gnd_net_),
            .in1(N__40283),
            .in2(_gnd_net_),
            .in3(N__79961),
            .lcout(\Commands_frame_decoder.source_offset4data_1_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_RNIGRIF1_2_LC_7_13_2 .C_ON=1'b0;
    defparam \uart_pc.state_RNIGRIF1_2_LC_7_13_2 .SEQ_MODE=4'b0000;
    defparam \uart_pc.state_RNIGRIF1_2_LC_7_13_2 .LUT_INIT=16'b0101010011111100;
    LogicCell40 \uart_pc.state_RNIGRIF1_2_LC_7_13_2  (
            .in0(N__40370),
            .in1(N__40107),
            .in2(N__41645),
            .in3(N__40427),
            .lcout(\uart_pc.timer_Count_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_RNIITIF1_4_LC_7_13_3 .C_ON=1'b0;
    defparam \uart_pc.state_RNIITIF1_4_LC_7_13_3 .SEQ_MODE=4'b0000;
    defparam \uart_pc.state_RNIITIF1_4_LC_7_13_3 .LUT_INIT=16'b0101000100010001;
    LogicCell40 \uart_pc.state_RNIITIF1_4_LC_7_13_3  (
            .in0(N__40531),
            .in1(N__41629),
            .in2(N__40439),
            .in3(N__40369),
            .lcout(\uart_pc.un1_state_4_0 ),
            .ltout(\uart_pc.un1_state_4_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.bit_Count_RNO_0_2_LC_7_13_4 .C_ON=1'b0;
    defparam \uart_pc.bit_Count_RNO_0_2_LC_7_13_4 .SEQ_MODE=4'b0000;
    defparam \uart_pc.bit_Count_RNO_0_2_LC_7_13_4 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \uart_pc.bit_Count_RNO_0_2_LC_7_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__40266),
            .in3(N__41566),
            .lcout(\uart_pc.CO0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_RNO_0_2_LC_7_13_6 .C_ON=1'b0;
    defparam \uart_pc.state_RNO_0_2_LC_7_13_6 .SEQ_MODE=4'b0000;
    defparam \uart_pc.state_RNO_0_2_LC_7_13_6 .LUT_INIT=16'b0000000000111010;
    LogicCell40 \uart_pc.state_RNO_0_2_LC_7_13_6  (
            .in0(N__40114),
            .in1(N__40237),
            .in2(N__40143),
            .in3(N__79962),
            .lcout(),
            .ltout(\uart_pc.state_srsts_i_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_2_LC_7_13_7 .C_ON=1'b0;
    defparam \uart_pc.state_2_LC_7_13_7 .SEQ_MODE=4'b1000;
    defparam \uart_pc.state_2_LC_7_13_7 .LUT_INIT=16'b1101000011110000;
    LogicCell40 \uart_pc.state_2_LC_7_13_7  (
            .in0(N__40428),
            .in1(N__40142),
            .in2(N__40122),
            .in3(N__40371),
            .lcout(\uart_pc.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87117),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_xy_ki_esr_4_LC_7_14_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_ki_esr_4_LC_7_14_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_ki_esr_4_LC_7_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_xy_ki_esr_4_LC_7_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85027),
            .lcout(xy_ki_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87133),
            .ce(N__78666),
            .sr(N__79600));
    defparam \uart_pc.timer_Count_RNIRP8S_1_LC_7_15_0 .C_ON=1'b1;
    defparam \uart_pc.timer_Count_RNIRP8S_1_LC_7_15_0 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNIRP8S_1_LC_7_15_0 .LUT_INIT=16'b0001000100010001;
    LogicCell40 \uart_pc.timer_Count_RNIRP8S_1_LC_7_15_0  (
            .in0(N__41868),
            .in1(N__40089),
            .in2(N__41873),
            .in3(_gnd_net_),
            .lcout(\uart_pc.un1_state_2_0_a3_0 ),
            .ltout(),
            .carryin(bfn_7_15_0_),
            .carryout(\uart_pc.un4_timer_Count_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNO_0_2_LC_7_15_1 .C_ON=1'b1;
    defparam \uart_pc.timer_Count_RNO_0_2_LC_7_15_1 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNO_0_2_LC_7_15_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_pc.timer_Count_RNO_0_2_LC_7_15_1  (
            .in0(_gnd_net_),
            .in1(N__40312),
            .in2(_gnd_net_),
            .in3(N__40590),
            .lcout(\uart_pc.timer_Count_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(\uart_pc.un4_timer_Count_1_cry_1 ),
            .carryout(\uart_pc.un4_timer_Count_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNO_0_3_LC_7_15_2 .C_ON=1'b1;
    defparam \uart_pc.timer_Count_RNO_0_3_LC_7_15_2 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNO_0_3_LC_7_15_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_pc.timer_Count_RNO_0_3_LC_7_15_2  (
            .in0(_gnd_net_),
            .in1(N__40423),
            .in2(_gnd_net_),
            .in3(N__40587),
            .lcout(\uart_pc.timer_Count_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(\uart_pc.un4_timer_Count_1_cry_2 ),
            .carryout(\uart_pc.un4_timer_Count_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNO_0_4_LC_7_15_3 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_RNO_0_4_LC_7_15_3 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNO_0_4_LC_7_15_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uart_pc.timer_Count_RNO_0_4_LC_7_15_3  (
            .in0(_gnd_net_),
            .in1(N__40365),
            .in2(_gnd_net_),
            .in3(N__40584),
            .lcout(\uart_pc.timer_Count_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_RNIBLRB2_4_LC_7_15_4 .C_ON=1'b0;
    defparam \uart_pc.state_RNIBLRB2_4_LC_7_15_4 .SEQ_MODE=4'b0000;
    defparam \uart_pc.state_RNIBLRB2_4_LC_7_15_4 .LUT_INIT=16'b1101111111001100;
    LogicCell40 \uart_pc.state_RNIBLRB2_4_LC_7_15_4  (
            .in0(N__40577),
            .in1(N__40552),
            .in2(N__40506),
            .in3(N__41651),
            .lcout(\uart_pc.un1_state_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_3_LC_7_15_5 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_3_LC_7_15_5 .SEQ_MODE=4'b1000;
    defparam \uart_pc.timer_Count_3_LC_7_15_5 .LUT_INIT=16'b0000000010101000;
    LogicCell40 \uart_pc.timer_Count_3_LC_7_15_5  (
            .in0(N__40449),
            .in1(N__41956),
            .in2(N__41914),
            .in3(N__79977),
            .lcout(\uart_pc.timer_CountZ1Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87151),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_4_LC_7_15_6 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_4_LC_7_15_6 .SEQ_MODE=4'b1000;
    defparam \uart_pc.timer_Count_4_LC_7_15_6 .LUT_INIT=16'b0101010000000000;
    LogicCell40 \uart_pc.timer_Count_4_LC_7_15_6  (
            .in0(N__79975),
            .in1(N__41906),
            .in2(N__41961),
            .in3(N__40392),
            .lcout(\uart_pc.timer_CountZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87151),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_2_LC_7_15_7 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_2_LC_7_15_7 .SEQ_MODE=4'b1000;
    defparam \uart_pc.timer_Count_2_LC_7_15_7 .LUT_INIT=16'b0000000010101000;
    LogicCell40 \uart_pc.timer_Count_2_LC_7_15_7  (
            .in0(N__40329),
            .in1(N__41955),
            .in2(N__41913),
            .in3(N__79976),
            .lcout(\uart_pc.timer_CountZ1Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87151),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI8NB61_2_11_LC_7_16_1 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI8NB61_2_11_LC_7_16_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI8NB61_2_11_LC_7_16_1 .LUT_INIT=16'b0111011100010001;
    LogicCell40 \pid_front.error_p_reg_esr_RNI8NB61_2_11_LC_7_16_1  (
            .in0(N__49182),
            .in1(N__49128),
            .in2(_gnd_net_),
            .in3(N__49223),
            .lcout(\pid_front.g0_1_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_esr_RNIUHO16_12_LC_7_16_4 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_esr_RNIUHO16_12_LC_7_16_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_esr_RNIUHO16_12_LC_7_16_4 .LUT_INIT=16'b0100010011001100;
    LogicCell40 \pid_front.pid_prereg_esr_RNIUHO16_12_LC_7_16_4  (
            .in0(N__45654),
            .in1(N__45690),
            .in2(_gnd_net_),
            .in3(N__45608),
            .lcout(\pid_front.N_76 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_esr_RNIOL7G1_8_LC_7_16_6 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_esr_RNIOL7G1_8_LC_7_16_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_esr_RNIOL7G1_8_LC_7_16_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \pid_front.pid_prereg_esr_RNIOL7G1_8_LC_7_16_6  (
            .in0(N__45653),
            .in1(N__43425),
            .in2(N__41835),
            .in3(N__45548),
            .lcout(\pid_front.N_99 ),
            .ltout(\pid_front.N_99_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_esr_RNI3Q532_4_LC_7_16_7 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_esr_RNI3Q532_4_LC_7_16_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_esr_RNI3Q532_4_LC_7_16_7 .LUT_INIT=16'b0101000001000000;
    LogicCell40 \pid_front.pid_prereg_esr_RNI3Q532_4_LC_7_16_7  (
            .in0(N__45384),
            .in1(N__43224),
            .in2(N__40632),
            .in3(N__43256),
            .lcout(\pid_front.N_75 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_0_LC_7_18_0 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_0_LC_7_18_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_0_LC_7_18_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_0_LC_7_18_0  (
            .in0(_gnd_net_),
            .in1(N__66243),
            .in2(_gnd_net_),
            .in3(N__66261),
            .lcout(\pid_side.error_i_acumm_preregZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87195),
            .ce(N__69901),
            .sr(N__79624));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNIKAP4_8_LC_7_18_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNIKAP4_8_LC_7_18_1 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNIKAP4_8_LC_7_18_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_RNIKAP4_8_LC_7_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48498),
            .lcout(drone_H_disp_side_i_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNILBP4_9_LC_7_18_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNILBP4_9_LC_7_18_2 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNILBP4_9_LC_7_18_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_RNILBP4_9_LC_7_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48489),
            .lcout(drone_H_disp_side_i_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNIT4RD_10_LC_7_18_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNIT4RD_10_LC_7_18_3 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNIT4RD_10_LC_7_18_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_RNIT4RD_10_LC_7_18_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48195),
            .lcout(drone_H_disp_side_i_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_axb_12_LC_7_18_5 .C_ON=1'b0;
    defparam \pid_alt.error_axb_12_LC_7_18_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_axb_12_LC_7_18_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_alt.error_axb_12_LC_7_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40683),
            .lcout(\pid_alt.error_axbZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_axb_13_LC_7_18_6 .C_ON=1'b0;
    defparam \pid_alt.error_axb_13_LC_7_18_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_axb_13_LC_7_18_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_alt.error_axb_13_LC_7_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40677),
            .lcout(\pid_alt.error_axbZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_axb_14_LC_7_18_7 .C_ON=1'b0;
    defparam \pid_alt.error_axb_14_LC_7_18_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_axb_14_LC_7_18_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pid_alt.error_axb_14_LC_7_18_7  (
            .in0(N__40671),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_axbZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_10_LC_7_19_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_10_LC_7_19_0 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_10_LC_7_19_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_10_LC_7_19_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59106),
            .lcout(\dron_frame_decoder_1.drone_altitude_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87212),
            .ce(N__47733),
            .sr(N__79631));
    defparam \dron_frame_decoder_1.source_Altitude_esr_11_LC_7_19_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_11_LC_7_19_1 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_11_LC_7_19_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_11_LC_7_19_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59025),
            .lcout(\dron_frame_decoder_1.drone_altitude_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87212),
            .ce(N__47733),
            .sr(N__79631));
    defparam \dron_frame_decoder_1.source_Altitude_esr_12_LC_7_19_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_12_LC_7_19_2 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_12_LC_7_19_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_12_LC_7_19_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58930),
            .lcout(drone_altitude_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87212),
            .ce(N__47733),
            .sr(N__79631));
    defparam \dron_frame_decoder_1.source_Altitude_esr_13_LC_7_19_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_13_LC_7_19_3 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_13_LC_7_19_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_13_LC_7_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58841),
            .lcout(drone_altitude_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87212),
            .ce(N__47733),
            .sr(N__79631));
    defparam \dron_frame_decoder_1.source_Altitude_esr_14_LC_7_19_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_14_LC_7_19_4 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_14_LC_7_19_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_14_LC_7_19_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58757),
            .lcout(drone_altitude_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87212),
            .ce(N__47733),
            .sr(N__79631));
    defparam \dron_frame_decoder_1.source_Altitude_esr_15_LC_7_19_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_15_LC_7_19_5 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_15_LC_7_19_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_15_LC_7_19_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58643),
            .lcout(drone_altitude_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87212),
            .ce(N__47733),
            .sr(N__79631));
    defparam \dron_frame_decoder_1.source_Altitude_esr_8_LC_7_19_6 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_8_LC_7_19_6 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_8_LC_7_19_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_8_LC_7_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59333),
            .lcout(\dron_frame_decoder_1.drone_altitude_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87212),
            .ce(N__47733),
            .sr(N__79631));
    defparam \dron_frame_decoder_1.source_Altitude_esr_9_LC_7_19_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_9_LC_7_19_7 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_9_LC_7_19_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_9_LC_7_19_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59205),
            .lcout(\dron_frame_decoder_1.drone_altitude_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87212),
            .ce(N__47733),
            .sr(N__79631));
    defparam \pid_front.pid_prereg_esr_RNIIH1A1_24_LC_7_20_3 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_esr_RNIIH1A1_24_LC_7_20_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_esr_RNIIH1A1_24_LC_7_20_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_front.pid_prereg_esr_RNIIH1A1_24_LC_7_20_3  (
            .in0(N__43677),
            .in1(N__43695),
            .in2(N__43650),
            .in3(N__43443),
            .lcout(\pid_front.un11lto30_i_a2_5_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_1_cry_1_c_LC_8_1_0 .C_ON=1'b1;
    defparam \reset_module_System.count_1_cry_1_c_LC_8_1_0 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_1_cry_1_c_LC_8_1_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \reset_module_System.count_1_cry_1_c_LC_8_1_0  (
            .in0(_gnd_net_),
            .in1(N__41049),
            .in2(N__40950),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_1_0_),
            .carryout(\reset_module_System.count_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNO_0_2_LC_8_1_1 .C_ON=1'b1;
    defparam \reset_module_System.count_RNO_0_2_LC_8_1_1 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNO_0_2_LC_8_1_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_RNO_0_2_LC_8_1_1  (
            .in0(_gnd_net_),
            .in1(N__40820),
            .in2(_gnd_net_),
            .in3(N__40803),
            .lcout(\reset_module_System.count_1_2 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_1 ),
            .carryout(\reset_module_System.count_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_3_LC_8_1_2 .C_ON=1'b1;
    defparam \reset_module_System.count_3_LC_8_1_2 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_3_LC_8_1_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_3_LC_8_1_2  (
            .in0(_gnd_net_),
            .in1(N__40800),
            .in2(_gnd_net_),
            .in3(N__40788),
            .lcout(\reset_module_System.countZ0Z_3 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_2 ),
            .carryout(\reset_module_System.count_1_cry_3 ),
            .clk(N__86989),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_4_LC_8_1_3 .C_ON=1'b1;
    defparam \reset_module_System.count_4_LC_8_1_3 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_4_LC_8_1_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_4_LC_8_1_3  (
            .in0(_gnd_net_),
            .in1(N__40784),
            .in2(_gnd_net_),
            .in3(N__40773),
            .lcout(\reset_module_System.countZ0Z_4 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_3 ),
            .carryout(\reset_module_System.count_1_cry_4 ),
            .clk(N__86989),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_5_LC_8_1_4 .C_ON=1'b1;
    defparam \reset_module_System.count_5_LC_8_1_4 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_5_LC_8_1_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_5_LC_8_1_4  (
            .in0(_gnd_net_),
            .in1(N__40770),
            .in2(_gnd_net_),
            .in3(N__40758),
            .lcout(\reset_module_System.countZ0Z_5 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_4 ),
            .carryout(\reset_module_System.count_1_cry_5 ),
            .clk(N__86989),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_6_LC_8_1_5 .C_ON=1'b1;
    defparam \reset_module_System.count_6_LC_8_1_5 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_6_LC_8_1_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_6_LC_8_1_5  (
            .in0(_gnd_net_),
            .in1(N__40755),
            .in2(_gnd_net_),
            .in3(N__40743),
            .lcout(\reset_module_System.countZ0Z_6 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_5 ),
            .carryout(\reset_module_System.count_1_cry_6 ),
            .clk(N__86989),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_7_LC_8_1_6 .C_ON=1'b1;
    defparam \reset_module_System.count_7_LC_8_1_6 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_7_LC_8_1_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_7_LC_8_1_6  (
            .in0(_gnd_net_),
            .in1(N__40740),
            .in2(_gnd_net_),
            .in3(N__40728),
            .lcout(\reset_module_System.countZ0Z_7 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_6 ),
            .carryout(\reset_module_System.count_1_cry_7 ),
            .clk(N__86989),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_8_LC_8_1_7 .C_ON=1'b1;
    defparam \reset_module_System.count_8_LC_8_1_7 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_8_LC_8_1_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_8_LC_8_1_7  (
            .in0(_gnd_net_),
            .in1(N__40725),
            .in2(_gnd_net_),
            .in3(N__40713),
            .lcout(\reset_module_System.countZ0Z_8 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_7 ),
            .carryout(\reset_module_System.count_1_cry_8 ),
            .clk(N__86989),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_9_LC_8_2_0 .C_ON=1'b1;
    defparam \reset_module_System.count_9_LC_8_2_0 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_9_LC_8_2_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_9_LC_8_2_0  (
            .in0(_gnd_net_),
            .in1(N__40709),
            .in2(_gnd_net_),
            .in3(N__40695),
            .lcout(\reset_module_System.countZ0Z_9 ),
            .ltout(),
            .carryin(bfn_8_2_0_),
            .carryout(\reset_module_System.count_1_cry_9 ),
            .clk(N__86998),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_10_LC_8_2_1 .C_ON=1'b1;
    defparam \reset_module_System.count_10_LC_8_2_1 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_10_LC_8_2_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_10_LC_8_2_1  (
            .in0(_gnd_net_),
            .in1(N__41163),
            .in2(_gnd_net_),
            .in3(N__40923),
            .lcout(\reset_module_System.countZ0Z_10 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_9 ),
            .carryout(\reset_module_System.count_1_cry_10 ),
            .clk(N__86998),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_11_LC_8_2_2 .C_ON=1'b1;
    defparam \reset_module_System.count_11_LC_8_2_2 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_11_LC_8_2_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_11_LC_8_2_2  (
            .in0(_gnd_net_),
            .in1(N__41151),
            .in2(_gnd_net_),
            .in3(N__40920),
            .lcout(\reset_module_System.countZ0Z_11 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_10 ),
            .carryout(\reset_module_System.count_1_cry_11 ),
            .clk(N__86998),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_12_LC_8_2_3 .C_ON=1'b1;
    defparam \reset_module_System.count_12_LC_8_2_3 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_12_LC_8_2_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_12_LC_8_2_3  (
            .in0(_gnd_net_),
            .in1(N__40913),
            .in2(_gnd_net_),
            .in3(N__40902),
            .lcout(\reset_module_System.countZ0Z_12 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_11 ),
            .carryout(\reset_module_System.count_1_cry_12 ),
            .clk(N__86998),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_13_LC_8_2_4 .C_ON=1'b1;
    defparam \reset_module_System.count_13_LC_8_2_4 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_13_LC_8_2_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_13_LC_8_2_4  (
            .in0(_gnd_net_),
            .in1(N__41087),
            .in2(_gnd_net_),
            .in3(N__40899),
            .lcout(\reset_module_System.countZ0Z_13 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_12 ),
            .carryout(\reset_module_System.count_1_cry_13 ),
            .clk(N__86998),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_14_LC_8_2_5 .C_ON=1'b1;
    defparam \reset_module_System.count_14_LC_8_2_5 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_14_LC_8_2_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_14_LC_8_2_5  (
            .in0(_gnd_net_),
            .in1(N__40896),
            .in2(_gnd_net_),
            .in3(N__40884),
            .lcout(\reset_module_System.countZ0Z_14 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_13 ),
            .carryout(\reset_module_System.count_1_cry_14 ),
            .clk(N__86998),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_15_LC_8_2_6 .C_ON=1'b1;
    defparam \reset_module_System.count_15_LC_8_2_6 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_15_LC_8_2_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_15_LC_8_2_6  (
            .in0(_gnd_net_),
            .in1(N__41117),
            .in2(_gnd_net_),
            .in3(N__40881),
            .lcout(\reset_module_System.countZ0Z_15 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_14 ),
            .carryout(\reset_module_System.count_1_cry_15 ),
            .clk(N__86998),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_16_LC_8_2_7 .C_ON=1'b1;
    defparam \reset_module_System.count_16_LC_8_2_7 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_16_LC_8_2_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_16_LC_8_2_7  (
            .in0(_gnd_net_),
            .in1(N__40874),
            .in2(_gnd_net_),
            .in3(N__40863),
            .lcout(\reset_module_System.countZ0Z_16 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_15 ),
            .carryout(\reset_module_System.count_1_cry_16 ),
            .clk(N__86998),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_17_LC_8_3_0 .C_ON=1'b1;
    defparam \reset_module_System.count_17_LC_8_3_0 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_17_LC_8_3_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_17_LC_8_3_0  (
            .in0(_gnd_net_),
            .in1(N__40859),
            .in2(_gnd_net_),
            .in3(N__40845),
            .lcout(\reset_module_System.countZ0Z_17 ),
            .ltout(),
            .carryin(bfn_8_3_0_),
            .carryout(\reset_module_System.count_1_cry_17 ),
            .clk(N__87003),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_18_LC_8_3_1 .C_ON=1'b1;
    defparam \reset_module_System.count_18_LC_8_3_1 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_18_LC_8_3_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_18_LC_8_3_1  (
            .in0(_gnd_net_),
            .in1(N__40841),
            .in2(_gnd_net_),
            .in3(N__40827),
            .lcout(\reset_module_System.countZ0Z_18 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_17 ),
            .carryout(\reset_module_System.count_1_cry_18 ),
            .clk(N__87003),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_19_LC_8_3_2 .C_ON=1'b1;
    defparam \reset_module_System.count_19_LC_8_3_2 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_19_LC_8_3_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_19_LC_8_3_2  (
            .in0(_gnd_net_),
            .in1(N__41133),
            .in2(_gnd_net_),
            .in3(N__41187),
            .lcout(\reset_module_System.countZ0Z_19 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_18 ),
            .carryout(\reset_module_System.count_1_cry_19 ),
            .clk(N__87003),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_20_LC_8_3_3 .C_ON=1'b1;
    defparam \reset_module_System.count_20_LC_8_3_3 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_20_LC_8_3_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_20_LC_8_3_3  (
            .in0(_gnd_net_),
            .in1(N__41183),
            .in2(_gnd_net_),
            .in3(N__41169),
            .lcout(\reset_module_System.countZ0Z_20 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_19 ),
            .carryout(\reset_module_System.count_1_cry_20 ),
            .clk(N__87003),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_21_LC_8_3_4 .C_ON=1'b0;
    defparam \reset_module_System.count_21_LC_8_3_4 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_21_LC_8_3_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \reset_module_System.count_21_LC_8_3_4  (
            .in0(_gnd_net_),
            .in1(N__41105),
            .in2(_gnd_net_),
            .in3(N__41166),
            .lcout(\reset_module_System.countZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87003),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNIP8RT_10_LC_8_3_6 .C_ON=1'b0;
    defparam \reset_module_System.count_RNIP8RT_10_LC_8_3_6 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNIP8RT_10_LC_8_3_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \reset_module_System.count_RNIP8RT_10_LC_8_3_6  (
            .in0(_gnd_net_),
            .in1(N__41162),
            .in2(_gnd_net_),
            .in3(N__41150),
            .lcout(\reset_module_System.reset6_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNI34OR1_21_LC_8_4_0 .C_ON=1'b0;
    defparam \reset_module_System.count_RNI34OR1_21_LC_8_4_0 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNI34OR1_21_LC_8_4_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \reset_module_System.count_RNI34OR1_21_LC_8_4_0  (
            .in0(N__41132),
            .in1(N__41121),
            .in2(N__41106),
            .in3(N__41091),
            .lcout(\reset_module_System.reset6_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone_sync.aux_0__0__0_LC_8_4_3 .C_ON=1'b0;
    defparam \uart_drone_sync.aux_0__0__0_LC_8_4_3 .SEQ_MODE=4'b1000;
    defparam \uart_drone_sync.aux_0__0__0_LC_8_4_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone_sync.aux_0__0__0_LC_8_4_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41076),
            .lcout(\uart_drone_sync.aux_0__0__0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87010),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNO_0_1_LC_8_5_2 .C_ON=1'b0;
    defparam \reset_module_System.count_RNO_0_1_LC_8_5_2 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNO_0_1_LC_8_5_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \reset_module_System.count_RNO_0_1_LC_8_5_2  (
            .in0(_gnd_net_),
            .in1(N__41055),
            .in2(_gnd_net_),
            .in3(N__40945),
            .lcout(),
            .ltout(\reset_module_System.count_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_1_LC_8_5_3 .C_ON=1'b0;
    defparam \reset_module_System.count_1_LC_8_5_3 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_1_LC_8_5_3 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \reset_module_System.count_1_LC_8_5_3  (
            .in0(N__41017),
            .in1(N__41001),
            .in2(N__40983),
            .in3(N__40980),
            .lcout(\reset_module_System.countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87018),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_5_LC_8_6_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_5_LC_8_6_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_5_LC_8_6_0 .LUT_INIT=16'b0000010100100010;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_5_LC_8_6_0  (
            .in0(N__61619),
            .in1(N__42145),
            .in2(N__44553),
            .in3(N__61419),
            .lcout(\ppm_encoder_1.pulses2count_9_i_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_5_LC_8_6_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_5_LC_8_6_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_5_LC_8_6_2 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.throttle_5_LC_8_6_2  (
            .in0(N__41256),
            .in1(N__41292),
            .in2(N__65296),
            .in3(N__42146),
            .lcout(\ppm_encoder_1.throttleZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87025),
            .ce(),
            .sr(N__79560));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_9_LC_8_6_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_9_LC_8_6_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_9_LC_8_6_3 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_9_LC_8_6_3  (
            .in0(N__61418),
            .in1(N__61618),
            .in2(_gnd_net_),
            .in3(N__47116),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_2Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_9_LC_8_6_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_9_LC_8_6_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_9_LC_8_6_4 .LUT_INIT=16'b0011101011001010;
    LogicCell40 \ppm_encoder_1.throttle_9_LC_8_6_4  (
            .in0(N__47117),
            .in1(N__41235),
            .in2(N__65297),
            .in3(N__41208),
            .lcout(\ppm_encoder_1.throttleZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87025),
            .ce(),
            .sr(N__79560));
    defparam \ppm_encoder_1.rudder_6_LC_8_6_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_6_LC_8_6_6 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.rudder_6_LC_8_6_6 .LUT_INIT=16'b0111011100100010;
    LogicCell40 \ppm_encoder_1.rudder_6_LC_8_6_6  (
            .in0(N__65248),
            .in1(N__42357),
            .in2(_gnd_net_),
            .in3(N__57781),
            .lcout(\ppm_encoder_1.rudderZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87025),
            .ce(),
            .sr(N__79560));
    defparam \ppm_encoder_1.throttle_11_LC_8_7_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_11_LC_8_7_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_11_LC_8_7_1 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.throttle_11_LC_8_7_1  (
            .in0(N__41502),
            .in1(N__41469),
            .in2(N__65290),
            .in3(N__57361),
            .lcout(\ppm_encoder_1.throttleZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87035),
            .ce(),
            .sr(N__79565));
    defparam \ppm_encoder_1.throttle_3_LC_8_7_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_3_LC_8_7_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_3_LC_8_7_7 .LUT_INIT=16'b1001111110010000;
    LogicCell40 \ppm_encoder_1.throttle_3_LC_8_7_7  (
            .in0(N__41325),
            .in1(N__41304),
            .in2(N__65291),
            .in3(N__68584),
            .lcout(\ppm_encoder_1.throttleZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87035),
            .ce(),
            .sr(N__79565));
    defparam \ppm_encoder_1.un1_throttle_cry_0_c_LC_8_8_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_0_c_LC_8_8_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_0_c_LC_8_8_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_0_c_LC_8_8_0  (
            .in0(_gnd_net_),
            .in1(N__53156),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_8_0_),
            .carryout(\ppm_encoder_1.un1_throttle_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_0_THRU_LUT4_0_LC_8_8_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_0_THRU_LUT4_0_LC_8_8_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_0_THRU_LUT4_0_LC_8_8_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_0_THRU_LUT4_0_LC_8_8_1  (
            .in0(_gnd_net_),
            .in1(N__50315),
            .in2(N__56523),
            .in3(N__41193),
            .lcout(\ppm_encoder_1.un1_throttle_cry_0_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_0 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_1_THRU_LUT4_0_LC_8_8_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_1_THRU_LUT4_0_LC_8_8_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_1_THRU_LUT4_0_LC_8_8_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_1_THRU_LUT4_0_LC_8_8_2  (
            .in0(_gnd_net_),
            .in1(N__44570),
            .in2(_gnd_net_),
            .in3(N__41190),
            .lcout(\ppm_encoder_1.un1_throttle_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_1 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_2_THRU_LUT4_0_LC_8_8_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_2_THRU_LUT4_0_LC_8_8_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_2_THRU_LUT4_0_LC_8_8_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_2_THRU_LUT4_0_LC_8_8_3  (
            .in0(_gnd_net_),
            .in1(N__41321),
            .in2(N__56524),
            .in3(N__41298),
            .lcout(\ppm_encoder_1.un1_throttle_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_2 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_3_THRU_LUT4_0_LC_8_8_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_3_THRU_LUT4_0_LC_8_8_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_3_THRU_LUT4_0_LC_8_8_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_3_THRU_LUT4_0_LC_8_8_4  (
            .in0(_gnd_net_),
            .in1(N__42315),
            .in2(_gnd_net_),
            .in3(N__41295),
            .lcout(\ppm_encoder_1.un1_throttle_cry_3_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_3 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_4_THRU_LUT4_0_LC_8_8_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_4_THRU_LUT4_0_LC_8_8_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_4_THRU_LUT4_0_LC_8_8_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_4_THRU_LUT4_0_LC_8_8_5  (
            .in0(_gnd_net_),
            .in1(N__41291),
            .in2(_gnd_net_),
            .in3(N__41247),
            .lcout(\ppm_encoder_1.un1_throttle_cry_4_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_4 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_5_THRU_LUT4_0_LC_8_8_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_5_THRU_LUT4_0_LC_8_8_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_5_THRU_LUT4_0_LC_8_8_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_5_THRU_LUT4_0_LC_8_8_6  (
            .in0(_gnd_net_),
            .in1(N__56459),
            .in2(N__41439),
            .in3(N__41244),
            .lcout(\ppm_encoder_1.un1_throttle_cry_5_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_5 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_6_THRU_LUT4_0_LC_8_8_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_6_THRU_LUT4_0_LC_8_8_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_6_THRU_LUT4_0_LC_8_8_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_6_THRU_LUT4_0_LC_8_8_7  (
            .in0(_gnd_net_),
            .in1(N__47189),
            .in2(_gnd_net_),
            .in3(N__41241),
            .lcout(\ppm_encoder_1.un1_throttle_cry_6_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_6 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_7_THRU_LUT4_0_LC_8_9_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_7_THRU_LUT4_0_LC_8_9_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_7_THRU_LUT4_0_LC_8_9_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_7_THRU_LUT4_0_LC_8_9_0  (
            .in0(_gnd_net_),
            .in1(N__41409),
            .in2(_gnd_net_),
            .in3(N__41238),
            .lcout(\ppm_encoder_1.un1_throttle_cry_7_THRU_CO ),
            .ltout(),
            .carryin(bfn_8_9_0_),
            .carryout(\ppm_encoder_1.un1_throttle_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_8_THRU_LUT4_0_LC_8_9_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_8_THRU_LUT4_0_LC_8_9_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_8_THRU_LUT4_0_LC_8_9_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_8_THRU_LUT4_0_LC_8_9_1  (
            .in0(_gnd_net_),
            .in1(N__41231),
            .in2(_gnd_net_),
            .in3(N__41199),
            .lcout(\ppm_encoder_1.un1_throttle_cry_8_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_8 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_9_THRU_LUT4_0_LC_8_9_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_9_THRU_LUT4_0_LC_8_9_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_9_THRU_LUT4_0_LC_8_9_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_9_THRU_LUT4_0_LC_8_9_2  (
            .in0(_gnd_net_),
            .in1(N__44657),
            .in2(_gnd_net_),
            .in3(N__41196),
            .lcout(\ppm_encoder_1.un1_throttle_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_9 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_10_THRU_LUT4_0_LC_8_9_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_10_THRU_LUT4_0_LC_8_9_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_10_THRU_LUT4_0_LC_8_9_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_10_THRU_LUT4_0_LC_8_9_3  (
            .in0(_gnd_net_),
            .in1(N__41501),
            .in2(_gnd_net_),
            .in3(N__41460),
            .lcout(\ppm_encoder_1.un1_throttle_cry_10_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_10 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_11_THRU_LUT4_0_LC_8_9_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_11_THRU_LUT4_0_LC_8_9_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_11_THRU_LUT4_0_LC_8_9_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_11_THRU_LUT4_0_LC_8_9_4  (
            .in0(_gnd_net_),
            .in1(N__47258),
            .in2(_gnd_net_),
            .in3(N__41457),
            .lcout(\ppm_encoder_1.un1_throttle_cry_11_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_11 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_12_THRU_LUT4_0_LC_8_9_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_12_THRU_LUT4_0_LC_8_9_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_12_THRU_LUT4_0_LC_8_9_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_12_THRU_LUT4_0_LC_8_9_5  (
            .in0(_gnd_net_),
            .in1(N__44621),
            .in2(N__56507),
            .in3(N__41454),
            .lcout(\ppm_encoder_1.un1_throttle_cry_12_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_12 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_esr_14_LC_8_9_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_esr_14_LC_8_9_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_esr_14_LC_8_9_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.throttle_esr_14_LC_8_9_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41451),
            .lcout(\ppm_encoder_1.throttleZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87055),
            .ce(N__50158),
            .sr(N__79574));
    defparam \ppm_encoder_1.throttle_6_LC_8_10_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_6_LC_8_10_1 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.throttle_6_LC_8_10_1 .LUT_INIT=16'b1001100111110000;
    LogicCell40 \ppm_encoder_1.throttle_6_LC_8_10_1  (
            .in0(N__41448),
            .in1(N__41435),
            .in2(N__61762),
            .in3(N__65267),
            .lcout(\ppm_encoder_1.throttleZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87063),
            .ce(),
            .sr(N__79582));
    defparam \ppm_encoder_1.throttle_8_LC_8_10_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_8_LC_8_10_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_8_LC_8_10_2 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.throttle_8_LC_8_10_2  (
            .in0(N__41407),
            .in1(N__41379),
            .in2(N__65303),
            .in3(N__60703),
            .lcout(\ppm_encoder_1.throttleZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87063),
            .ce(),
            .sr(N__79582));
    defparam \scaler_4.source_data_1_4_LC_8_10_3 .C_ON=1'b0;
    defparam \scaler_4.source_data_1_4_LC_8_10_3 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_4_LC_8_10_3 .LUT_INIT=16'b0111001011011000;
    LogicCell40 \scaler_4.source_data_1_4_LC_8_10_3  (
            .in0(N__41363),
            .in1(N__42749),
            .in2(N__50177),
            .in3(N__42722),
            .lcout(scaler_4_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87063),
            .ce(),
            .sr(N__79582));
    defparam \scaler_4.source_data_1_esr_ctle_14_LC_8_10_4 .C_ON=1'b0;
    defparam \scaler_4.source_data_1_esr_ctle_14_LC_8_10_4 .SEQ_MODE=4'b0000;
    defparam \scaler_4.source_data_1_esr_ctle_14_LC_8_10_4 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \scaler_4.source_data_1_esr_ctle_14_LC_8_10_4  (
            .in0(N__79954),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41362),
            .lcout(\scaler_4.debug_CH3_20A_c_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_RNIES9Q1_2_LC_8_10_5 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_RNIES9Q1_2_LC_8_10_5 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNIES9Q1_2_LC_8_10_5 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \uart_drone.timer_Count_RNIES9Q1_2_LC_8_10_5  (
            .in0(N__47943),
            .in1(N__47893),
            .in2(_gnd_net_),
            .in3(N__79953),
            .lcout(\uart_drone.timer_Count_RNIES9Q1Z0Z_2 ),
            .ltout(\uart_drone.timer_Count_RNIES9Q1Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_RNIRC5U2_2_LC_8_10_6 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_RNIRC5U2_2_LC_8_10_6 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNIRC5U2_2_LC_8_10_6 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \uart_drone.timer_Count_RNIRC5U2_2_LC_8_10_6  (
            .in0(N__47894),
            .in1(_gnd_net_),
            .in2(N__41718),
            .in3(_gnd_net_),
            .lcout(\uart_drone.data_rdyc_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.bit_Count_0_LC_8_10_7 .C_ON=1'b0;
    defparam \uart_pc.bit_Count_0_LC_8_10_7 .SEQ_MODE=4'b1000;
    defparam \uart_pc.bit_Count_0_LC_8_10_7 .LUT_INIT=16'b0011001101000000;
    LogicCell40 \uart_pc.bit_Count_0_LC_8_10_7  (
            .in0(N__41707),
            .in1(N__41678),
            .in2(N__41652),
            .in3(N__41565),
            .lcout(\uart_pc.bit_CountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87063),
            .ce(),
            .sr(N__79582));
    defparam \Commands_frame_decoder.source_CH4data_esr_0_LC_8_11_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH4data_esr_0_LC_8_11_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH4data_esr_0_LC_8_11_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH4data_esr_0_LC_8_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__83794),
            .lcout(frame_decoder_CH4data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87075),
            .ce(N__41532),
            .sr(N__79589));
    defparam \Commands_frame_decoder.source_CH4data_esr_1_LC_8_11_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH4data_esr_1_LC_8_11_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH4data_esr_1_LC_8_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH4data_esr_1_LC_8_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84161),
            .lcout(frame_decoder_CH4data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87075),
            .ce(N__41532),
            .sr(N__79589));
    defparam \Commands_frame_decoder.source_CH4data_esr_2_LC_8_11_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH4data_esr_2_LC_8_11_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH4data_esr_2_LC_8_11_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH4data_esr_2_LC_8_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__77549),
            .lcout(frame_decoder_CH4data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87075),
            .ce(N__41532),
            .sr(N__79589));
    defparam \Commands_frame_decoder.source_CH4data_esr_3_LC_8_11_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH4data_esr_3_LC_8_11_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH4data_esr_3_LC_8_11_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH4data_esr_3_LC_8_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__83988),
            .lcout(frame_decoder_CH4data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87075),
            .ce(N__41532),
            .sr(N__79589));
    defparam \Commands_frame_decoder.source_CH4data_esr_4_LC_8_11_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH4data_esr_4_LC_8_11_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH4data_esr_4_LC_8_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH4data_esr_4_LC_8_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84979),
            .lcout(frame_decoder_CH4data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87075),
            .ce(N__41532),
            .sr(N__79589));
    defparam \Commands_frame_decoder.source_CH4data_esr_5_LC_8_11_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH4data_esr_5_LC_8_11_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH4data_esr_5_LC_8_11_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Commands_frame_decoder.source_CH4data_esr_5_LC_8_11_5  (
            .in0(N__85199),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(frame_decoder_CH4data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87075),
            .ce(N__41532),
            .sr(N__79589));
    defparam \Commands_frame_decoder.source_CH4data_esr_6_LC_8_11_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH4data_esr_6_LC_8_11_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH4data_esr_6_LC_8_11_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH4data_esr_6_LC_8_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73638),
            .lcout(frame_decoder_CH4data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87075),
            .ce(N__41532),
            .sr(N__79589));
    defparam \Commands_frame_decoder.source_offset4data_esr_0_LC_8_12_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset4data_esr_0_LC_8_12_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset4data_esr_0_LC_8_12_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset4data_esr_0_LC_8_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__83796),
            .lcout(frame_decoder_OFF4data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87087),
            .ce(N__41748),
            .sr(N__79594));
    defparam \Commands_frame_decoder.source_offset4data_esr_1_LC_8_12_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset4data_esr_1_LC_8_12_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset4data_esr_1_LC_8_12_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset4data_esr_1_LC_8_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84147),
            .lcout(frame_decoder_OFF4data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87087),
            .ce(N__41748),
            .sr(N__79594));
    defparam \Commands_frame_decoder.source_offset4data_esr_2_LC_8_12_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset4data_esr_2_LC_8_12_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset4data_esr_2_LC_8_12_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset4data_esr_2_LC_8_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__77520),
            .lcout(frame_decoder_OFF4data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87087),
            .ce(N__41748),
            .sr(N__79594));
    defparam \Commands_frame_decoder.source_offset4data_esr_3_LC_8_12_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset4data_esr_3_LC_8_12_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset4data_esr_3_LC_8_12_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Commands_frame_decoder.source_offset4data_esr_3_LC_8_12_3  (
            .in0(N__83968),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(frame_decoder_OFF4data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87087),
            .ce(N__41748),
            .sr(N__79594));
    defparam \Commands_frame_decoder.source_offset4data_esr_4_LC_8_12_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset4data_esr_4_LC_8_12_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset4data_esr_4_LC_8_12_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset4data_esr_4_LC_8_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85026),
            .lcout(frame_decoder_OFF4data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87087),
            .ce(N__41748),
            .sr(N__79594));
    defparam \Commands_frame_decoder.source_offset4data_esr_5_LC_8_12_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset4data_esr_5_LC_8_12_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset4data_esr_5_LC_8_12_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset4data_esr_5_LC_8_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85158),
            .lcout(frame_decoder_OFF4data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87087),
            .ce(N__41748),
            .sr(N__79594));
    defparam \Commands_frame_decoder.source_offset4data_esr_6_LC_8_12_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset4data_esr_6_LC_8_12_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset4data_esr_6_LC_8_12_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset4data_esr_6_LC_8_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73639),
            .lcout(frame_decoder_OFF4data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87087),
            .ce(N__41748),
            .sr(N__79594));
    defparam \Commands_frame_decoder.source_offset4data_ess_7_LC_8_12_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset4data_ess_7_LC_8_12_7 .SEQ_MODE=4'b1001;
    defparam \Commands_frame_decoder.source_offset4data_ess_7_LC_8_12_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset4data_ess_7_LC_8_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85364),
            .lcout(frame_decoder_OFF4data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87087),
            .ce(N__41748),
            .sr(N__79594));
    defparam \dron_frame_decoder_1.WDT_0_LC_8_13_0 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_0_LC_8_13_0 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_0_LC_8_13_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_0_LC_8_13_0  (
            .in0(_gnd_net_),
            .in1(N__41733),
            .in2(N__42873),
            .in3(N__42872),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_0 ),
            .ltout(),
            .carryin(bfn_8_13_0_),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_0 ),
            .clk(N__87103),
            .ce(),
            .sr(N__41811));
    defparam \dron_frame_decoder_1.WDT_1_LC_8_13_1 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_1_LC_8_13_1 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_1_LC_8_13_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_1_LC_8_13_1  (
            .in0(_gnd_net_),
            .in1(N__41727),
            .in2(_gnd_net_),
            .in3(N__41721),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_1 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_0 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_1 ),
            .clk(N__87103),
            .ce(),
            .sr(N__41811));
    defparam \dron_frame_decoder_1.WDT_2_LC_8_13_2 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_2_LC_8_13_2 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_2_LC_8_13_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_2_LC_8_13_2  (
            .in0(_gnd_net_),
            .in1(N__41787),
            .in2(_gnd_net_),
            .in3(N__41781),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_2 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_1 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_2 ),
            .clk(N__87103),
            .ce(),
            .sr(N__41811));
    defparam \dron_frame_decoder_1.WDT_3_LC_8_13_3 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_3_LC_8_13_3 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_3_LC_8_13_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_3_LC_8_13_3  (
            .in0(_gnd_net_),
            .in1(N__41778),
            .in2(_gnd_net_),
            .in3(N__41772),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_3 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_2 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_3 ),
            .clk(N__87103),
            .ce(),
            .sr(N__41811));
    defparam \dron_frame_decoder_1.WDT_4_LC_8_13_4 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_4_LC_8_13_4 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_4_LC_8_13_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_4_LC_8_13_4  (
            .in0(_gnd_net_),
            .in1(N__42888),
            .in2(_gnd_net_),
            .in3(N__41769),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_4 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_3 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_4 ),
            .clk(N__87103),
            .ce(),
            .sr(N__41811));
    defparam \dron_frame_decoder_1.WDT_5_LC_8_13_5 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_5_LC_8_13_5 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_5_LC_8_13_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_5_LC_8_13_5  (
            .in0(_gnd_net_),
            .in1(N__42915),
            .in2(_gnd_net_),
            .in3(N__41766),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_5 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_4 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_5 ),
            .clk(N__87103),
            .ce(),
            .sr(N__41811));
    defparam \dron_frame_decoder_1.WDT_6_LC_8_13_6 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_6_LC_8_13_6 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_6_LC_8_13_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_6_LC_8_13_6  (
            .in0(_gnd_net_),
            .in1(N__42858),
            .in2(_gnd_net_),
            .in3(N__41763),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_6 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_5 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_6 ),
            .clk(N__87103),
            .ce(),
            .sr(N__41811));
    defparam \dron_frame_decoder_1.WDT_7_LC_8_13_7 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_7_LC_8_13_7 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_7_LC_8_13_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_7_LC_8_13_7  (
            .in0(_gnd_net_),
            .in1(N__42846),
            .in2(_gnd_net_),
            .in3(N__41760),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_7 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_6 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_7 ),
            .clk(N__87103),
            .ce(),
            .sr(N__41811));
    defparam \dron_frame_decoder_1.WDT_8_LC_8_14_0 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_8_LC_8_14_0 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_8_LC_8_14_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_8_LC_8_14_0  (
            .in0(_gnd_net_),
            .in1(N__42929),
            .in2(_gnd_net_),
            .in3(N__41757),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_8 ),
            .ltout(),
            .carryin(bfn_8_14_0_),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_8 ),
            .clk(N__87118),
            .ce(),
            .sr(N__41810));
    defparam \dron_frame_decoder_1.WDT_9_LC_8_14_1 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_9_LC_8_14_1 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_9_LC_8_14_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_9_LC_8_14_1  (
            .in0(_gnd_net_),
            .in1(N__42902),
            .in2(_gnd_net_),
            .in3(N__41754),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_9 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_8 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_9 ),
            .clk(N__87118),
            .ce(),
            .sr(N__41810));
    defparam \dron_frame_decoder_1.WDT_10_LC_8_14_2 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_10_LC_8_14_2 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_10_LC_8_14_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_10_LC_8_14_2  (
            .in0(_gnd_net_),
            .in1(N__42833),
            .in2(_gnd_net_),
            .in3(N__41751),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_10 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_9 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_10 ),
            .clk(N__87118),
            .ce(),
            .sr(N__41810));
    defparam \dron_frame_decoder_1.WDT_11_LC_8_14_3 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_11_LC_8_14_3 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_11_LC_8_14_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_11_LC_8_14_3  (
            .in0(_gnd_net_),
            .in1(N__42807),
            .in2(_gnd_net_),
            .in3(N__41826),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_11 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_10 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_11 ),
            .clk(N__87118),
            .ce(),
            .sr(N__41810));
    defparam \dron_frame_decoder_1.WDT_12_LC_8_14_4 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_12_LC_8_14_4 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_12_LC_8_14_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_12_LC_8_14_4  (
            .in0(_gnd_net_),
            .in1(N__42768),
            .in2(_gnd_net_),
            .in3(N__41823),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_12 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_11 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_12 ),
            .clk(N__87118),
            .ce(),
            .sr(N__41810));
    defparam \dron_frame_decoder_1.WDT_13_LC_8_14_5 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_13_LC_8_14_5 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_13_LC_8_14_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_13_LC_8_14_5  (
            .in0(_gnd_net_),
            .in1(N__42792),
            .in2(_gnd_net_),
            .in3(N__41820),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_13 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_12 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_13 ),
            .clk(N__87118),
            .ce(),
            .sr(N__41810));
    defparam \dron_frame_decoder_1.WDT_14_LC_8_14_6 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_14_LC_8_14_6 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_14_LC_8_14_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_14_LC_8_14_6  (
            .in0(_gnd_net_),
            .in1(N__43064),
            .in2(_gnd_net_),
            .in3(N__41817),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_14 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_13 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_14 ),
            .clk(N__87118),
            .ce(),
            .sr(N__41810));
    defparam \dron_frame_decoder_1.WDT_15_LC_8_14_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.WDT_15_LC_8_14_7 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_15_LC_8_14_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \dron_frame_decoder_1.WDT_15_LC_8_14_7  (
            .in0(_gnd_net_),
            .in1(N__43047),
            .in2(_gnd_net_),
            .in3(N__41814),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87118),
            .ce(),
            .sr(N__41810));
    defparam \pid_front.un11lto30_i_a2_0_c_LC_8_15_0 .C_ON=1'b1;
    defparam \pid_front.un11lto30_i_a2_0_c_LC_8_15_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.un11lto30_i_a2_0_c_LC_8_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_front.un11lto30_i_a2_0_c_LC_8_15_0  (
            .in0(_gnd_net_),
            .in1(N__43104),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_15_0_),
            .carryout(\pid_front.un11lto30_i_a2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un11lto30_i_a2_1_c_LC_8_15_1 .C_ON=1'b1;
    defparam \pid_front.un11lto30_i_a2_1_c_LC_8_15_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.un11lto30_i_a2_1_c_LC_8_15_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_front.un11lto30_i_a2_1_c_LC_8_15_1  (
            .in0(_gnd_net_),
            .in1(N__42036),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pid_front.un11lto30_i_a2 ),
            .carryout(\pid_front.un11lto30_i_a2_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un11lto30_i_a2_2_c_LC_8_15_2 .C_ON=1'b1;
    defparam \pid_front.un11lto30_i_a2_2_c_LC_8_15_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.un11lto30_i_a2_2_c_LC_8_15_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_front.un11lto30_i_a2_2_c_LC_8_15_2  (
            .in0(_gnd_net_),
            .in1(N__42045),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pid_front.un11lto30_i_a2_0 ),
            .carryout(\pid_front.un11lto30_i_a2_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un11lto30_i_a2_3_c_LC_8_15_3 .C_ON=1'b1;
    defparam \pid_front.un11lto30_i_a2_3_c_LC_8_15_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.un11lto30_i_a2_3_c_LC_8_15_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_front.un11lto30_i_a2_3_c_LC_8_15_3  (
            .in0(_gnd_net_),
            .in1(N__42027),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pid_front.un11lto30_i_a2_1 ),
            .carryout(\pid_front.un11lto30_i_a2_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un11lto30_i_a2_4_c_LC_8_15_4 .C_ON=1'b1;
    defparam \pid_front.un11lto30_i_a2_4_c_LC_8_15_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.un11lto30_i_a2_4_c_LC_8_15_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_front.un11lto30_i_a2_4_c_LC_8_15_4  (
            .in0(_gnd_net_),
            .in1(N__41846),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pid_front.un11lto30_i_a2_2 ),
            .carryout(\pid_front.un11lto30_i_a2_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un11lto30_i_a2_5_c_LC_8_15_5 .C_ON=1'b1;
    defparam \pid_front.un11lto30_i_a2_5_c_LC_8_15_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.un11lto30_i_a2_5_c_LC_8_15_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_front.un11lto30_i_a2_5_c_LC_8_15_5  (
            .in0(_gnd_net_),
            .in1(N__42003),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pid_front.un11lto30_i_a2_3 ),
            .carryout(\pid_front.un11lto30_i_a2_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un11lto30_i_a2_6_c_LC_8_15_6 .C_ON=1'b1;
    defparam \pid_front.un11lto30_i_a2_6_c_LC_8_15_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.un11lto30_i_a2_6_c_LC_8_15_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_front.un11lto30_i_a2_6_c_LC_8_15_6  (
            .in0(_gnd_net_),
            .in1(N__41994),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pid_front.un11lto30_i_a2_4 ),
            .carryout(\pid_front.un11lto30_i_a2_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un11lto30_i_a2_7_c_LC_8_15_7 .C_ON=1'b1;
    defparam \pid_front.un11lto30_i_a2_7_c_LC_8_15_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.un11lto30_i_a2_7_c_LC_8_15_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_front.un11lto30_i_a2_7_c_LC_8_15_7  (
            .in0(_gnd_net_),
            .in1(N__43016),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pid_front.un11lto30_i_a2_5 ),
            .carryout(\pid_front.un11lto30_i_a2_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un11lto30_i_a2_7_c_RNI57AF1_LC_8_16_0 .C_ON=1'b0;
    defparam \pid_front.un11lto30_i_a2_7_c_RNI57AF1_LC_8_16_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.un11lto30_i_a2_7_c_RNI57AF1_LC_8_16_0 .LUT_INIT=16'b0000100000001111;
    LogicCell40 \pid_front.un11lto30_i_a2_7_c_RNI57AF1_LC_8_16_0  (
            .in0(N__45655),
            .in1(N__45598),
            .in2(N__45383),
            .in3(N__41964),
            .lcout(\pid_front.source_pid_1_sqmuxa_1_0_o2_sx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_esr_RNIMHT91_16_LC_8_16_1 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_esr_RNIMHT91_16_LC_8_16_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_esr_RNIMHT91_16_LC_8_16_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_front.pid_prereg_esr_RNIMHT91_16_LC_8_16_1  (
            .in0(N__43353),
            .in1(N__43539),
            .in2(N__43557),
            .in3(N__43527),
            .lcout(\pid_front.un11lto30_i_a2_3_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_0_LC_8_16_3 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_0_LC_8_16_3 .SEQ_MODE=4'b1000;
    defparam \uart_pc.timer_Count_0_LC_8_16_3 .LUT_INIT=16'b0000000000110010;
    LogicCell40 \uart_pc.timer_Count_0_LC_8_16_3  (
            .in0(N__41960),
            .in1(N__41872),
            .in2(N__41915),
            .in3(N__79994),
            .lcout(\uart_pc.timer_CountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87152),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_esr_RNI295P1_15_LC_8_16_7 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_esr_RNI295P1_15_LC_8_16_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_esr_RNI295P1_15_LC_8_16_7 .LUT_INIT=16'b0000010100000000;
    LogicCell40 \pid_front.pid_prereg_esr_RNI295P1_15_LC_8_16_7  (
            .in0(N__42018),
            .in1(_gnd_net_),
            .in2(N__43374),
            .in3(N__41847),
            .lcout(\pid_front.source_pid_1_sqmuxa_1_0_a2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_esr_RNI4ABT_6_LC_8_17_0 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_esr_RNI4ABT_6_LC_8_17_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_esr_RNI4ABT_6_LC_8_17_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \pid_front.pid_prereg_esr_RNI4ABT_6_LC_8_17_0  (
            .in0(N__43186),
            .in1(N__43157),
            .in2(N__45500),
            .in3(N__45254),
            .lcout(\pid_front.source_pid_1_sqmuxa_1_0_a2_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un11lto30_i_a2_2_c_RNO_LC_8_17_2 .C_ON=1'b0;
    defparam \pid_front.un11lto30_i_a2_2_c_RNO_LC_8_17_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.un11lto30_i_a2_2_c_RNO_LC_8_17_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_front.un11lto30_i_a2_2_c_RNO_LC_8_17_2  (
            .in0(N__45535),
            .in1(N__43414),
            .in2(N__45499),
            .in3(N__45253),
            .lcout(\pid_front.N_11_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un11lto30_i_a2_1_c_RNO_LC_8_17_3 .C_ON=1'b0;
    defparam \pid_front.un11lto30_i_a2_1_c_RNO_LC_8_17_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.un11lto30_i_a2_1_c_RNO_LC_8_17_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_front.un11lto30_i_a2_1_c_RNO_LC_8_17_3  (
            .in0(N__43156),
            .in1(N__43212),
            .in2(N__43188),
            .in3(N__43242),
            .lcout(\pid_front.un11lto30_i_a2_0_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_esr_RNI6TRI_0_LC_8_17_4 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_esr_RNI6TRI_0_LC_8_17_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_esr_RNI6TRI_0_LC_8_17_4 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \pid_front.pid_prereg_esr_RNI6TRI_0_LC_8_17_4  (
            .in0(N__43243),
            .in1(N__45588),
            .in2(_gnd_net_),
            .in3(N__43337),
            .lcout(\pid_front.source_pid_1_sqmuxa_1_0_a4_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un11lto30_i_a2_3_c_RNO_LC_8_17_5 .C_ON=1'b0;
    defparam \pid_front.un11lto30_i_a2_3_c_RNO_LC_8_17_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.un11lto30_i_a2_3_c_RNO_LC_8_17_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_front.un11lto30_i_a2_3_c_RNO_LC_8_17_5  (
            .in0(N__45587),
            .in1(N__43370),
            .in2(N__45638),
            .in3(N__42016),
            .lcout(\pid_front.un11lto30_i_a2_2_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_14_LC_8_17_6 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_14_LC_8_17_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_14_LC_8_17_6 .LUT_INIT=16'b0011101011001010;
    LogicCell40 \pid_front.pid_prereg_14_LC_8_17_6  (
            .in0(N__42017),
            .in1(N__48699),
            .in2(N__60196),
            .in3(N__43383),
            .lcout(\pid_front.pid_preregZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87167),
            .ce(),
            .sr(N__79625));
    defparam \pid_front.error_p_reg_esr_RNIV7CQ2_8_LC_8_18_0 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIV7CQ2_8_LC_8_18_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIV7CQ2_8_LC_8_18_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_front.error_p_reg_esr_RNIV7CQ2_8_LC_8_18_0  (
            .in0(N__46035),
            .in1(N__48018),
            .in2(N__47799),
            .in3(N__55042),
            .lcout(\pid_front.error_p_reg_esr_RNIV7CQ2Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_prereg_esr_9_LC_8_18_1 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_9_LC_8_18_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_9_LC_8_18_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_9_LC_8_18_1  (
            .in0(N__55043),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_i_acumm_preregZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87181),
            .ce(N__56084),
            .sr(N__79632));
    defparam \pid_front.pid_prereg_esr_RNI211A1_20_LC_8_18_3 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_esr_RNI211A1_20_LC_8_18_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_esr_RNI211A1_20_LC_8_18_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_front.pid_prereg_esr_RNI211A1_20_LC_8_18_3  (
            .in0(N__43467),
            .in1(N__43485),
            .in2(N__43458),
            .in3(N__43509),
            .lcout(\pid_front.un11lto30_i_a2_4_and ),
            .ltout(\pid_front.un11lto30_i_a2_4_and_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_esr_RNID3QC5_15_LC_8_18_4 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_esr_RNID3QC5_15_LC_8_18_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_esr_RNID3QC5_15_LC_8_18_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \pid_front.pid_prereg_esr_RNID3QC5_15_LC_8_18_4  (
            .in0(N__41993),
            .in1(N__43023),
            .in2(N__41976),
            .in3(N__41973),
            .lcout(\pid_front.N_98 ),
            .ltout(\pid_front.N_98_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_esr_RNIA6N08_0_LC_8_18_5 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_esr_RNIA6N08_0_LC_8_18_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_esr_RNIA6N08_0_LC_8_18_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \pid_front.pid_prereg_esr_RNIA6N08_0_LC_8_18_5  (
            .in0(N__42084),
            .in1(N__43113),
            .in2(N__42078),
            .in3(N__43127),
            .lcout(\pid_front.N_389 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI20QN6_19_LC_8_19_0 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI20QN6_19_LC_8_19_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI20QN6_19_LC_8_19_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \pid_front.error_p_reg_esr_RNI20QN6_19_LC_8_19_0  (
            .in0(_gnd_net_),
            .in1(N__45992),
            .in2(_gnd_net_),
            .in3(N__45974),
            .lcout(\pid_front.error_p_reg_esr_RNI20QN6Z0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIF0FB3_0_19_LC_8_19_1 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIF0FB3_0_19_LC_8_19_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIF0FB3_0_19_LC_8_19_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_front.error_p_reg_esr_RNIF0FB3_0_19_LC_8_19_1  (
            .in0(N__48206),
            .in1(N__49262),
            .in2(_gnd_net_),
            .in3(N__55250),
            .lcout(\pid_front.un1_pid_prereg_0_9 ),
            .ltout(\pid_front.un1_pid_prereg_0_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIQOPM6_18_LC_8_19_2 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIQOPM6_18_LC_8_19_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIQOPM6_18_LC_8_19_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \pid_front.error_p_reg_esr_RNIQOPM6_18_LC_8_19_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__42075),
            .in3(N__42068),
            .lcout(\pid_front.error_p_reg_esr_RNIQOPM6Z0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIF0FB3_19_LC_8_19_3 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIF0FB3_19_LC_8_19_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIF0FB3_19_LC_8_19_3 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_front.error_p_reg_esr_RNIF0FB3_19_LC_8_19_3  (
            .in0(N__48207),
            .in1(N__49263),
            .in2(_gnd_net_),
            .in3(N__55251),
            .lcout(\pid_front.un1_pid_prereg_0_10 ),
            .ltout(\pid_front.un1_pid_prereg_0_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNISOJED_18_LC_8_19_4 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNISOJED_18_LC_8_19_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNISOJED_18_LC_8_19_4 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \pid_front.error_p_reg_esr_RNISOJED_18_LC_8_19_4  (
            .in0(N__42057),
            .in1(N__42069),
            .in2(N__42072),
            .in3(N__45973),
            .lcout(\pid_front.error_p_reg_esr_RNISOJEDZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIBOAB3_18_LC_8_19_5 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIBOAB3_18_LC_8_19_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIBOAB3_18_LC_8_19_5 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_front.error_p_reg_esr_RNIBOAB3_18_LC_8_19_5  (
            .in0(N__51720),
            .in1(N__70539),
            .in2(_gnd_net_),
            .in3(N__55287),
            .lcout(\pid_front.un1_pid_prereg_0_8 ),
            .ltout(\pid_front.un1_pid_prereg_0_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI80EDD_17_LC_8_19_6 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI80EDD_17_LC_8_19_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI80EDD_17_LC_8_19_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \pid_front.error_p_reg_esr_RNI80EDD_17_LC_8_19_6  (
            .in0(N__51966),
            .in1(N__51696),
            .in2(N__42060),
            .in3(N__42056),
            .lcout(\pid_front.error_p_reg_esr_RNI80EDDZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIJVAC3_0_20_LC_8_19_7 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIJVAC3_0_20_LC_8_19_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIJVAC3_0_20_LC_8_19_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_front.error_p_reg_esr_RNIJVAC3_0_20_LC_8_19_7  (
            .in0(N__48381),
            .in1(N__48354),
            .in2(_gnd_net_),
            .in3(N__55728),
            .lcout(\pid_front.un1_pid_prereg_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNINM162_0_22_LC_8_20_0 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNINM162_0_22_LC_8_20_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNINM162_0_22_LC_8_20_0 .LUT_INIT=16'b0001100011100111;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNINM162_0_22_LC_8_20_0  (
            .in0(N__87418),
            .in1(N__48314),
            .in2(N__46335),
            .in3(N__55634),
            .lcout(\pid_front.un1_pid_prereg_0_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNINM162_22_LC_8_20_1 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNINM162_22_LC_8_20_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNINM162_22_LC_8_20_1 .LUT_INIT=16'b1011101010100010;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNINM162_22_LC_8_20_1  (
            .in0(N__55635),
            .in1(N__46312),
            .in2(N__48334),
            .in3(N__87419),
            .lcout(\pid_front.un1_pid_prereg_0_22 ),
            .ltout(\pid_front.un1_pid_prereg_0_22_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNISQ6O8_22_LC_8_20_2 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNISQ6O8_22_LC_8_20_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNISQ6O8_22_LC_8_20_2 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNISQ6O8_22_LC_8_20_2  (
            .in0(N__42114),
            .in1(N__42126),
            .in2(N__42129),
            .in3(N__42166),
            .lcout(\pid_front.error_d_reg_prev_esr_RNISQ6O8Z0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNICA2C4_22_LC_8_20_3 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNICA2C4_22_LC_8_20_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNICA2C4_22_LC_8_20_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNICA2C4_22_LC_8_20_3  (
            .in0(_gnd_net_),
            .in1(N__42113),
            .in2(_gnd_net_),
            .in3(N__42125),
            .lcout(\pid_front.error_d_reg_prev_esr_RNICA2C4Z0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNILJ062_22_LC_8_20_4 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNILJ062_22_LC_8_20_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNILJ062_22_LC_8_20_4 .LUT_INIT=16'b1110111100001000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNILJ062_22_LC_8_20_4  (
            .in0(N__87417),
            .in1(N__48313),
            .in2(N__46334),
            .in3(N__56295),
            .lcout(\pid_front.un1_pid_prereg_0_20 ),
            .ltout(\pid_front.un1_pid_prereg_0_20_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIKE2O8_22_LC_8_20_5 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIKE2O8_22_LC_8_20_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIKE2O8_22_LC_8_20_5 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIKE2O8_22_LC_8_20_5  (
            .in0(N__43731),
            .in1(N__42112),
            .in2(N__42102),
            .in3(N__43746),
            .lcout(\pid_front.error_d_reg_prev_esr_RNIKE2O8Z0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIGG4C4_22_LC_8_20_6 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIGG4C4_22_LC_8_20_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIGG4C4_22_LC_8_20_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIGG4C4_22_LC_8_20_6  (
            .in0(_gnd_net_),
            .in1(N__42095),
            .in2(_gnd_net_),
            .in3(N__42167),
            .lcout(\pid_front.error_d_reg_prev_esr_RNIGG4C4Z0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_22_LC_8_20_7 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_22_LC_8_20_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_22_LC_8_20_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_22_LC_8_20_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__87420),
            .lcout(\pid_front.error_d_reg_prevZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87213),
            .ce(N__70483),
            .sr(N__70354));
    defparam \pid_front.error_d_reg_prev_esr_RNI36BO8_22_LC_8_21_0 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNI36BO8_22_LC_8_21_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNI36BO8_22_LC_8_21_0 .LUT_INIT=16'b0110011001100110;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNI36BO8_22_LC_8_21_0  (
            .in0(N__42218),
            .in1(N__42185),
            .in2(N__42171),
            .in3(N__42099),
            .lcout(\pid_front.error_d_reg_prev_esr_RNI36BO8Z0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIPP262_22_LC_8_21_1 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIPP262_22_LC_8_21_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIPP262_22_LC_8_21_1 .LUT_INIT=16'b1110111100001000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIPP262_22_LC_8_21_1  (
            .in0(N__87424),
            .in1(N__48318),
            .in2(N__46336),
            .in3(N__56210),
            .lcout(\pid_front.un1_pid_prereg_0_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIQR362_0_22_LC_8_21_2 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIQR362_0_22_LC_8_21_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIQR362_0_22_LC_8_21_2 .LUT_INIT=16'b0010010011011011;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIQR362_0_22_LC_8_21_2  (
            .in0(N__87422),
            .in1(N__46322),
            .in2(N__48335),
            .in3(N__55520),
            .lcout(\pid_front.un1_pid_prereg_0_25 ),
            .ltout(\pid_front.un1_pid_prereg_0_25_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIJL6C4_22_LC_8_21_3 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIJL6C4_22_LC_8_21_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIJL6C4_22_LC_8_21_3 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIJL6C4_22_LC_8_21_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__42222),
            .in3(N__42217),
            .lcout(\pid_front.error_d_reg_prev_esr_RNIJL6C4Z0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNI7DEO8_22_LC_8_21_4 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNI7DEO8_22_LC_8_21_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNI7DEO8_22_LC_8_21_4 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNI7DEO8_22_LC_8_21_4  (
            .in0(N__42219),
            .in1(N__42189),
            .in2(N__42206),
            .in3(N__42186),
            .lcout(\pid_front.error_d_reg_prev_esr_RNI7DEO8Z0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIQR362_22_LC_8_21_5 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIQR362_22_LC_8_21_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIQR362_22_LC_8_21_5 .LUT_INIT=16'b1010111010001010;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIQR362_22_LC_8_21_5  (
            .in0(N__55521),
            .in1(N__48320),
            .in2(N__46338),
            .in3(N__87421),
            .lcout(\pid_front.un1_pid_prereg_0_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_esr_RNO_0_30_LC_8_21_6 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_esr_RNO_0_30_LC_8_21_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_esr_RNO_0_30_LC_8_21_6 .LUT_INIT=16'b1000011101111000;
    LogicCell40 \pid_front.pid_prereg_esr_RNO_0_30_LC_8_21_6  (
            .in0(N__42202),
            .in1(N__42187),
            .in2(N__42207),
            .in3(N__42188),
            .lcout(\pid_front.un1_pid_prereg_0_axb_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIPP262_0_22_LC_8_21_7 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIPP262_0_22_LC_8_21_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIPP262_0_22_LC_8_21_7 .LUT_INIT=16'b0001100011100111;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIPP262_0_22_LC_8_21_7  (
            .in0(N__87423),
            .in1(N__48319),
            .in2(N__46337),
            .in3(N__56211),
            .lcout(\pid_front.un1_pid_prereg_0_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.state_RNIVIRQ_0_0_LC_8_22_7 .C_ON=1'b0;
    defparam \pid_front.state_RNIVIRQ_0_0_LC_8_22_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.state_RNIVIRQ_0_0_LC_8_22_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \pid_front.state_RNIVIRQ_0_0_LC_8_22_7  (
            .in0(_gnd_net_),
            .in1(N__67519),
            .in2(_gnd_net_),
            .in3(N__79941),
            .lcout(\pid_front.state_ns_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI8NB61_1_11_LC_8_24_5 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI8NB61_1_11_LC_8_24_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI8NB61_1_11_LC_8_24_5 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_front.error_p_reg_esr_RNI8NB61_1_11_LC_8_24_5  (
            .in0(N__49177),
            .in1(N__49118),
            .in2(_gnd_net_),
            .in3(N__49224),
            .lcout(\pid_front.error_p_reg_esr_RNI8NB61_1Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNISKK21_5_LC_9_2_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNISKK21_5_LC_9_2_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNISKK21_5_LC_9_2_0 .LUT_INIT=16'b1111000001111000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNISKK21_5_LC_9_2_0  (
            .in0(N__63806),
            .in1(N__57710),
            .in2(N__59666),
            .in3(N__64256),
            .lcout(\ppm_encoder_1.N_261_i_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIJL0E1_5_LC_9_2_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIJL0E1_5_LC_9_2_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIJL0E1_5_LC_9_2_1 .LUT_INIT=16'b0011101100001010;
    LogicCell40 \ppm_encoder_1.throttle_RNIJL0E1_5_LC_9_2_1  (
            .in0(N__58012),
            .in1(N__44552),
            .in2(N__42153),
            .in3(N__57185),
            .lcout(\ppm_encoder_1.un2_throttle_iv_0_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNIC96O_5_LC_9_2_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNIC96O_5_LC_9_2_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNIC96O_5_LC_9_2_2 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \ppm_encoder_1.elevator_RNIC96O_5_LC_9_2_2  (
            .in0(N__42233),
            .in1(N__52826),
            .in2(_gnd_net_),
            .in3(N__52943),
            .lcout(\ppm_encoder_1.elevator_RNIC96OZ0Z_5 ),
            .ltout(\ppm_encoder_1.elevator_RNIC96OZ0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.rudder_esr_RNI2S0I2_5_LC_9_2_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_esr_RNI2S0I2_5_LC_9_2_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.rudder_esr_RNI2S0I2_5_LC_9_2_3 .LUT_INIT=16'b1111111111110100;
    LogicCell40 \ppm_encoder_1.rudder_esr_RNI2S0I2_5_LC_9_2_3  (
            .in0(N__60455),
            .in1(N__63807),
            .in2(N__42249),
            .in3(N__57068),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_1_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNI003R4_5_LC_9_2_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI003R4_5_LC_9_2_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI003R4_5_LC_9_2_4 .LUT_INIT=16'b1010100101010110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI003R4_5_LC_9_2_4  (
            .in0(N__59661),
            .in1(N__42246),
            .in2(N__42240),
            .in3(N__56946),
            .lcout(),
            .ltout(\ppm_encoder_1.un1_init_pulses_0_axb_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNISKNT5_5_LC_9_2_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNISKNT5_5_LC_9_2_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNISKNT5_5_LC_9_2_5 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNISKNT5_5_LC_9_2_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__42237),
            .in3(N__44309),
            .lcout(\ppm_encoder_1.init_pulses_RNISKNT5Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_5_LC_9_2_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_5_LC_9_2_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.elevator_5_LC_9_2_6 .LUT_INIT=16'b0011101011001010;
    LogicCell40 \ppm_encoder_1.elevator_5_LC_9_2_6  (
            .in0(N__42234),
            .in1(N__45087),
            .in2(N__65307),
            .in3(N__45111),
            .lcout(\ppm_encoder_1.elevatorZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__86990),
            .ce(),
            .sr(N__79558));
    defparam \ppm_encoder_1.init_pulses_RNI1OK21_0_8_LC_9_3_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI1OK21_0_8_LC_9_3_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI1OK21_0_8_LC_9_3_0 .LUT_INIT=16'b1001110011001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI1OK21_0_8_LC_9_3_0  (
            .in0(N__64263),
            .in1(N__60235),
            .in2(N__60942),
            .in3(N__61056),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNI0NK21_0_7_LC_9_3_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI0NK21_0_7_LC_9_3_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI0NK21_0_7_LC_9_3_1 .LUT_INIT=16'b1111000001111000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI0NK21_0_7_LC_9_3_1  (
            .in0(N__61055),
            .in1(N__60933),
            .in2(N__56715),
            .in3(N__64262),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNIFC6O_8_LC_9_3_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNIFC6O_8_LC_9_3_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNIFC6O_8_LC_9_3_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \ppm_encoder_1.elevator_RNIFC6O_8_LC_9_3_2  (
            .in0(N__47163),
            .in1(N__52827),
            .in2(_gnd_net_),
            .in3(N__52944),
            .lcout(),
            .ltout(\ppm_encoder_1.elevator_RNIFC6OZ0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.rudder_RNI00TI2_8_LC_9_3_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_RNI00TI2_8_LC_9_3_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.rudder_RNI00TI2_8_LC_9_3_3 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \ppm_encoder_1.rudder_RNI00TI2_8_LC_9_3_3  (
            .in0(N__60683),
            .in1(N__60934),
            .in2(N__42225),
            .in3(N__57069),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_2_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNI7DVR4_8_LC_9_3_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI7DVR4_8_LC_9_3_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI7DVR4_8_LC_9_3_4 .LUT_INIT=16'b0110011001101001;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI7DVR4_8_LC_9_3_4  (
            .in0(N__60231),
            .in1(N__56949),
            .in2(N__42270),
            .in3(N__42264),
            .lcout(),
            .ltout(\ppm_encoder_1.un1_init_pulses_0_axb_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNI85KU5_8_LC_9_3_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI85KU5_8_LC_9_3_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI85KU5_8_LC_9_3_5 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI85KU5_8_LC_9_3_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__42267),
            .in3(N__44258),
            .lcout(\ppm_encoder_1.init_pulses_RNI85KU5Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIPR0E1_8_LC_9_3_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIPR0E1_8_LC_9_3_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIPR0E1_8_LC_9_3_6 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \ppm_encoder_1.throttle_RNIPR0E1_8_LC_9_3_6  (
            .in0(N__47445),
            .in1(N__58013),
            .in2(N__60716),
            .in3(N__57186),
            .lcout(\ppm_encoder_1.un2_throttle_iv_0_1_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNI1OK21_8_LC_9_3_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI1OK21_8_LC_9_3_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI1OK21_8_LC_9_3_7 .LUT_INIT=16'b1111000001111000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI1OK21_8_LC_9_3_7  (
            .in0(N__61054),
            .in1(N__60932),
            .in2(N__60239),
            .in3(N__64261),
            .lcout(\ppm_encoder_1.N_264_i_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNIO4K62_3_LC_9_4_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNIO4K62_3_LC_9_4_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNIO4K62_3_LC_9_4_0 .LUT_INIT=16'b1111111110111010;
    LogicCell40 \ppm_encoder_1.elevator_RNIO4K62_3_LC_9_4_0  (
            .in0(N__63797),
            .in1(N__63594),
            .in2(N__52865),
            .in3(N__57059),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_2_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIG2MF4_3_LC_9_4_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIG2MF4_3_LC_9_4_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIG2MF4_3_LC_9_4_1 .LUT_INIT=16'b0110011001101001;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIG2MF4_3_LC_9_4_1  (
            .in0(N__53230),
            .in1(N__56935),
            .in2(N__42258),
            .in3(N__44325),
            .lcout(),
            .ltout(\ppm_encoder_1.un1_init_pulses_0_axb_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIALAI5_3_LC_9_4_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIALAI5_3_LC_9_4_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIALAI5_3_LC_9_4_2 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIALAI5_3_LC_9_4_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__42255),
            .in3(N__44156),
            .lcout(\ppm_encoder_1.init_pulses_RNIALAI5Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIQIK21_3_LC_9_4_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIQIK21_3_LC_9_4_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIQIK21_3_LC_9_4_3 .LUT_INIT=16'b1111000001111000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIQIK21_3_LC_9_4_3  (
            .in0(N__63795),
            .in1(N__57702),
            .in2(N__53232),
            .in3(N__64167),
            .lcout(\ppm_encoder_1.N_256_i_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIRQ2R4_4_LC_9_4_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIRQ2R4_4_LC_9_4_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIRQ2R4_4_LC_9_4_5 .LUT_INIT=16'b0110011001101001;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIRQ2R4_4_LC_9_4_5  (
            .in0(N__59715),
            .in1(N__56936),
            .in2(N__42336),
            .in3(N__50193),
            .lcout(),
            .ltout(\ppm_encoder_1.un1_init_pulses_0_axb_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIMENT5_4_LC_9_4_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIMENT5_4_LC_9_4_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIMENT5_4_LC_9_4_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIMENT5_4_LC_9_4_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__42252),
            .in3(N__44126),
            .lcout(\ppm_encoder_1.init_pulses_RNIMENT5Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIRJK21_4_LC_9_4_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIRJK21_4_LC_9_4_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIRJK21_4_LC_9_4_7 .LUT_INIT=16'b1111000001111000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIRJK21_4_LC_9_4_7  (
            .in0(N__63796),
            .in1(N__57703),
            .in2(N__59718),
            .in3(N__64168),
            .lcout(\ppm_encoder_1.N_260_i_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_4_LC_9_5_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_4_LC_9_5_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_4_LC_9_5_0 .LUT_INIT=16'b0001000011010000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_4_LC_9_5_0  (
            .in0(N__44774),
            .in1(N__61581),
            .in2(N__61452),
            .in3(N__47092),
            .lcout(\ppm_encoder_1.pulses2count_9_i_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIHJ0E1_4_LC_9_5_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIHJ0E1_4_LC_9_5_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIHJ0E1_4_LC_9_5_2 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \ppm_encoder_1.throttle_RNIHJ0E1_4_LC_9_5_2  (
            .in0(N__44773),
            .in1(N__58011),
            .in2(N__42288),
            .in3(N__57157),
            .lcout(\ppm_encoder_1.un2_throttle_iv_0_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_4_LC_9_5_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_4_LC_9_5_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_4_LC_9_5_3 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.throttle_4_LC_9_5_3  (
            .in0(N__42327),
            .in1(N__42314),
            .in2(N__65299),
            .in3(N__42287),
            .lcout(\ppm_encoder_1.throttleZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87011),
            .ce(),
            .sr(N__79561));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_4_LC_9_5_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_4_LC_9_5_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_4_LC_9_5_4 .LUT_INIT=16'b0000010100000000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_4_LC_9_5_4  (
            .in0(N__42286),
            .in1(_gnd_net_),
            .in2(N__61451),
            .in3(N__61580),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_2Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_4_LC_9_5_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_4_LC_9_5_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.elevator_4_LC_9_5_5 .LUT_INIT=16'b0011101011001010;
    LogicCell40 \ppm_encoder_1.elevator_4_LC_9_5_5  (
            .in0(N__47093),
            .in1(N__44790),
            .in2(N__65298),
            .in3(N__44814),
            .lcout(\ppm_encoder_1.elevatorZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87011),
            .ce(),
            .sr(N__79561));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNIUCMN_1_LC_9_5_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNIUCMN_1_LC_9_5_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNIUCMN_1_LC_9_5_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_RNIUCMN_1_LC_9_5_6  (
            .in0(N__61430),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57158),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_RNIUCMNZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_rudder_cry_6_c_LC_9_6_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_rudder_cry_6_c_LC_9_6_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_rudder_cry_6_c_LC_9_6_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.un1_rudder_cry_6_c_LC_9_6_0  (
            .in0(_gnd_net_),
            .in1(N__42356),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_6_0_),
            .carryout(\ppm_encoder_1.un1_rudder_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_rudder_cry_6_THRU_LUT4_0_LC_9_6_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_rudder_cry_6_THRU_LUT4_0_LC_9_6_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_rudder_cry_6_THRU_LUT4_0_LC_9_6_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_rudder_cry_6_THRU_LUT4_0_LC_9_6_1  (
            .in0(_gnd_net_),
            .in1(N__44459),
            .in2(_gnd_net_),
            .in3(N__42273),
            .lcout(\ppm_encoder_1.un1_rudder_cry_6_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_rudder_cry_6 ),
            .carryout(\ppm_encoder_1.un1_rudder_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_rudder_cry_7_THRU_LUT4_0_LC_9_6_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_rudder_cry_7_THRU_LUT4_0_LC_9_6_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_rudder_cry_7_THRU_LUT4_0_LC_9_6_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_rudder_cry_7_THRU_LUT4_0_LC_9_6_2  (
            .in0(_gnd_net_),
            .in1(N__44432),
            .in2(_gnd_net_),
            .in3(N__42393),
            .lcout(\ppm_encoder_1.un1_rudder_cry_7_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_rudder_cry_7 ),
            .carryout(\ppm_encoder_1.un1_rudder_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_rudder_cry_8_THRU_LUT4_0_LC_9_6_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_rudder_cry_8_THRU_LUT4_0_LC_9_6_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_rudder_cry_8_THRU_LUT4_0_LC_9_6_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_rudder_cry_8_THRU_LUT4_0_LC_9_6_3  (
            .in0(_gnd_net_),
            .in1(N__44415),
            .in2(_gnd_net_),
            .in3(N__42390),
            .lcout(\ppm_encoder_1.un1_rudder_cry_8_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_rudder_cry_8 ),
            .carryout(\ppm_encoder_1.un1_rudder_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_rudder_cry_9_THRU_LUT4_0_LC_9_6_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_rudder_cry_9_THRU_LUT4_0_LC_9_6_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_rudder_cry_9_THRU_LUT4_0_LC_9_6_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_rudder_cry_9_THRU_LUT4_0_LC_9_6_4  (
            .in0(_gnd_net_),
            .in1(N__44510),
            .in2(_gnd_net_),
            .in3(N__42387),
            .lcout(\ppm_encoder_1.un1_rudder_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_rudder_cry_9 ),
            .carryout(\ppm_encoder_1.un1_rudder_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_rudder_cry_10_THRU_LUT4_0_LC_9_6_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_rudder_cry_10_THRU_LUT4_0_LC_9_6_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_rudder_cry_10_THRU_LUT4_0_LC_9_6_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_rudder_cry_10_THRU_LUT4_0_LC_9_6_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__44204),
            .in3(N__42384),
            .lcout(\ppm_encoder_1.un1_rudder_cry_10_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_rudder_cry_10 ),
            .carryout(\ppm_encoder_1.un1_rudder_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_rudder_cry_11_THRU_LUT4_0_LC_9_6_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_rudder_cry_11_THRU_LUT4_0_LC_9_6_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_rudder_cry_11_THRU_LUT4_0_LC_9_6_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_rudder_cry_11_THRU_LUT4_0_LC_9_6_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__44489),
            .in3(N__42381),
            .lcout(\ppm_encoder_1.un1_rudder_cry_11_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_rudder_cry_11 ),
            .carryout(\ppm_encoder_1.un1_rudder_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_rudder_cry_12_THRU_LUT4_0_LC_9_6_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_rudder_cry_12_THRU_LUT4_0_LC_9_6_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_rudder_cry_12_THRU_LUT4_0_LC_9_6_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_rudder_cry_12_THRU_LUT4_0_LC_9_6_7  (
            .in0(_gnd_net_),
            .in1(N__53708),
            .in2(N__56575),
            .in3(N__42378),
            .lcout(\ppm_encoder_1.un1_rudder_cry_12_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_rudder_cry_12 ),
            .carryout(\ppm_encoder_1.un1_rudder_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.rudder_esr_14_LC_9_7_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_esr_14_LC_9_7_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.rudder_esr_14_LC_9_7_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ppm_encoder_1.rudder_esr_14_LC_9_7_0  (
            .in0(_gnd_net_),
            .in1(N__42435),
            .in2(_gnd_net_),
            .in3(N__42375),
            .lcout(\ppm_encoder_1.rudderZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87026),
            .ce(N__50159),
            .sr(N__79569));
    defparam \scaler_4.un2_source_data_0_cry_1_c_LC_9_8_0 .C_ON=1'b1;
    defparam \scaler_4.un2_source_data_0_cry_1_c_LC_9_8_0 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un2_source_data_0_cry_1_c_LC_9_8_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \scaler_4.un2_source_data_0_cry_1_c_LC_9_8_0  (
            .in0(_gnd_net_),
            .in1(N__42663),
            .in2(N__42372),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_8_0_),
            .carryout(\scaler_4.un2_source_data_0_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.source_data_1_esr_6_LC_9_8_1 .C_ON=1'b1;
    defparam \scaler_4.source_data_1_esr_6_LC_9_8_1 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_6_LC_9_8_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.source_data_1_esr_6_LC_9_8_1  (
            .in0(_gnd_net_),
            .in1(N__42620),
            .in2(N__42673),
            .in3(N__42339),
            .lcout(scaler_4_data_6),
            .ltout(),
            .carryin(\scaler_4.un2_source_data_0_cry_1 ),
            .carryout(\scaler_4.un2_source_data_0_cry_2 ),
            .clk(N__87036),
            .ce(N__42426),
            .sr(N__79575));
    defparam \scaler_4.source_data_1_esr_7_LC_9_8_2 .C_ON=1'b1;
    defparam \scaler_4.source_data_1_esr_7_LC_9_8_2 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_7_LC_9_8_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.source_data_1_esr_7_LC_9_8_2  (
            .in0(_gnd_net_),
            .in1(N__42587),
            .in2(N__42624),
            .in3(N__42459),
            .lcout(scaler_4_data_7),
            .ltout(),
            .carryin(\scaler_4.un2_source_data_0_cry_2 ),
            .carryout(\scaler_4.un2_source_data_0_cry_3 ),
            .clk(N__87036),
            .ce(N__42426),
            .sr(N__79575));
    defparam \scaler_4.source_data_1_esr_8_LC_9_8_3 .C_ON=1'b1;
    defparam \scaler_4.source_data_1_esr_8_LC_9_8_3 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_8_LC_9_8_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.source_data_1_esr_8_LC_9_8_3  (
            .in0(_gnd_net_),
            .in1(N__42554),
            .in2(N__42591),
            .in3(N__42456),
            .lcout(scaler_4_data_8),
            .ltout(),
            .carryin(\scaler_4.un2_source_data_0_cry_3 ),
            .carryout(\scaler_4.un2_source_data_0_cry_4 ),
            .clk(N__87036),
            .ce(N__42426),
            .sr(N__79575));
    defparam \scaler_4.source_data_1_esr_9_LC_9_8_4 .C_ON=1'b1;
    defparam \scaler_4.source_data_1_esr_9_LC_9_8_4 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_9_LC_9_8_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.source_data_1_esr_9_LC_9_8_4  (
            .in0(_gnd_net_),
            .in1(N__42521),
            .in2(N__42558),
            .in3(N__42453),
            .lcout(scaler_4_data_9),
            .ltout(),
            .carryin(\scaler_4.un2_source_data_0_cry_4 ),
            .carryout(\scaler_4.un2_source_data_0_cry_5 ),
            .clk(N__87036),
            .ce(N__42426),
            .sr(N__79575));
    defparam \scaler_4.source_data_1_esr_10_LC_9_8_5 .C_ON=1'b1;
    defparam \scaler_4.source_data_1_esr_10_LC_9_8_5 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_10_LC_9_8_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.source_data_1_esr_10_LC_9_8_5  (
            .in0(_gnd_net_),
            .in1(N__42488),
            .in2(N__42525),
            .in3(N__42450),
            .lcout(scaler_4_data_10),
            .ltout(),
            .carryin(\scaler_4.un2_source_data_0_cry_5 ),
            .carryout(\scaler_4.un2_source_data_0_cry_6 ),
            .clk(N__87036),
            .ce(N__42426),
            .sr(N__79575));
    defparam \scaler_4.source_data_1_esr_11_LC_9_8_6 .C_ON=1'b1;
    defparam \scaler_4.source_data_1_esr_11_LC_9_8_6 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_11_LC_9_8_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.source_data_1_esr_11_LC_9_8_6  (
            .in0(_gnd_net_),
            .in1(N__42980),
            .in2(N__42492),
            .in3(N__42447),
            .lcout(scaler_4_data_11),
            .ltout(),
            .carryin(\scaler_4.un2_source_data_0_cry_6 ),
            .carryout(\scaler_4.un2_source_data_0_cry_7 ),
            .clk(N__87036),
            .ce(N__42426),
            .sr(N__79575));
    defparam \scaler_4.source_data_1_esr_12_LC_9_8_7 .C_ON=1'b1;
    defparam \scaler_4.source_data_1_esr_12_LC_9_8_7 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_12_LC_9_8_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.source_data_1_esr_12_LC_9_8_7  (
            .in0(_gnd_net_),
            .in1(N__42965),
            .in2(N__42984),
            .in3(N__42444),
            .lcout(scaler_4_data_12),
            .ltout(),
            .carryin(\scaler_4.un2_source_data_0_cry_7 ),
            .carryout(\scaler_4.un2_source_data_0_cry_8 ),
            .clk(N__87036),
            .ce(N__42426),
            .sr(N__79575));
    defparam \scaler_4.source_data_1_esr_13_LC_9_9_0 .C_ON=1'b1;
    defparam \scaler_4.source_data_1_esr_13_LC_9_9_0 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_13_LC_9_9_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.source_data_1_esr_13_LC_9_9_0  (
            .in0(_gnd_net_),
            .in1(N__42966),
            .in2(N__42942),
            .in3(N__42441),
            .lcout(scaler_4_data_13),
            .ltout(),
            .carryin(bfn_9_9_0_),
            .carryout(\scaler_4.un2_source_data_0_cry_9 ),
            .clk(N__87046),
            .ce(N__42421),
            .sr(N__79583));
    defparam \scaler_4.source_data_1_esr_14_LC_9_9_1 .C_ON=1'b0;
    defparam \scaler_4.source_data_1_esr_14_LC_9_9_1 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_14_LC_9_9_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \scaler_4.source_data_1_esr_14_LC_9_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42438),
            .lcout(scaler_4_data_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87046),
            .ce(N__42421),
            .sr(N__79583));
    defparam \uart_drone.bit_Count_0_LC_9_10_0 .C_ON=1'b0;
    defparam \uart_drone.bit_Count_0_LC_9_10_0 .SEQ_MODE=4'b1000;
    defparam \uart_drone.bit_Count_0_LC_9_10_0 .LUT_INIT=16'b0010011000100010;
    LogicCell40 \uart_drone.bit_Count_0_LC_9_10_0  (
            .in0(N__62053),
            .in1(N__50522),
            .in2(N__50862),
            .in3(N__44963),
            .lcout(\uart_drone.bit_CountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87056),
            .ce(),
            .sr(N__79590));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_LC_9_11_0 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_LC_9_11_0 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_LC_9_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_LC_9_11_0  (
            .in0(_gnd_net_),
            .in1(N__42747),
            .in2(N__42721),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_11_0_),
            .carryout(\scaler_4.un3_source_data_0_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_RNI40BL_LC_9_11_1 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_RNI40BL_LC_9_11_1 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_RNI40BL_LC_9_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_RNI40BL_LC_9_11_1  (
            .in0(_gnd_net_),
            .in1(N__42690),
            .in2(N__42684),
            .in3(N__42642),
            .lcout(\scaler_4.un2_source_data_0 ),
            .ltout(),
            .carryin(\scaler_4.un3_source_data_0_cry_0 ),
            .carryout(\scaler_4.un3_source_data_0_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_1_c_RNI74CL_LC_9_11_2 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_1_c_RNI74CL_LC_9_11_2 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_1_c_RNI74CL_LC_9_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_1_c_RNI74CL_LC_9_11_2  (
            .in0(_gnd_net_),
            .in1(N__42639),
            .in2(N__42633),
            .in3(N__42609),
            .lcout(\scaler_4.un3_source_data_0_cry_1_c_RNI74CL ),
            .ltout(),
            .carryin(\scaler_4.un3_source_data_0_cry_1 ),
            .carryout(\scaler_4.un3_source_data_0_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_2_c_RNIA8DL_LC_9_11_3 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_2_c_RNIA8DL_LC_9_11_3 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_2_c_RNIA8DL_LC_9_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_2_c_RNIA8DL_LC_9_11_3  (
            .in0(_gnd_net_),
            .in1(N__42606),
            .in2(N__42600),
            .in3(N__42576),
            .lcout(\scaler_4.un3_source_data_0_cry_2_c_RNIA8DL ),
            .ltout(),
            .carryin(\scaler_4.un3_source_data_0_cry_2 ),
            .carryout(\scaler_4.un3_source_data_0_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_3_c_RNIDCEL_LC_9_11_4 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_3_c_RNIDCEL_LC_9_11_4 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_3_c_RNIDCEL_LC_9_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_3_c_RNIDCEL_LC_9_11_4  (
            .in0(_gnd_net_),
            .in1(N__42573),
            .in2(N__42567),
            .in3(N__42543),
            .lcout(\scaler_4.un3_source_data_0_cry_3_c_RNIDCEL ),
            .ltout(),
            .carryin(\scaler_4.un3_source_data_0_cry_3 ),
            .carryout(\scaler_4.un3_source_data_0_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_4_c_RNIGGFL_LC_9_11_5 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_4_c_RNIGGFL_LC_9_11_5 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_4_c_RNIGGFL_LC_9_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_4_c_RNIGGFL_LC_9_11_5  (
            .in0(_gnd_net_),
            .in1(N__42540),
            .in2(N__42534),
            .in3(N__42510),
            .lcout(\scaler_4.un3_source_data_0_cry_4_c_RNIGGFL ),
            .ltout(),
            .carryin(\scaler_4.un3_source_data_0_cry_4 ),
            .carryout(\scaler_4.un3_source_data_0_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_5_c_RNIJKGL_LC_9_11_6 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_5_c_RNIJKGL_LC_9_11_6 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_5_c_RNIJKGL_LC_9_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_5_c_RNIJKGL_LC_9_11_6  (
            .in0(_gnd_net_),
            .in1(N__42507),
            .in2(N__42501),
            .in3(N__42477),
            .lcout(\scaler_4.un3_source_data_0_cry_5_c_RNIJKGL ),
            .ltout(),
            .carryin(\scaler_4.un3_source_data_0_cry_5 ),
            .carryout(\scaler_4.un3_source_data_0_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_6_c_RNIOUNN_LC_9_11_7 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_6_c_RNIOUNN_LC_9_11_7 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_6_c_RNIOUNN_LC_9_11_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_6_c_RNIOUNN_LC_9_11_7  (
            .in0(_gnd_net_),
            .in1(N__42474),
            .in2(_gnd_net_),
            .in3(N__42969),
            .lcout(\scaler_4.un3_source_data_0_cry_6_c_RNIOUNN ),
            .ltout(),
            .carryin(\scaler_4.un3_source_data_0_cry_6 ),
            .carryout(\scaler_4.un3_source_data_0_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_7_c_RNIP0PN_LC_9_12_0 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_7_c_RNIP0PN_LC_9_12_0 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_7_c_RNIP0PN_LC_9_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_7_c_RNIP0PN_LC_9_12_0  (
            .in0(_gnd_net_),
            .in1(N__53886),
            .in2(N__56550),
            .in3(N__42948),
            .lcout(\scaler_4.un3_source_data_0_cry_7_c_RNIP0PN ),
            .ltout(),
            .carryin(bfn_9_12_0_),
            .carryout(\scaler_4.un3_source_data_0_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_8_c_RNIS918_LC_9_12_1 .C_ON=1'b0;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_8_c_RNIS918_LC_9_12_1 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_8_c_RNIS918_LC_9_12_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_8_c_RNIS918_LC_9_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42945),
            .lcout(\scaler_4.un3_source_data_0_cry_8_c_RNIS918 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.WDT_RNIM3K1_4_LC_9_13_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.WDT_RNIM3K1_4_LC_9_13_0 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.WDT_RNIM3K1_4_LC_9_13_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \dron_frame_decoder_1.WDT_RNIM3K1_4_LC_9_13_0  (
            .in0(N__42930),
            .in1(N__42914),
            .in2(N__42903),
            .in3(N__42887),
            .lcout(\dron_frame_decoder_1.WDT10lto9_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.WDT_RNIA9RK1_11_LC_9_13_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.WDT_RNIA9RK1_11_LC_9_13_1 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.WDT_RNIA9RK1_11_LC_9_13_1 .LUT_INIT=16'b0000001100000111;
    LogicCell40 \dron_frame_decoder_1.WDT_RNIA9RK1_11_LC_9_13_1  (
            .in0(N__42766),
            .in1(N__42789),
            .in2(N__43065),
            .in3(N__42805),
            .lcout(),
            .ltout(\dron_frame_decoder_1.WDT10_0_i_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.WDT_RNIBUTU2_15_LC_9_13_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.WDT_RNIBUTU2_15_LC_9_13_2 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.WDT_RNIBUTU2_15_LC_9_13_2 .LUT_INIT=16'b0111001111110011;
    LogicCell40 \dron_frame_decoder_1.WDT_RNIBUTU2_15_LC_9_13_2  (
            .in0(N__42790),
            .in1(N__43045),
            .in2(N__42876),
            .in3(N__42813),
            .lcout(\dron_frame_decoder_1.WDT10_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.WDT_RNI9TKF_6_LC_9_13_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.WDT_RNI9TKF_6_LC_9_13_3 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.WDT_RNI9TKF_6_LC_9_13_3 .LUT_INIT=16'b1110000011110000;
    LogicCell40 \dron_frame_decoder_1.WDT_RNI9TKF_6_LC_9_13_3  (
            .in0(N__42857),
            .in1(N__42845),
            .in2(N__42834),
            .in3(N__42819),
            .lcout(\dron_frame_decoder_1.WDT10lt12_0 ),
            .ltout(\dron_frame_decoder_1.WDT10lt12_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.WDT_RNINA9N1_11_LC_9_13_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.WDT_RNINA9N1_11_LC_9_13_4 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.WDT_RNINA9N1_11_LC_9_13_4 .LUT_INIT=16'b1100110011001000;
    LogicCell40 \dron_frame_decoder_1.WDT_RNINA9N1_11_LC_9_13_4  (
            .in0(N__42806),
            .in1(N__42791),
            .in2(N__42771),
            .in3(N__42767),
            .lcout(),
            .ltout(\dron_frame_decoder_1.WDT10lt14_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.WDT_RNIPI9R2_15_LC_9_13_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.WDT_RNIPI9R2_15_LC_9_13_5 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.WDT_RNIPI9R2_15_LC_9_13_5 .LUT_INIT=16'b0000000000110111;
    LogicCell40 \dron_frame_decoder_1.WDT_RNIPI9R2_15_LC_9_13_5  (
            .in0(N__43063),
            .in1(N__43046),
            .in2(N__43029),
            .in3(N__50958),
            .lcout(\dron_frame_decoder_1.N_218 ),
            .ltout(\dron_frame_decoder_1.N_218_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_2_LC_9_13_6 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_2_LC_9_13_6 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.state_2_LC_9_13_6 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \dron_frame_decoder_1.state_2_LC_9_13_6  (
            .in0(N__50960),
            .in1(N__51077),
            .in2(N__43026),
            .in3(N__47823),
            .lcout(\dron_frame_decoder_1.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87088),
            .ce(),
            .sr(N__79605));
    defparam \dron_frame_decoder_1.state_RNITC181_2_LC_9_13_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNITC181_2_LC_9_13_7 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNITC181_2_LC_9_13_7 .LUT_INIT=16'b1111111101000000;
    LogicCell40 \dron_frame_decoder_1.state_RNITC181_2_LC_9_13_7  (
            .in0(N__47822),
            .in1(N__50959),
            .in2(N__51078),
            .in3(N__79965),
            .lcout(\dron_frame_decoder_1.N_700_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.source_pid_1_esr_6_LC_9_14_3 .C_ON=1'b0;
    defparam \pid_front.source_pid_1_esr_6_LC_9_14_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.source_pid_1_esr_6_LC_9_14_3 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \pid_front.source_pid_1_esr_6_LC_9_14_3  (
            .in0(N__45350),
            .in1(N__45457),
            .in2(_gnd_net_),
            .in3(N__43187),
            .lcout(front_order_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87104),
            .ce(N__45213),
            .sr(N__45180));
    defparam \pid_front.source_pid_1_esr_7_LC_9_14_4 .C_ON=1'b0;
    defparam \pid_front.source_pid_1_esr_7_LC_9_14_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.source_pid_1_esr_7_LC_9_14_4 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \pid_front.source_pid_1_esr_7_LC_9_14_4  (
            .in0(N__45455),
            .in1(N__45351),
            .in2(_gnd_net_),
            .in3(N__43158),
            .lcout(front_order_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87104),
            .ce(N__45213),
            .sr(N__45180));
    defparam \pid_front.source_pid_1_esr_9_LC_9_14_6 .C_ON=1'b0;
    defparam \pid_front.source_pid_1_esr_9_LC_9_14_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.source_pid_1_esr_9_LC_9_14_6 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \pid_front.source_pid_1_esr_9_LC_9_14_6  (
            .in0(N__45456),
            .in1(N__45352),
            .in2(_gnd_net_),
            .in3(N__43424),
            .lcout(front_order_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87104),
            .ce(N__45213),
            .sr(N__45180));
    defparam \pid_front.pid_prereg_esr_RNIN7IV_28_LC_9_14_7 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_esr_RNIN7IV_28_LC_9_14_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_esr_RNIN7IV_28_LC_9_14_7 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \pid_front.pid_prereg_esr_RNIN7IV_28_LC_9_14_7  (
            .in0(N__45349),
            .in1(N__43593),
            .in2(_gnd_net_),
            .in3(N__43620),
            .lcout(\pid_front.un11lto30_i_a2_6_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_esr_RNIDDR99_30_LC_9_15_1 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_esr_RNIDDR99_30_LC_9_15_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_esr_RNIDDR99_30_LC_9_15_1 .LUT_INIT=16'b1111111110101011;
    LogicCell40 \pid_front.pid_prereg_esr_RNIDDR99_30_LC_9_15_1  (
            .in0(N__43095),
            .in1(N__45697),
            .in2(N__45379),
            .in3(N__43005),
            .lcout(),
            .ltout(\pid_front.N_102_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.state_RNIH9GOH_1_LC_9_15_2 .C_ON=1'b0;
    defparam \pid_front.state_RNIH9GOH_1_LC_9_15_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.state_RNIH9GOH_1_LC_9_15_2 .LUT_INIT=16'b1111111110001010;
    LogicCell40 \pid_front.state_RNIH9GOH_1_LC_9_15_2  (
            .in0(N__60112),
            .in1(N__42999),
            .in2(N__42990),
            .in3(N__66038),
            .lcout(\pid_front.un1_reset_0_i ),
            .ltout(\pid_front.un1_reset_0_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.state_RNIEI7TH_1_LC_9_15_3 .C_ON=1'b0;
    defparam \pid_front.state_RNIEI7TH_1_LC_9_15_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.state_RNIEI7TH_1_LC_9_15_3 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \pid_front.state_RNIEI7TH_1_LC_9_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__42987),
            .in3(N__60113),
            .lcout(\pid_front.state_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.source_pid_1_esr_4_LC_9_15_4 .C_ON=1'b0;
    defparam \pid_front.source_pid_1_esr_4_LC_9_15_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.source_pid_1_esr_4_LC_9_15_4 .LUT_INIT=16'b1111111111001101;
    LogicCell40 \pid_front.source_pid_1_esr_4_LC_9_15_4  (
            .in0(N__45378),
            .in1(N__43098),
            .in2(N__45462),
            .in3(N__43257),
            .lcout(front_order_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87119),
            .ce(N__45211),
            .sr(N__45167));
    defparam \pid_front.source_pid_1_esr_5_LC_9_15_5 .C_ON=1'b0;
    defparam \pid_front.source_pid_1_esr_5_LC_9_15_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.source_pid_1_esr_5_LC_9_15_5 .LUT_INIT=16'b1010001010100000;
    LogicCell40 \pid_front.source_pid_1_esr_5_LC_9_15_5  (
            .in0(N__43223),
            .in1(N__43131),
            .in2(N__45381),
            .in3(N__45453),
            .lcout(front_order_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87119),
            .ce(N__45211),
            .sr(N__45167));
    defparam \pid_front.source_pid_1_esr_0_LC_9_15_6 .C_ON=1'b0;
    defparam \pid_front.source_pid_1_esr_0_LC_9_15_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.source_pid_1_esr_0_LC_9_15_6 .LUT_INIT=16'b0011001000000000;
    LogicCell40 \pid_front.source_pid_1_esr_0_LC_9_15_6  (
            .in0(N__45377),
            .in1(N__43096),
            .in2(N__45461),
            .in3(N__43341),
            .lcout(front_order_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87119),
            .ce(N__45211),
            .sr(N__45167));
    defparam \pid_front.source_pid_1_esr_1_LC_9_15_7 .C_ON=1'b0;
    defparam \pid_front.source_pid_1_esr_1_LC_9_15_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.source_pid_1_esr_1_LC_9_15_7 .LUT_INIT=16'b0101010000000000;
    LogicCell40 \pid_front.source_pid_1_esr_1_LC_9_15_7  (
            .in0(N__43097),
            .in1(N__45454),
            .in2(N__45380),
            .in3(N__43317),
            .lcout(front_order_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87119),
            .ce(N__45211),
            .sr(N__45167));
    defparam \pid_front.pid_prereg_esr_RNIVFPG_1_LC_9_16_2 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_esr_RNIVFPG_1_LC_9_16_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_esr_RNIVFPG_1_LC_9_16_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_front.pid_prereg_esr_RNIVFPG_1_LC_9_16_2  (
            .in0(N__43313),
            .in1(N__43216),
            .in2(N__43281),
            .in3(N__43295),
            .lcout(\pid_front.source_pid_1_sqmuxa_1_0_a4_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un11lto30_i_a2_0_c_RNO_LC_9_16_3 .C_ON=1'b0;
    defparam \pid_front.un11lto30_i_a2_0_c_RNO_LC_9_16_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.un11lto30_i_a2_0_c_RNO_LC_9_16_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_front.un11lto30_i_a2_0_c_RNO_LC_9_16_3  (
            .in0(N__43294),
            .in1(N__43312),
            .in2(N__43280),
            .in3(N__43336),
            .lcout(\pid_front.source_pid10lt4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.source_pid_1_esr_2_LC_9_16_4 .C_ON=1'b0;
    defparam \pid_front.source_pid_1_esr_2_LC_9_16_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.source_pid_1_esr_2_LC_9_16_4 .LUT_INIT=16'b0011001000000000;
    LogicCell40 \pid_front.source_pid_1_esr_2_LC_9_16_4  (
            .in0(N__45365),
            .in1(N__43093),
            .in2(N__45459),
            .in3(N__43296),
            .lcout(front_order_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87134),
            .ce(N__45214),
            .sr(N__45176));
    defparam \pid_front.source_pid_1_esr_3_LC_9_16_6 .C_ON=1'b0;
    defparam \pid_front.source_pid_1_esr_3_LC_9_16_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.source_pid_1_esr_3_LC_9_16_6 .LUT_INIT=16'b0011001000000000;
    LogicCell40 \pid_front.source_pid_1_esr_3_LC_9_16_6  (
            .in0(N__45366),
            .in1(N__43094),
            .in2(N__45460),
            .in3(N__43276),
            .lcout(front_order_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87134),
            .ce(N__45214),
            .sr(N__45176));
    defparam \pid_front.un1_pid_prereg_0_cry_0_c_THRU_CRY_0_LC_9_17_0 .C_ON=1'b1;
    defparam \pid_front.un1_pid_prereg_0_cry_0_c_THRU_CRY_0_LC_9_17_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.un1_pid_prereg_0_cry_0_c_THRU_CRY_0_LC_9_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_front.un1_pid_prereg_0_cry_0_c_THRU_CRY_0_LC_9_17_0  (
            .in0(_gnd_net_),
            .in1(N__49547),
            .in2(N__49551),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_17_0_),
            .carryout(\pid_front.un1_pid_prereg_0_cry_0_c_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_esr_0_LC_9_17_1 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_0_LC_9_17_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_0_LC_9_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_0_LC_9_17_1  (
            .in0(_gnd_net_),
            .in1(N__49791),
            .in2(N__54849),
            .in3(N__43320),
            .lcout(\pid_front.pid_preregZ0Z_0 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_0_cry_0_c_THRU_CO ),
            .carryout(\pid_front.un1_pid_prereg_0_cry_0 ),
            .clk(N__87153),
            .ce(N__56087),
            .sr(N__79633));
    defparam \pid_front.pid_prereg_esr_1_LC_9_17_2 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_1_LC_9_17_2 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_1_LC_9_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_1_LC_9_17_2  (
            .in0(_gnd_net_),
            .in1(N__49827),
            .in2(N__54813),
            .in3(N__43299),
            .lcout(\pid_front.pid_preregZ0Z_1 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_0_cry_0 ),
            .carryout(\pid_front.un1_pid_prereg_0_cry_1 ),
            .clk(N__87153),
            .ce(N__56087),
            .sr(N__79633));
    defparam \pid_front.pid_prereg_esr_2_LC_9_17_3 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_2_LC_9_17_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_2_LC_9_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_2_LC_9_17_3  (
            .in0(_gnd_net_),
            .in1(N__52347),
            .in2(N__54765),
            .in3(N__43284),
            .lcout(\pid_front.pid_preregZ0Z_2 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_0_cry_1 ),
            .carryout(\pid_front.un1_pid_prereg_0_cry_2 ),
            .clk(N__87153),
            .ce(N__56087),
            .sr(N__79633));
    defparam \pid_front.pid_prereg_esr_3_LC_9_17_4 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_3_LC_9_17_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_3_LC_9_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_3_LC_9_17_4  (
            .in0(_gnd_net_),
            .in1(N__52304),
            .in2(N__51396),
            .in3(N__43260),
            .lcout(\pid_front.pid_preregZ0Z_3 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_0_cry_2 ),
            .carryout(\pid_front.un1_pid_prereg_0_cry_3 ),
            .clk(N__87153),
            .ce(N__56087),
            .sr(N__79633));
    defparam \pid_front.pid_prereg_esr_4_LC_9_17_5 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_4_LC_9_17_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_4_LC_9_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_4_LC_9_17_5  (
            .in0(_gnd_net_),
            .in1(N__45126),
            .in2(N__51371),
            .in3(N__43227),
            .lcout(\pid_front.pid_preregZ0Z_4 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_0_cry_3 ),
            .carryout(\pid_front.un1_pid_prereg_0_cry_4 ),
            .clk(N__87153),
            .ce(N__56087),
            .sr(N__79633));
    defparam \pid_front.pid_prereg_esr_5_LC_9_17_6 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_5_LC_9_17_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_5_LC_9_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_5_LC_9_17_6  (
            .in0(_gnd_net_),
            .in1(N__45800),
            .in2(N__45810),
            .in3(N__43191),
            .lcout(\pid_front.pid_preregZ0Z_5 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_0_cry_4 ),
            .carryout(\pid_front.un1_pid_prereg_0_cry_5 ),
            .clk(N__87153),
            .ce(N__56087),
            .sr(N__79633));
    defparam \pid_front.pid_prereg_esr_6_LC_9_17_7 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_6_LC_9_17_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_6_LC_9_17_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_6_LC_9_17_7  (
            .in0(_gnd_net_),
            .in1(N__45729),
            .in2(N__45756),
            .in3(N__43161),
            .lcout(\pid_front.pid_preregZ0Z_6 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_0_cry_5 ),
            .carryout(\pid_front.un1_pid_prereg_0_cry_6 ),
            .clk(N__87153),
            .ce(N__56087),
            .sr(N__79633));
    defparam \pid_front.pid_prereg_esr_7_LC_9_18_0 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_7_LC_9_18_0 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_7_LC_9_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_7_LC_9_18_0  (
            .in0(_gnd_net_),
            .in1(N__46191),
            .in2(N__45927),
            .in3(N__43137),
            .lcout(\pid_front.pid_preregZ0Z_7 ),
            .ltout(),
            .carryin(bfn_9_18_0_),
            .carryout(\pid_front.un1_pid_prereg_0_cry_7 ),
            .clk(N__87168),
            .ce(N__56086),
            .sr(N__79640));
    defparam \pid_front.pid_prereg_esr_8_LC_9_18_1 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_8_LC_9_18_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_8_LC_9_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_8_LC_9_18_1  (
            .in0(_gnd_net_),
            .in1(N__48141),
            .in2(N__48167),
            .in3(N__43134),
            .lcout(\pid_front.pid_preregZ0Z_8 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_0_cry_7 ),
            .carryout(\pid_front.un1_pid_prereg_0_cry_8 ),
            .clk(N__87168),
            .ce(N__56086),
            .sr(N__79640));
    defparam \pid_front.pid_prereg_esr_9_LC_9_18_2 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_9_LC_9_18_2 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_9_LC_9_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_9_LC_9_18_2  (
            .in0(_gnd_net_),
            .in1(N__43431),
            .in2(N__47798),
            .in3(N__43398),
            .lcout(\pid_front.pid_preregZ0Z_9 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_0_cry_8 ),
            .carryout(\pid_front.un1_pid_prereg_0_cry_9 ),
            .clk(N__87168),
            .ce(N__56086),
            .sr(N__79640));
    defparam \pid_front.pid_prereg_esr_10_LC_9_18_3 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_10_LC_9_18_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_10_LC_9_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_10_LC_9_18_3  (
            .in0(_gnd_net_),
            .in1(N__45825),
            .in2(N__46023),
            .in3(N__43395),
            .lcout(\pid_front.pid_preregZ0Z_10 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_0_cry_9 ),
            .carryout(\pid_front.un1_pid_prereg_0_cry_10 ),
            .clk(N__87168),
            .ce(N__56086),
            .sr(N__79640));
    defparam \pid_front.pid_prereg_esr_11_LC_9_18_4 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_11_LC_9_18_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_11_LC_9_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_11_LC_9_18_4  (
            .in0(_gnd_net_),
            .in1(N__46754),
            .in2(N__46065),
            .in3(N__43392),
            .lcout(\pid_front.pid_preregZ0Z_11 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_0_cry_10 ),
            .carryout(\pid_front.un1_pid_prereg_0_cry_11 ),
            .clk(N__87168),
            .ce(N__56086),
            .sr(N__79640));
    defparam \pid_front.pid_prereg_esr_12_LC_9_18_5 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_12_LC_9_18_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_12_LC_9_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_12_LC_9_18_5  (
            .in0(_gnd_net_),
            .in1(N__43854),
            .in2(N__46716),
            .in3(N__43389),
            .lcout(\pid_front.pid_preregZ0Z_12 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_0_cry_11 ),
            .carryout(\pid_front.un1_pid_prereg_0_cry_12 ),
            .clk(N__87168),
            .ce(N__56086),
            .sr(N__79640));
    defparam \pid_front.pid_prereg_esr_13_LC_9_18_6 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_13_LC_9_18_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_13_LC_9_18_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_13_LC_9_18_6  (
            .in0(_gnd_net_),
            .in1(N__51878),
            .in2(N__43710),
            .in3(N__43386),
            .lcout(\pid_front.pid_preregZ0Z_13 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_0_cry_12 ),
            .carryout(\pid_front.un1_pid_prereg_0_cry_13 ),
            .clk(N__87168),
            .ce(N__56086),
            .sr(N__79640));
    defparam \pid_front.un1_pid_prereg_0_cry_13_THRU_LUT4_0_LC_9_18_7 .C_ON=1'b1;
    defparam \pid_front.un1_pid_prereg_0_cry_13_THRU_LUT4_0_LC_9_18_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.un1_pid_prereg_0_cry_13_THRU_LUT4_0_LC_9_18_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.un1_pid_prereg_0_cry_13_THRU_LUT4_0_LC_9_18_7  (
            .in0(_gnd_net_),
            .in1(N__48695),
            .in2(_gnd_net_),
            .in3(N__43377),
            .lcout(\pid_front.un1_pid_prereg_0_cry_13_THRU_CO ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_0_cry_13 ),
            .carryout(\pid_front.un1_pid_prereg_0_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_esr_15_LC_9_19_0 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_15_LC_9_19_0 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_15_LC_9_19_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_15_LC_9_19_0  (
            .in0(_gnd_net_),
            .in1(N__46400),
            .in2(N__46362),
            .in3(N__43356),
            .lcout(\pid_front.pid_preregZ0Z_15 ),
            .ltout(),
            .carryin(bfn_9_19_0_),
            .carryout(\pid_front.un1_pid_prereg_0_cry_15 ),
            .clk(N__87182),
            .ce(N__56085),
            .sr(N__79648));
    defparam \pid_front.pid_prereg_esr_16_LC_9_19_1 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_16_LC_9_19_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_16_LC_9_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_16_LC_9_19_1  (
            .in0(_gnd_net_),
            .in1(N__43821),
            .in2(N__43809),
            .in3(N__43344),
            .lcout(\pid_front.pid_preregZ0Z_16 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_0_cry_15 ),
            .carryout(\pid_front.un1_pid_prereg_0_cry_16 ),
            .clk(N__87182),
            .ce(N__56085),
            .sr(N__79648));
    defparam \pid_front.pid_prereg_esr_17_LC_9_19_2 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_17_LC_9_19_2 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_17_LC_9_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_17_LC_9_19_2  (
            .in0(_gnd_net_),
            .in1(N__44037),
            .in2(N__43794),
            .in3(N__43542),
            .lcout(\pid_front.pid_preregZ0Z_17 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_0_cry_16 ),
            .carryout(\pid_front.un1_pid_prereg_0_cry_17 ),
            .clk(N__87182),
            .ce(N__56085),
            .sr(N__79648));
    defparam \pid_front.pid_prereg_esr_18_LC_9_19_3 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_18_LC_9_19_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_18_LC_9_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_18_LC_9_19_3  (
            .in0(_gnd_net_),
            .in1(N__43986),
            .in2(N__44022),
            .in3(N__43530),
            .lcout(\pid_front.pid_preregZ0Z_18 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_0_cry_17 ),
            .carryout(\pid_front.un1_pid_prereg_0_cry_18 ),
            .clk(N__87182),
            .ce(N__56085),
            .sr(N__79648));
    defparam \pid_front.pid_prereg_esr_19_LC_9_19_4 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_19_LC_9_19_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_19_LC_9_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_19_LC_9_19_4  (
            .in0(_gnd_net_),
            .in1(N__51777),
            .in2(N__43974),
            .in3(N__43518),
            .lcout(\pid_front.pid_preregZ0Z_19 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_0_cry_18 ),
            .carryout(\pid_front.un1_pid_prereg_0_cry_19 ),
            .clk(N__87182),
            .ce(N__56085),
            .sr(N__79648));
    defparam \pid_front.pid_prereg_esr_20_LC_9_19_5 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_20_LC_9_19_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_20_LC_9_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_20_LC_9_19_5  (
            .in0(_gnd_net_),
            .in1(N__43515),
            .in2(N__51951),
            .in3(N__43503),
            .lcout(\pid_front.pid_preregZ0Z_20 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_0_cry_19 ),
            .carryout(\pid_front.un1_pid_prereg_0_cry_20 ),
            .clk(N__87182),
            .ce(N__56085),
            .sr(N__79648));
    defparam \pid_front.pid_prereg_esr_21_LC_9_19_6 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_21_LC_9_19_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_21_LC_9_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_21_LC_9_19_6  (
            .in0(_gnd_net_),
            .in1(N__43500),
            .in2(N__43494),
            .in3(N__43479),
            .lcout(\pid_front.pid_preregZ0Z_21 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_0_cry_20 ),
            .carryout(\pid_front.un1_pid_prereg_0_cry_21 ),
            .clk(N__87182),
            .ce(N__56085),
            .sr(N__79648));
    defparam \pid_front.pid_prereg_esr_22_LC_9_19_7 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_22_LC_9_19_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_22_LC_9_19_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_22_LC_9_19_7  (
            .in0(_gnd_net_),
            .in1(N__45960),
            .in2(N__43476),
            .in3(N__43461),
            .lcout(\pid_front.pid_preregZ0Z_22 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_0_cry_21 ),
            .carryout(\pid_front.un1_pid_prereg_0_cry_22 ),
            .clk(N__87182),
            .ce(N__56085),
            .sr(N__79648));
    defparam \pid_front.pid_prereg_esr_23_LC_9_20_0 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_23_LC_9_20_0 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_23_LC_9_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_23_LC_9_20_0  (
            .in0(_gnd_net_),
            .in1(N__46137),
            .in2(N__46110),
            .in3(N__43446),
            .lcout(\pid_front.pid_preregZ0Z_23 ),
            .ltout(),
            .carryin(bfn_9_20_0_),
            .carryout(\pid_front.un1_pid_prereg_0_cry_23 ),
            .clk(N__87196),
            .ce(N__56083),
            .sr(N__79656));
    defparam \pid_front.pid_prereg_esr_24_LC_9_20_1 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_24_LC_9_20_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_24_LC_9_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_24_LC_9_20_1  (
            .in0(_gnd_net_),
            .in1(N__43752),
            .in2(N__46005),
            .in3(N__43434),
            .lcout(\pid_front.pid_preregZ0Z_24 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_0_cry_23 ),
            .carryout(\pid_front.un1_pid_prereg_0_cry_24 ),
            .clk(N__87196),
            .ce(N__56083),
            .sr(N__79656));
    defparam \pid_front.pid_prereg_esr_25_LC_9_20_2 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_25_LC_9_20_2 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_25_LC_9_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_25_LC_9_20_2  (
            .in0(_gnd_net_),
            .in1(N__43773),
            .in2(N__43566),
            .in3(N__43686),
            .lcout(\pid_front.pid_preregZ0Z_25 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_0_cry_24 ),
            .carryout(\pid_front.un1_pid_prereg_0_cry_25 ),
            .clk(N__87196),
            .ce(N__56083),
            .sr(N__79656));
    defparam \pid_front.pid_prereg_esr_26_LC_9_20_3 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_26_LC_9_20_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_26_LC_9_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_26_LC_9_20_3  (
            .in0(_gnd_net_),
            .in1(N__43683),
            .in2(N__43719),
            .in3(N__43668),
            .lcout(\pid_front.pid_preregZ0Z_26 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_0_cry_25 ),
            .carryout(\pid_front.un1_pid_prereg_0_cry_26 ),
            .clk(N__87196),
            .ce(N__56083),
            .sr(N__79656));
    defparam \pid_front.pid_prereg_esr_27_LC_9_20_4 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_27_LC_9_20_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_27_LC_9_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_27_LC_9_20_4  (
            .in0(_gnd_net_),
            .in1(N__43665),
            .in2(N__43659),
            .in3(N__43638),
            .lcout(\pid_front.pid_preregZ0Z_27 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_0_cry_26 ),
            .carryout(\pid_front.un1_pid_prereg_0_cry_27 ),
            .clk(N__87196),
            .ce(N__56083),
            .sr(N__79656));
    defparam \pid_front.pid_prereg_esr_28_LC_9_20_5 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_28_LC_9_20_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_28_LC_9_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_28_LC_9_20_5  (
            .in0(_gnd_net_),
            .in1(N__43635),
            .in2(N__43629),
            .in3(N__43611),
            .lcout(\pid_front.pid_preregZ0Z_28 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_0_cry_27 ),
            .carryout(\pid_front.un1_pid_prereg_0_cry_28 ),
            .clk(N__87196),
            .ce(N__56083),
            .sr(N__79656));
    defparam \pid_front.pid_prereg_esr_29_LC_9_20_6 .C_ON=1'b1;
    defparam \pid_front.pid_prereg_esr_29_LC_9_20_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_29_LC_9_20_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.pid_prereg_esr_29_LC_9_20_6  (
            .in0(_gnd_net_),
            .in1(N__43608),
            .in2(N__43602),
            .in3(N__43581),
            .lcout(\pid_front.pid_preregZ0Z_29 ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_0_cry_28 ),
            .carryout(\pid_front.un1_pid_prereg_0_cry_29 ),
            .clk(N__87196),
            .ce(N__56083),
            .sr(N__79656));
    defparam \pid_front.pid_prereg_esr_30_LC_9_20_7 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_esr_30_LC_9_20_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_30_LC_9_20_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_front.pid_prereg_esr_30_LC_9_20_7  (
            .in0(_gnd_net_),
            .in1(N__43578),
            .in2(_gnd_net_),
            .in3(N__43572),
            .lcout(\pid_front.pid_preregZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87196),
            .ce(N__56083),
            .sr(N__79656));
    defparam \pid_front.error_d_reg_prev_esr_RNIJGV52_0_22_LC_9_21_0 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIJGV52_0_22_LC_9_21_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIJGV52_0_22_LC_9_21_0 .LUT_INIT=16'b0001100011100111;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIJGV52_0_22_LC_9_21_0  (
            .in0(N__87414),
            .in1(N__48337),
            .in2(N__46331),
            .in3(N__55664),
            .lcout(\pid_front.un1_pid_prereg_0_17 ),
            .ltout(\pid_front.un1_pid_prereg_0_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNI4UTB4_22_LC_9_21_1 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNI4UTB4_22_LC_9_21_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNI4UTB4_22_LC_9_21_1 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNI4UTB4_22_LC_9_21_1  (
            .in0(N__46250),
            .in1(_gnd_net_),
            .in2(N__43569),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_d_reg_prev_esr_RNI4UTB4Z0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIJGV52_22_LC_9_21_2 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIJGV52_22_LC_9_21_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIJGV52_22_LC_9_21_2 .LUT_INIT=16'b1110111100001000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIJGV52_22_LC_9_21_2  (
            .in0(N__87415),
            .in1(N__48338),
            .in2(N__46332),
            .in3(N__55665),
            .lcout(\pid_front.un1_pid_prereg_0_18 ),
            .ltout(\pid_front.un1_pid_prereg_0_18_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIC2UN8_22_LC_9_21_3 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIC2UN8_22_LC_9_21_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIC2UN8_22_LC_9_21_3 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIC2UN8_22_LC_9_21_3  (
            .in0(N__46251),
            .in1(N__43767),
            .in2(N__43776),
            .in3(N__43745),
            .lcout(\pid_front.error_d_reg_prev_esr_RNIC2UN8Z0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIFJ8U9_22_LC_9_21_4 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIFJ8U9_22_LC_9_21_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIFJ8U9_22_LC_9_21_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIFJ8U9_22_LC_9_21_4  (
            .in0(N__45954),
            .in1(N__46249),
            .in2(N__46155),
            .in3(N__43763),
            .lcout(\pid_front.error_d_reg_prev_esr_RNIFJ8U9Z0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIVTNC2_0_14_LC_9_21_5 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIVTNC2_0_14_LC_9_21_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIVTNC2_0_14_LC_9_21_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \pid_front.error_p_reg_esr_RNIVTNC2_0_14_LC_9_21_5  (
            .in0(N__54303),
            .in1(N__82776),
            .in2(N__54269),
            .in3(N__46161),
            .lcout(\pid_front.g0_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNILJ062_0_22_LC_9_21_6 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNILJ062_0_22_LC_9_21_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNILJ062_0_22_LC_9_21_6 .LUT_INIT=16'b0001100011100111;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNILJ062_0_22_LC_9_21_6  (
            .in0(N__87416),
            .in1(N__48339),
            .in2(N__46333),
            .in3(N__56291),
            .lcout(\pid_front.un1_pid_prereg_0_19 ),
            .ltout(\pid_front.un1_pid_prereg_0_19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNI840C4_22_LC_9_21_7 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNI840C4_22_LC_9_21_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNI840C4_22_LC_9_21_7 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNI840C4_22_LC_9_21_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__43734),
            .in3(N__43730),
            .lcout(\pid_front.error_d_reg_prev_esr_RNI840C4Z0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI1IK9E_12_LC_9_22_0 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI1IK9E_12_LC_9_22_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI1IK9E_12_LC_9_22_0 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_front.error_p_reg_esr_RNI1IK9E_12_LC_9_22_0  (
            .in0(N__54933),
            .in1(N__43830),
            .in2(N__51885),
            .in3(N__43911),
            .lcout(\pid_front.error_p_reg_esr_RNI1IK9EZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNILTVH2_0_12_LC_9_22_1 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNILTVH2_0_12_LC_9_22_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNILTVH2_0_12_LC_9_22_1 .LUT_INIT=16'b0101000001110001;
    LogicCell40 \pid_front.error_p_reg_esr_RNILTVH2_0_12_LC_9_22_1  (
            .in0(N__48969),
            .in1(N__48907),
            .in2(N__43842),
            .in3(N__49247),
            .lcout(),
            .ltout(\pid_front.un1_pid_prereg_167_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNI1KIM4_12_LC_9_22_2 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNI1KIM4_12_LC_9_22_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNI1KIM4_12_LC_9_22_2 .LUT_INIT=16'b1010111100100011;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNI1KIM4_12_LC_9_22_2  (
            .in0(N__51915),
            .in1(N__48671),
            .in2(N__43698),
            .in3(N__49625),
            .lcout(\pid_front.un1_pid_prereg_167_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIK2AG3_12_LC_9_22_3 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIK2AG3_12_LC_9_22_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIK2AG3_12_LC_9_22_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \pid_front.error_p_reg_esr_RNIK2AG3_12_LC_9_22_3  (
            .in0(N__43829),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54932),
            .lcout(),
            .ltout(\pid_front.un1_pid_prereg_153_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIHM5CD_10_LC_9_22_4 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIHM5CD_10_LC_9_22_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIHM5CD_10_LC_9_22_4 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIHM5CD_10_LC_9_22_4  (
            .in0(N__54972),
            .in1(N__46737),
            .in2(N__43857),
            .in3(N__43910),
            .lcout(\pid_front.error_d_reg_prev_esr_RNIHM5CDZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_fast_esr_RNIOTBC_0_12_LC_9_22_5 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_fast_esr_RNIOTBC_0_12_LC_9_22_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_fast_esr_RNIOTBC_0_12_LC_9_22_5 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \pid_front.error_d_reg_fast_esr_RNIOTBC_0_12_LC_9_22_5  (
            .in0(N__46583),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48528),
            .lcout(\pid_front.N_2191_i ),
            .ltout(\pid_front.N_2191_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNILTVH2_12_LC_9_22_6 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNILTVH2_12_LC_9_22_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNILTVH2_12_LC_9_22_6 .LUT_INIT=16'b0001111011100001;
    LogicCell40 \pid_front.error_p_reg_esr_RNILTVH2_12_LC_9_22_6  (
            .in0(N__49248),
            .in1(N__48908),
            .in2(N__43833),
            .in3(N__48970),
            .lcout(\pid_front.error_p_reg_esr_RNILTVH2Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIJVCRE_13_LC_9_22_7 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIJVCRE_13_LC_9_22_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIJVCRE_13_LC_9_22_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \pid_front.error_p_reg_esr_RNIJVCRE_13_LC_9_22_7  (
            .in0(N__46378),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46415),
            .lcout(\pid_front.error_p_reg_esr_RNIJVCREZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIHFPHL_13_LC_9_23_0 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIHFPHL_13_LC_9_23_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIHFPHL_13_LC_9_23_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_front.error_p_reg_esr_RNIHFPHL_13_LC_9_23_0  (
            .in0(N__46422),
            .in1(N__44068),
            .in2(N__46386),
            .in3(N__44048),
            .lcout(\pid_front.error_p_reg_esr_RNIHFPHLZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIJS6B3_0_15_LC_9_23_1 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIJS6B3_0_15_LC_9_23_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIJS6B3_0_15_LC_9_23_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_front.error_p_reg_esr_RNIJS6B3_0_15_LC_9_23_1  (
            .in0(N__43947),
            .in1(N__43959),
            .in2(_gnd_net_),
            .in3(N__55350),
            .lcout(\pid_front.un1_pid_prereg_0_1 ),
            .ltout(\pid_front.un1_pid_prereg_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIUFCM6_14_LC_9_23_2 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIUFCM6_14_LC_9_23_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIUFCM6_14_LC_9_23_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \pid_front.error_p_reg_esr_RNIUFCM6_14_LC_9_23_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__43797),
            .in3(N__44069),
            .lcout(\pid_front.error_p_reg_esr_RNIUFCM6Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIH0C61_14_LC_9_23_3 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIH0C61_14_LC_9_23_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIH0C61_14_LC_9_23_3 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_front.error_p_reg_esr_RNIH0C61_14_LC_9_23_3  (
            .in0(N__54255),
            .in1(N__54302),
            .in2(_gnd_net_),
            .in3(N__82770),
            .lcout(\pid_front.error_p_reg_esr_RNIH0C61Z0Z_14 ),
            .ltout(\pid_front.error_p_reg_esr_RNIH0C61Z0Z_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIBJ5B3_0_14_LC_9_23_4 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIBJ5B3_0_14_LC_9_23_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIBJ5B3_0_14_LC_9_23_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_p_reg_esr_RNIBJ5B3_0_14_LC_9_23_4  (
            .in0(_gnd_net_),
            .in1(N__43898),
            .in2(N__43779),
            .in3(N__55378),
            .lcout(\pid_front.error_p_reg_esr_RNIBJ5B3_0Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIBJ5B3_14_LC_9_23_5 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIBJ5B3_14_LC_9_23_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIBJ5B3_14_LC_9_23_5 .LUT_INIT=16'b1111101010100000;
    LogicCell40 \pid_front.error_p_reg_esr_RNIBJ5B3_14_LC_9_23_5  (
            .in0(N__55379),
            .in1(_gnd_net_),
            .in2(N__43902),
            .in3(N__43917),
            .lcout(\pid_front.un1_pid_prereg_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNI5JRF4_10_LC_9_23_7 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNI5JRF4_10_LC_9_23_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNI5JRF4_10_LC_9_23_7 .LUT_INIT=16'b1111110111000100;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNI5JRF4_10_LC_9_23_7  (
            .in0(N__46533),
            .in1(N__46460),
            .in2(N__46500),
            .in3(N__46539),
            .lcout(\pid_front.error_d_reg_prev_esr_RNI5JRF4Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIETB61_4_13_LC_9_24_0 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIETB61_4_13_LC_9_24_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIETB61_4_13_LC_9_24_0 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_front.error_p_reg_esr_RNIETB61_4_13_LC_9_24_0  (
            .in0(N__48885),
            .in1(N__48795),
            .in2(_gnd_net_),
            .in3(N__48767),
            .lcout(\pid_front.error_p_reg_esr_RNIETB61_4Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_13_LC_9_24_1 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_13_LC_9_24_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_13_LC_9_24_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_front.error_d_reg_prev_esr_13_LC_9_24_1  (
            .in0(N__48768),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_d_reg_prevZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87252),
            .ce(N__70490),
            .sr(N__70348));
    defparam \pid_front.error_p_reg_esr_RNIK3C61_0_15_LC_9_24_2 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIK3C61_0_15_LC_9_24_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIK3C61_0_15_LC_9_24_2 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_front.error_p_reg_esr_RNIK3C61_0_15_LC_9_24_2  (
            .in0(N__43889),
            .in1(N__43865),
            .in2(_gnd_net_),
            .in3(N__87322),
            .lcout(\pid_front.error_p_reg_esr_RNIK3C61_0Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_15_LC_9_24_3 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_15_LC_9_24_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_15_LC_9_24_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_front.error_d_reg_prev_esr_15_LC_9_24_3  (
            .in0(N__87324),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_d_reg_prevZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87252),
            .ce(N__70490),
            .sr(N__70348));
    defparam \pid_front.error_p_reg_esr_RNIK3C61_15_LC_9_24_4 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIK3C61_15_LC_9_24_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIK3C61_15_LC_9_24_4 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_front.error_p_reg_esr_RNIK3C61_15_LC_9_24_4  (
            .in0(N__43890),
            .in1(N__43866),
            .in2(_gnd_net_),
            .in3(N__87323),
            .lcout(\pid_front.error_p_reg_esr_RNIK3C61Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIN6C61_0_16_LC_9_24_5 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIN6C61_0_16_LC_9_24_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIN6C61_0_16_LC_9_24_5 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_front.error_p_reg_esr_RNIN6C61_0_16_LC_9_24_5  (
            .in0(N__44105),
            .in1(N__44081),
            .in2(_gnd_net_),
            .in3(N__87295),
            .lcout(\pid_front.error_p_reg_esr_RNIN6C61_0Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_16_LC_9_24_6 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_16_LC_9_24_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_16_LC_9_24_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_front.error_d_reg_prev_esr_16_LC_9_24_6  (
            .in0(N__87297),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_d_reg_prevZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87252),
            .ce(N__70490),
            .sr(N__70348));
    defparam \pid_front.error_p_reg_esr_RNIN6C61_16_LC_9_24_7 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIN6C61_16_LC_9_24_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIN6C61_16_LC_9_24_7 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_front.error_p_reg_esr_RNIN6C61_16_LC_9_24_7  (
            .in0(N__44106),
            .in1(N__44082),
            .in2(_gnd_net_),
            .in3(N__87296),
            .lcout(\pid_front.error_p_reg_esr_RNIN6C61Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNICIRCD_14_LC_9_25_0 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNICIRCD_14_LC_9_25_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNICIRCD_14_LC_9_25_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_front.error_p_reg_esr_RNICIRCD_14_LC_9_25_0  (
            .in0(N__44073),
            .in1(N__43997),
            .in2(N__44055),
            .in3(N__43931),
            .lcout(\pid_front.error_p_reg_esr_RNICIRCDZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIR58B3_0_16_LC_9_25_1 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIR58B3_0_16_LC_9_25_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIR58B3_0_16_LC_9_25_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_front.error_p_reg_esr_RNIR58B3_0_16_LC_9_25_1  (
            .in0(N__51737),
            .in1(N__44006),
            .in2(_gnd_net_),
            .in3(N__56173),
            .lcout(\pid_front.un1_pid_prereg_0_3 ),
            .ltout(\pid_front.un1_pid_prereg_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIE2FM6_15_LC_9_25_2 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIE2FM6_15_LC_9_25_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIE2FM6_15_LC_9_25_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \pid_front.error_p_reg_esr_RNIE2FM6_15_LC_9_25_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__44025),
            .in3(N__43930),
            .lcout(\pid_front.error_p_reg_esr_RNIE2FM6Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIR58B3_16_LC_9_25_3 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIR58B3_16_LC_9_25_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIR58B3_16_LC_9_25_3 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_front.error_p_reg_esr_RNIR58B3_16_LC_9_25_3  (
            .in0(N__51738),
            .in1(N__44007),
            .in2(_gnd_net_),
            .in3(N__56174),
            .lcout(\pid_front.un1_pid_prereg_0_4 ),
            .ltout(\pid_front.un1_pid_prereg_0_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNICN0DD_15_LC_9_25_4 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNICN0DD_15_LC_9_25_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNICN0DD_15_LC_9_25_4 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \pid_front.error_p_reg_esr_RNICN0DD_15_LC_9_25_4  (
            .in0(N__43932),
            .in1(N__43998),
            .in2(N__43989),
            .in3(N__51791),
            .lcout(\pid_front.error_p_reg_esr_RNICN0DDZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI3F9B3_0_17_LC_9_25_5 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI3F9B3_0_17_LC_9_25_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI3F9B3_0_17_LC_9_25_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_front.error_p_reg_esr_RNI3F9B3_0_17_LC_9_25_5  (
            .in0(N__51843),
            .in1(N__51864),
            .in2(_gnd_net_),
            .in3(N__55312),
            .lcout(\pid_front.un1_pid_prereg_0_5 ),
            .ltout(\pid_front.un1_pid_prereg_0_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIUKHM6_16_LC_9_25_6 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIUKHM6_16_LC_9_25_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIUKHM6_16_LC_9_25_6 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \pid_front.error_p_reg_esr_RNIUKHM6_16_LC_9_25_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__43977),
            .in3(N__51812),
            .lcout(\pid_front.error_p_reg_esr_RNIUKHM6Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIJS6B3_15_LC_9_25_7 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIJS6B3_15_LC_9_25_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIJS6B3_15_LC_9_25_7 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_front.error_p_reg_esr_RNIJS6B3_15_LC_9_25_7  (
            .in0(N__43958),
            .in1(N__55346),
            .in2(_gnd_net_),
            .in3(N__43943),
            .lcout(\pid_front.un1_pid_prereg_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIC9HV_12_LC_10_1_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIC9HV_12_LC_10_1_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIC9HV_12_LC_10_1_0 .LUT_INIT=16'b1111000001111000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIC9HV_12_LC_10_1_0  (
            .in0(N__60940),
            .in1(N__61015),
            .in2(N__50436),
            .in3(N__64257),
            .lcout(\ppm_encoder_1.N_267_i_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIUKK21_5_LC_10_1_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIUKK21_5_LC_10_1_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIUKK21_5_LC_10_1_1 .LUT_INIT=16'b1001110011001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIUKK21_5_LC_10_1_1  (
            .in0(N__64258),
            .in1(N__59662),
            .in2(N__61042),
            .in3(N__60941),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_5_LC_10_1_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_5_LC_10_1_2 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_5_LC_10_1_2 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \ppm_encoder_1.init_pulses_5_LC_10_1_2  (
            .in0(N__55808),
            .in1(N__46782),
            .in2(N__55951),
            .in3(N__44298),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__86974),
            .ce(),
            .sr(N__79556));
    defparam \ppm_encoder_1.init_pulses_12_LC_10_1_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_12_LC_10_1_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.init_pulses_12_LC_10_1_3 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \ppm_encoder_1.init_pulses_12_LC_10_1_3  (
            .in0(N__55806),
            .in1(N__46860),
            .in2(N__55952),
            .in3(N__44217),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__86974),
            .ce(),
            .sr(N__79556));
    defparam \ppm_encoder_1.init_pulses_RNID4MT_11_LC_10_1_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNID4MT_11_LC_10_1_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNID4MT_11_LC_10_1_5 .LUT_INIT=16'b1011010011110000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNID4MT_11_LC_10_1_5  (
            .in0(N__64259),
            .in1(N__64586),
            .in2(N__53055),
            .in3(N__63430),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIG7MT_14_LC_10_1_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIG7MT_14_LC_10_1_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIG7MT_14_LC_10_1_6 .LUT_INIT=16'b1100110001101100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIG7MT_14_LC_10_1_6  (
            .in0(N__63431),
            .in1(N__57493),
            .in2(N__64601),
            .in3(N__64260),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_14_LC_10_1_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_14_LC_10_1_7 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_14_LC_10_1_7 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \ppm_encoder_1.init_pulses_14_LC_10_1_7  (
            .in0(N__55807),
            .in1(N__46842),
            .in2(N__55953),
            .in3(N__44367),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__86974),
            .ce(),
            .sr(N__79556));
    defparam \ppm_encoder_1.init_pulses_3_LC_10_2_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_3_LC_10_2_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.init_pulses_3_LC_10_2_0 .LUT_INIT=16'b0010001100100000;
    LogicCell40 \ppm_encoder_1.init_pulses_3_LC_10_2_0  (
            .in0(N__46806),
            .in1(N__55783),
            .in2(N__55936),
            .in3(N__44145),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__86977),
            .ce(),
            .sr(N__79559));
    defparam \ppm_encoder_1.init_pulses_4_LC_10_2_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_4_LC_10_2_1 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_4_LC_10_2_1 .LUT_INIT=16'b0000101100001000;
    LogicCell40 \ppm_encoder_1.init_pulses_4_LC_10_2_1  (
            .in0(N__46797),
            .in1(N__55894),
            .in2(N__55804),
            .in3(N__44115),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__86977),
            .ce(),
            .sr(N__79559));
    defparam \ppm_encoder_1.init_pulses_6_LC_10_2_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_6_LC_10_2_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.init_pulses_6_LC_10_2_2 .LUT_INIT=16'b0010001100100000;
    LogicCell40 \ppm_encoder_1.init_pulses_6_LC_10_2_2  (
            .in0(N__46773),
            .in1(N__55787),
            .in2(N__55937),
            .in3(N__44286),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__86977),
            .ce(),
            .sr(N__79559));
    defparam \ppm_encoder_1.init_pulses_7_LC_10_2_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_7_LC_10_2_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.init_pulses_7_LC_10_2_3 .LUT_INIT=16'b0000101100001000;
    LogicCell40 \ppm_encoder_1.init_pulses_7_LC_10_2_3  (
            .in0(N__46911),
            .in1(N__55895),
            .in2(N__55805),
            .in3(N__44277),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__86977),
            .ce(),
            .sr(N__79559));
    defparam \ppm_encoder_1.init_pulses_8_LC_10_2_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_8_LC_10_2_4 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_8_LC_10_2_4 .LUT_INIT=16'b0010001100100000;
    LogicCell40 \ppm_encoder_1.init_pulses_8_LC_10_2_4  (
            .in0(N__46890),
            .in1(N__55791),
            .in2(N__55938),
            .in3(N__44247),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__86977),
            .ce(),
            .sr(N__79559));
    defparam \ppm_encoder_1.init_pulses_11_LC_10_2_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_11_LC_10_2_5 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_11_LC_10_2_5 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \ppm_encoder_1.init_pulses_11_LC_10_2_5  (
            .in0(N__55782),
            .in1(N__46869),
            .in2(N__55939),
            .in3(N__44229),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__86977),
            .ce(),
            .sr(N__79559));
    defparam \ppm_encoder_1.rudder_11_LC_10_2_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_11_LC_10_2_7 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.rudder_11_LC_10_2_7 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.rudder_11_LC_10_2_7  (
            .in0(N__44205),
            .in1(N__44184),
            .in2(N__65306),
            .in3(N__53611),
            .lcout(\ppm_encoder_1.rudderZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__86977),
            .ce(),
            .sr(N__79559));
    defparam \ppm_encoder_1.init_pulses_RNIN39V4_0_LC_10_3_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNIN39V4_0_LC_10_3_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIN39V4_0_LC_10_3_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIN39V4_0_LC_10_3_0  (
            .in0(_gnd_net_),
            .in1(N__53190),
            .in2(N__53978),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_10_3_0_),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_1_LC_10_3_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_1_LC_10_3_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_1_LC_10_3_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_1_LC_10_3_1  (
            .in0(_gnd_net_),
            .in1(N__56730),
            .in2(N__56745),
            .in3(N__44172),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_1 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_0 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_2_LC_10_3_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_2_LC_10_3_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_2_LC_10_3_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_2_LC_10_3_2  (
            .in0(_gnd_net_),
            .in1(N__57723),
            .in2(N__57648),
            .in3(N__44169),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_2 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_1 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_3_LC_10_3_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_3_LC_10_3_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_3_LC_10_3_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_3_LC_10_3_3  (
            .in0(_gnd_net_),
            .in1(N__44166),
            .in2(N__44160),
            .in3(N__44139),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_3 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_2 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_4_LC_10_3_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_4_LC_10_3_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_4_LC_10_3_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_4_LC_10_3_4  (
            .in0(_gnd_net_),
            .in1(N__44136),
            .in2(N__44130),
            .in3(N__44109),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_4 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_3 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_5_LC_10_3_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_5_LC_10_3_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_5_LC_10_3_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_5_LC_10_3_5  (
            .in0(_gnd_net_),
            .in1(N__44319),
            .in2(N__44313),
            .in3(N__44289),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_5 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_4 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_6_LC_10_3_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_6_LC_10_3_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_6_LC_10_3_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_6_LC_10_3_6  (
            .in0(_gnd_net_),
            .in1(N__50208),
            .in2(N__50241),
            .in3(N__44280),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_6 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_5 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_7_LC_10_3_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_7_LC_10_3_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_7_LC_10_3_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_7_LC_10_3_7  (
            .in0(_gnd_net_),
            .in1(N__53463),
            .in2(N__53487),
            .in3(N__44271),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_7 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_6 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_8_LC_10_4_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_8_LC_10_4_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_8_LC_10_4_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_8_LC_10_4_0  (
            .in0(_gnd_net_),
            .in1(N__44268),
            .in2(N__44262),
            .in3(N__44238),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_8 ),
            .ltout(),
            .carryin(bfn_10_4_0_),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_9_LC_10_4_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_9_LC_10_4_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_9_LC_10_4_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_9_LC_10_4_1  (
            .in0(_gnd_net_),
            .in1(N__46971),
            .in2(N__47139),
            .in3(N__44235),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_9 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_8 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_10_LC_10_4_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_10_LC_10_4_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_10_LC_10_4_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_10_LC_10_4_2  (
            .in0(_gnd_net_),
            .in1(N__50082),
            .in2(N__50370),
            .in3(N__44232),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_10 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_9 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_11_LC_10_4_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_11_LC_10_4_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_11_LC_10_4_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_11_LC_10_4_3  (
            .in0(_gnd_net_),
            .in1(N__53076),
            .in2(N__53025),
            .in3(N__44220),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_11 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_10 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_12_LC_10_4_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_12_LC_10_4_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_12_LC_10_4_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_12_LC_10_4_4  (
            .in0(_gnd_net_),
            .in1(N__47295),
            .in2(N__47316),
            .in3(N__44208),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_12 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_11 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_13_LC_10_4_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_13_LC_10_4_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_13_LC_10_4_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_13_LC_10_4_5  (
            .in0(_gnd_net_),
            .in1(N__53415),
            .in2(N__53448),
            .in3(N__44370),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_13 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_12 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_14_LC_10_4_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_14_LC_10_4_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_14_LC_10_4_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_14_LC_10_4_6  (
            .in0(_gnd_net_),
            .in1(N__53304),
            .in2(N__53292),
            .in3(N__44355),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_14 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_13 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_15_LC_10_4_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_15_LC_10_4_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_15_LC_10_4_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_15_LC_10_4_7  (
            .in0(_gnd_net_),
            .in1(N__50022),
            .in2(N__50040),
            .in3(N__44352),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_15 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_14 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_16_LC_10_5_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_16_LC_10_5_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_16_LC_10_5_0 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_16_LC_10_5_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__44340),
            .in3(N__44349),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_16 ),
            .ltout(),
            .carryin(bfn_10_5_0_),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_17_LC_10_5_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_17_LC_10_5_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_17_LC_10_5_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_17_LC_10_5_1  (
            .in0(_gnd_net_),
            .in1(N__44331),
            .in2(_gnd_net_),
            .in3(N__44346),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_17 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_16 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_18_LC_10_5_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNO_0_18_LC_10_5_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_18_LC_10_5_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_18_LC_10_5_2  (
            .in0(_gnd_net_),
            .in1(N__60601),
            .in2(_gnd_net_),
            .in3(N__44343),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNII9MT_0_16_LC_10_5_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNII9MT_0_16_LC_10_5_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNII9MT_0_16_LC_10_5_3 .LUT_INIT=16'b1100110001101100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNII9MT_0_16_LC_10_5_3  (
            .in0(N__64590),
            .in1(N__63928),
            .in2(N__63456),
            .in3(N__64287),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIJAMT_0_17_LC_10_5_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIJAMT_0_17_LC_10_5_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIJAMT_0_17_LC_10_5_6 .LUT_INIT=16'b1001110011001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIJAMT_0_17_LC_10_5_6  (
            .in0(N__64286),
            .in1(N__64618),
            .in2(N__63457),
            .in3(N__64591),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_axb_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIFH0E1_3_LC_10_5_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIFH0E1_3_LC_10_5_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIFH0E1_3_LC_10_5_7 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \ppm_encoder_1.throttle_RNIFH0E1_3_LC_10_5_7  (
            .in0(N__57994),
            .in1(N__68171),
            .in2(N__68595),
            .in3(N__57156),
            .lcout(\ppm_encoder_1.un2_throttle_iv_0_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_5_LC_10_6_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_5_LC_10_6_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.aileron_5_LC_10_6_0 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \ppm_encoder_1.aileron_5_LC_10_6_0  (
            .in0(N__47337),
            .in1(N__53535),
            .in2(N__44551),
            .in3(N__65277),
            .lcout(\ppm_encoder_1.aileronZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87005),
            .ce(),
            .sr(N__79566));
    defparam \ppm_encoder_1.rudder_10_LC_10_6_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_10_LC_10_6_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.rudder_10_LC_10_6_2 .LUT_INIT=16'b0111101101001000;
    LogicCell40 \ppm_encoder_1.rudder_10_LC_10_6_2  (
            .in0(N__44520),
            .in1(N__65278),
            .in2(N__44514),
            .in3(N__60790),
            .lcout(\ppm_encoder_1.rudderZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87005),
            .ce(),
            .sr(N__79566));
    defparam \ppm_encoder_1.aileron_10_LC_10_6_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_10_LC_10_6_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.aileron_10_LC_10_6_3 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.aileron_10_LC_10_6_3  (
            .in0(N__53793),
            .in1(N__47490),
            .in2(N__65304),
            .in3(N__56803),
            .lcout(\ppm_encoder_1.aileronZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87005),
            .ce(),
            .sr(N__79566));
    defparam \ppm_encoder_1.rudder_12_LC_10_6_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_12_LC_10_6_4 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.rudder_12_LC_10_6_4 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \ppm_encoder_1.rudder_12_LC_10_6_4  (
            .in0(N__44496),
            .in1(N__44490),
            .in2(N__50483),
            .in3(N__65279),
            .lcout(\ppm_encoder_1.rudderZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87005),
            .ce(),
            .sr(N__79566));
    defparam \ppm_encoder_1.rudder_7_LC_10_6_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_7_LC_10_6_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.rudder_7_LC_10_6_5 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.rudder_7_LC_10_6_5  (
            .in0(N__44466),
            .in1(N__44460),
            .in2(N__65305),
            .in3(N__57862),
            .lcout(\ppm_encoder_1.rudderZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87005),
            .ce(),
            .sr(N__79566));
    defparam \ppm_encoder_1.rudder_8_LC_10_6_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_8_LC_10_6_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.rudder_8_LC_10_6_6 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \ppm_encoder_1.rudder_8_LC_10_6_6  (
            .in0(N__44442),
            .in1(N__44436),
            .in2(N__60682),
            .in3(N__65283),
            .lcout(\ppm_encoder_1.rudderZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87005),
            .ce(),
            .sr(N__79566));
    defparam \ppm_encoder_1.rudder_9_LC_10_7_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_9_LC_10_7_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.rudder_9_LC_10_7_0 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.rudder_9_LC_10_7_0  (
            .in0(N__44414),
            .in1(N__44400),
            .in2(N__65265),
            .in3(N__61795),
            .lcout(\ppm_encoder_1.rudderZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87013),
            .ce(),
            .sr(N__79570));
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNIJMMD_LC_10_7_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNIJMMD_LC_10_7_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNIJMMD_LC_10_7_1 .LUT_INIT=16'b0111011101110111;
    LogicCell40 \ppm_encoder_1.counter24_0_I_57_c_RNIJMMD_LC_10_7_1  (
            .in0(N__61162),
            .in1(N__61109),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\ppm_encoder_1.counter24_0_I_57_c_RNIJMMDZ0 ),
            .ltout(\ppm_encoder_1.counter24_0_I_57_c_RNIJMMDZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.ppm_output_reg_LC_10_7_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.ppm_output_reg_LC_10_7_2 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.ppm_output_reg_LC_10_7_2 .LUT_INIT=16'b1000101110101011;
    LogicCell40 \ppm_encoder_1.ppm_output_reg_LC_10_7_2  (
            .in0(N__44381),
            .in1(N__60513),
            .in2(N__44394),
            .in3(N__61218),
            .lcout(ppm_output_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87013),
            .ce(),
            .sr(N__79570));
    defparam \ppm_encoder_1.throttle_10_LC_10_7_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_10_LC_10_7_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_10_LC_10_7_3 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \ppm_encoder_1.throttle_10_LC_10_7_3  (
            .in0(N__44673),
            .in1(N__44661),
            .in2(N__60757),
            .in3(N__65172),
            .lcout(\ppm_encoder_1.throttleZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87013),
            .ce(),
            .sr(N__79570));
    defparam \ppm_encoder_1.throttle_13_LC_10_7_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_13_LC_10_7_5 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.throttle_13_LC_10_7_5 .LUT_INIT=16'b1001100111110000;
    LogicCell40 \ppm_encoder_1.throttle_13_LC_10_7_5  (
            .in0(N__44625),
            .in1(N__44598),
            .in2(N__61486),
            .in3(N__65173),
            .lcout(\ppm_encoder_1.throttleZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87013),
            .ce(),
            .sr(N__79570));
    defparam \ppm_encoder_1.throttle_2_LC_10_7_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_2_LC_10_7_6 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.throttle_2_LC_10_7_6 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.throttle_2_LC_10_7_6  (
            .in0(N__44586),
            .in1(N__44574),
            .in2(N__65266),
            .in3(N__53332),
            .lcout(\ppm_encoder_1.throttleZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87013),
            .ce(),
            .sr(N__79570));
    defparam \ppm_encoder_1.aileron_2_LC_10_8_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_2_LC_10_8_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.aileron_2_LC_10_8_0 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.aileron_2_LC_10_8_0  (
            .in0(N__47358),
            .in1(N__58181),
            .in2(N__65284),
            .in3(N__68836),
            .lcout(\ppm_encoder_1.aileronZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87020),
            .ce(),
            .sr(N__79576));
    defparam \ppm_encoder_1.elevator_11_LC_10_8_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_11_LC_10_8_1 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.elevator_11_LC_10_8_1 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \ppm_encoder_1.elevator_11_LC_10_8_1  (
            .in0(N__45477),
            .in1(N__45012),
            .in2(N__52630),
            .in3(N__65213),
            .lcout(\ppm_encoder_1.elevatorZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87020),
            .ce(),
            .sr(N__79576));
    defparam \ppm_encoder_1.elevator_3_LC_10_8_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_3_LC_10_8_2 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.elevator_3_LC_10_8_2 .LUT_INIT=16'b1001111110010000;
    LogicCell40 \ppm_encoder_1.elevator_3_LC_10_8_2  (
            .in0(N__44826),
            .in1(N__44853),
            .in2(N__65286),
            .in3(N__52852),
            .lcout(\ppm_encoder_1.elevatorZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87020),
            .ce(),
            .sr(N__79576));
    defparam \ppm_encoder_1.elevator_1_LC_10_8_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_1_LC_10_8_3 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.elevator_1_LC_10_8_3 .LUT_INIT=16'b1110001000101110;
    LogicCell40 \ppm_encoder_1.elevator_1_LC_10_8_3  (
            .in0(N__58028),
            .in1(N__65217),
            .in2(N__44922),
            .in3(N__44898),
            .lcout(\ppm_encoder_1.elevatorZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87020),
            .ce(),
            .sr(N__79576));
    defparam \ppm_encoder_1.elevator_12_LC_10_8_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_12_LC_10_8_4 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.elevator_12_LC_10_8_4 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.elevator_12_LC_10_8_4  (
            .in0(N__45567),
            .in1(N__45000),
            .in2(N__65285),
            .in3(N__47285),
            .lcout(\ppm_encoder_1.elevatorZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87020),
            .ce(),
            .sr(N__79576));
    defparam \ppm_encoder_1.elevator_2_LC_10_8_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_2_LC_10_8_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.elevator_2_LC_10_8_6 .LUT_INIT=16'b0111001011011000;
    LogicCell40 \ppm_encoder_1.elevator_2_LC_10_8_6  (
            .in0(N__65218),
            .in1(N__44886),
            .in2(N__58060),
            .in3(N__44865),
            .lcout(\ppm_encoder_1.elevatorZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87020),
            .ce(),
            .sr(N__79576));
    defparam \ppm_encoder_1.elevator_8_LC_10_9_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_8_LC_10_9_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.elevator_8_LC_10_9_0 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.elevator_8_LC_10_9_0  (
            .in0(N__45519),
            .in1(N__45066),
            .in2(N__65288),
            .in3(N__47159),
            .lcout(\ppm_encoder_1.elevatorZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87028),
            .ce(),
            .sr(N__79584));
    defparam \ppm_encoder_1.aileron_4_LC_10_9_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_4_LC_10_9_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.aileron_4_LC_10_9_1 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \ppm_encoder_1.aileron_4_LC_10_9_1  (
            .in0(N__47346),
            .in1(N__53768),
            .in2(N__44775),
            .in3(N__65222),
            .lcout(\ppm_encoder_1.aileronZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87028),
            .ce(),
            .sr(N__79584));
    defparam \ppm_encoder_1.elevator_9_LC_10_9_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_9_LC_10_9_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.elevator_9_LC_10_9_2 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.elevator_9_LC_10_9_2  (
            .in0(N__45036),
            .in1(N__45054),
            .in2(N__65289),
            .in3(N__47383),
            .lcout(\ppm_encoder_1.elevatorZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87028),
            .ce(),
            .sr(N__79584));
    defparam \ppm_encoder_1.aileron_9_LC_10_9_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_9_LC_10_9_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.aileron_9_LC_10_9_5 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \ppm_encoder_1.aileron_9_LC_10_9_5  (
            .in0(N__53730),
            .in1(N__47499),
            .in2(N__47414),
            .in3(N__65223),
            .lcout(\ppm_encoder_1.aileronZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87028),
            .ce(),
            .sr(N__79584));
    defparam \ppm_encoder_1.elevator_13_LC_10_9_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_13_LC_10_9_6 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.elevator_13_LC_10_9_6 .LUT_INIT=16'b1001111110010000;
    LogicCell40 \ppm_encoder_1.elevator_13_LC_10_9_6  (
            .in0(N__45720),
            .in1(N__44988),
            .in2(N__65287),
            .in3(N__50498),
            .lcout(\ppm_encoder_1.elevatorZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87028),
            .ce(),
            .sr(N__79584));
    defparam \ppm_encoder_1.elevator_10_LC_10_9_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_10_LC_10_9_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.elevator_10_LC_10_9_7 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \ppm_encoder_1.elevator_10_LC_10_9_7  (
            .in0(N__45024),
            .in1(N__45240),
            .in2(N__56779),
            .in3(N__65224),
            .lcout(\ppm_encoder_1.elevatorZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87028),
            .ce(),
            .sr(N__79584));
    defparam \uart_drone.state_RNO_0_3_LC_10_10_0 .C_ON=1'b0;
    defparam \uart_drone.state_RNO_0_3_LC_10_10_0 .SEQ_MODE=4'b0000;
    defparam \uart_drone.state_RNO_0_3_LC_10_10_0 .LUT_INIT=16'b0001001100110011;
    LogicCell40 \uart_drone.state_RNO_0_3_LC_10_10_0  (
            .in0(N__50786),
            .in1(N__44954),
            .in2(N__44751),
            .in3(N__50834),
            .lcout(),
            .ltout(\uart_drone.N_145_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_3_LC_10_10_1 .C_ON=1'b0;
    defparam \uart_drone.state_3_LC_10_10_1 .SEQ_MODE=4'b1000;
    defparam \uart_drone.state_3_LC_10_10_1 .LUT_INIT=16'b0000000000001011;
    LogicCell40 \uart_drone.state_3_LC_10_10_1  (
            .in0(N__44750),
            .in1(N__50717),
            .in2(N__44715),
            .in3(N__79991),
            .lcout(\uart_drone.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87038),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_RNI62411_4_LC_10_10_3 .C_ON=1'b0;
    defparam \uart_drone.state_RNI62411_4_LC_10_10_3 .SEQ_MODE=4'b0000;
    defparam \uart_drone.state_RNI62411_4_LC_10_10_3 .LUT_INIT=16'b0010001100000011;
    LogicCell40 \uart_drone.state_RNI62411_4_LC_10_10_3  (
            .in0(N__50833),
            .in1(N__44710),
            .in2(N__44964),
            .in3(N__50785),
            .lcout(\uart_drone.un1_state_4_0 ),
            .ltout(\uart_drone.un1_state_4_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.bit_Count_RNO_0_2_LC_10_10_4 .C_ON=1'b0;
    defparam \uart_drone.bit_Count_RNO_0_2_LC_10_10_4 .SEQ_MODE=4'b0000;
    defparam \uart_drone.bit_Count_RNO_0_2_LC_10_10_4 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \uart_drone.bit_Count_RNO_0_2_LC_10_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__44676),
            .in3(N__62046),
            .lcout(\uart_drone.CO0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.data_Aux_RNO_0_3_LC_10_10_5 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_RNO_0_3_LC_10_10_5 .SEQ_MODE=4'b0000;
    defparam \uart_drone.data_Aux_RNO_0_3_LC_10_10_5 .LUT_INIT=16'b0000100000001000;
    LogicCell40 \uart_drone.data_Aux_RNO_0_3_LC_10_10_5  (
            .in0(N__62047),
            .in1(N__62132),
            .in2(N__62204),
            .in3(_gnd_net_),
            .lcout(\uart_drone.data_Auxce_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.bit_Count_RNIJOJC1_2_LC_10_10_6 .C_ON=1'b0;
    defparam \uart_drone.bit_Count_RNIJOJC1_2_LC_10_10_6 .SEQ_MODE=4'b0000;
    defparam \uart_drone.bit_Count_RNIJOJC1_2_LC_10_10_6 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uart_drone.bit_Count_RNIJOJC1_2_LC_10_10_6  (
            .in0(N__62131),
            .in1(N__62186),
            .in2(_gnd_net_),
            .in3(N__62045),
            .lcout(\uart_drone.N_152 ),
            .ltout(\uart_drone.N_152_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_RNI63LK2_3_LC_10_10_7 .C_ON=1'b0;
    defparam \uart_drone.state_RNI63LK2_3_LC_10_10_7 .SEQ_MODE=4'b0000;
    defparam \uart_drone.state_RNI63LK2_3_LC_10_10_7 .LUT_INIT=16'b1111010100000000;
    LogicCell40 \uart_drone.state_RNI63LK2_3_LC_10_10_7  (
            .in0(N__44953),
            .in1(_gnd_net_),
            .in2(N__44925),
            .in3(N__50521),
            .lcout(\uart_drone.un1_state_7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_0_c_LC_10_11_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_0_c_LC_10_11_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_0_c_LC_10_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_0_c_LC_10_11_0  (
            .in0(_gnd_net_),
            .in1(N__53105),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_10_11_0_),
            .carryout(\ppm_encoder_1.un1_elevator_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_0_THRU_LUT4_0_LC_10_11_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_0_THRU_LUT4_0_LC_10_11_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_0_THRU_LUT4_0_LC_10_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_0_THRU_LUT4_0_LC_10_11_1  (
            .in0(_gnd_net_),
            .in1(N__44915),
            .in2(N__56547),
            .in3(N__44889),
            .lcout(\ppm_encoder_1.un1_elevator_cry_0_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_0 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_1_THRU_LUT4_0_LC_10_11_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_1_THRU_LUT4_0_LC_10_11_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_1_THRU_LUT4_0_LC_10_11_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_1_THRU_LUT4_0_LC_10_11_2  (
            .in0(_gnd_net_),
            .in1(N__44882),
            .in2(_gnd_net_),
            .in3(N__44856),
            .lcout(\ppm_encoder_1.un1_elevator_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_1 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_2_THRU_LUT4_0_LC_10_11_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_2_THRU_LUT4_0_LC_10_11_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_2_THRU_LUT4_0_LC_10_11_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_2_THRU_LUT4_0_LC_10_11_3  (
            .in0(_gnd_net_),
            .in1(N__44849),
            .in2(N__56548),
            .in3(N__44817),
            .lcout(\ppm_encoder_1.un1_elevator_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_2 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_3_THRU_LUT4_0_LC_10_11_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_3_THRU_LUT4_0_LC_10_11_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_3_THRU_LUT4_0_LC_10_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_3_THRU_LUT4_0_LC_10_11_4  (
            .in0(_gnd_net_),
            .in1(N__44813),
            .in2(_gnd_net_),
            .in3(N__44778),
            .lcout(\ppm_encoder_1.un1_elevator_cry_3_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_3 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_4_THRU_LUT4_0_LC_10_11_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_4_THRU_LUT4_0_LC_10_11_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_4_THRU_LUT4_0_LC_10_11_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_4_THRU_LUT4_0_LC_10_11_5  (
            .in0(_gnd_net_),
            .in1(N__45110),
            .in2(_gnd_net_),
            .in3(N__45075),
            .lcout(\ppm_encoder_1.un1_elevator_cry_4_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_4 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_5_THRU_LUT4_0_LC_10_11_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_5_THRU_LUT4_0_LC_10_11_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_5_THRU_LUT4_0_LC_10_11_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_5_THRU_LUT4_0_LC_10_11_6  (
            .in0(_gnd_net_),
            .in1(N__50573),
            .in2(N__56549),
            .in3(N__45072),
            .lcout(\ppm_encoder_1.un1_elevator_cry_5_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_5 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_6_THRU_LUT4_0_LC_10_11_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_6_THRU_LUT4_0_LC_10_11_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_6_THRU_LUT4_0_LC_10_11_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_6_THRU_LUT4_0_LC_10_11_7  (
            .in0(_gnd_net_),
            .in1(N__50276),
            .in2(_gnd_net_),
            .in3(N__45069),
            .lcout(\ppm_encoder_1.un1_elevator_cry_6_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_6 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_7_THRU_LUT4_0_LC_10_12_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_7_THRU_LUT4_0_LC_10_12_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_7_THRU_LUT4_0_LC_10_12_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_7_THRU_LUT4_0_LC_10_12_0  (
            .in0(_gnd_net_),
            .in1(N__45518),
            .in2(_gnd_net_),
            .in3(N__45057),
            .lcout(\ppm_encoder_1.un1_elevator_cry_7_THRU_CO ),
            .ltout(),
            .carryin(bfn_10_12_0_),
            .carryout(\ppm_encoder_1.un1_elevator_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_8_THRU_LUT4_0_LC_10_12_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_8_THRU_LUT4_0_LC_10_12_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_8_THRU_LUT4_0_LC_10_12_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_8_THRU_LUT4_0_LC_10_12_1  (
            .in0(_gnd_net_),
            .in1(N__45050),
            .in2(_gnd_net_),
            .in3(N__45027),
            .lcout(\ppm_encoder_1.un1_elevator_cry_8_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_8 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_9_THRU_LUT4_0_LC_10_12_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_9_THRU_LUT4_0_LC_10_12_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_9_THRU_LUT4_0_LC_10_12_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_9_THRU_LUT4_0_LC_10_12_2  (
            .in0(_gnd_net_),
            .in1(N__45236),
            .in2(_gnd_net_),
            .in3(N__45015),
            .lcout(\ppm_encoder_1.un1_elevator_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_9 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_10_THRU_LUT4_0_LC_10_12_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_10_THRU_LUT4_0_LC_10_12_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_10_THRU_LUT4_0_LC_10_12_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_10_THRU_LUT4_0_LC_10_12_3  (
            .in0(_gnd_net_),
            .in1(N__45476),
            .in2(_gnd_net_),
            .in3(N__45003),
            .lcout(\ppm_encoder_1.un1_elevator_cry_10_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_10 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_11_THRU_LUT4_0_LC_10_12_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_11_THRU_LUT4_0_LC_10_12_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_11_THRU_LUT4_0_LC_10_12_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_11_THRU_LUT4_0_LC_10_12_4  (
            .in0(_gnd_net_),
            .in1(N__45563),
            .in2(_gnd_net_),
            .in3(N__44991),
            .lcout(\ppm_encoder_1.un1_elevator_cry_11_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_11 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_12_THRU_LUT4_0_LC_10_12_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_12_THRU_LUT4_0_LC_10_12_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_12_THRU_LUT4_0_LC_10_12_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_12_THRU_LUT4_0_LC_10_12_5  (
            .in0(_gnd_net_),
            .in1(N__45713),
            .in2(N__56551),
            .in3(N__44979),
            .lcout(\ppm_encoder_1.un1_elevator_cry_12_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_12 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_esr_14_LC_10_12_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_esr_14_LC_10_12_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.elevator_esr_14_LC_10_12_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.elevator_esr_14_LC_10_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45723),
            .lcout(\ppm_encoder_1.elevatorZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87058),
            .ce(N__50153),
            .sr(N__79601));
    defparam \pid_front.source_pid_1_esr_13_LC_10_13_1 .C_ON=1'b0;
    defparam \pid_front.source_pid_1_esr_13_LC_10_13_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.source_pid_1_esr_13_LC_10_13_1 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \pid_front.source_pid_1_esr_13_LC_10_13_1  (
            .in0(N__45382),
            .in1(N__45702),
            .in2(_gnd_net_),
            .in3(N__45656),
            .lcout(front_order_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87065),
            .ce(N__45222),
            .sr(N__45168));
    defparam \pid_front.source_pid_1_esr_12_LC_10_14_2 .C_ON=1'b0;
    defparam \pid_front.source_pid_1_esr_12_LC_10_14_2 .SEQ_MODE=4'b1000;
    defparam \pid_front.source_pid_1_esr_12_LC_10_14_2 .LUT_INIT=16'b1111000000100000;
    LogicCell40 \pid_front.source_pid_1_esr_12_LC_10_14_2  (
            .in0(N__45698),
            .in1(N__45657),
            .in2(N__45609),
            .in3(N__45374),
            .lcout(front_order_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87077),
            .ce(N__45215),
            .sr(N__45169));
    defparam \pid_front.source_pid_1_esr_8_LC_10_14_4 .C_ON=1'b0;
    defparam \pid_front.source_pid_1_esr_8_LC_10_14_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.source_pid_1_esr_8_LC_10_14_4 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \pid_front.source_pid_1_esr_8_LC_10_14_4  (
            .in0(N__45458),
            .in1(N__45373),
            .in2(_gnd_net_),
            .in3(N__45549),
            .lcout(front_order_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87077),
            .ce(N__45215),
            .sr(N__45169));
    defparam \pid_front.source_pid_1_esr_11_LC_10_15_4 .C_ON=1'b0;
    defparam \pid_front.source_pid_1_esr_11_LC_10_15_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.source_pid_1_esr_11_LC_10_15_4 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \pid_front.source_pid_1_esr_11_LC_10_15_4  (
            .in0(N__45375),
            .in1(N__45446),
            .in2(_gnd_net_),
            .in3(N__45501),
            .lcout(front_order_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87090),
            .ce(N__45212),
            .sr(N__45166));
    defparam \pid_front.source_pid_1_esr_10_LC_10_15_7 .C_ON=1'b0;
    defparam \pid_front.source_pid_1_esr_10_LC_10_15_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.source_pid_1_esr_10_LC_10_15_7 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \pid_front.source_pid_1_esr_10_LC_10_15_7  (
            .in0(N__45445),
            .in1(N__45376),
            .in2(_gnd_net_),
            .in3(N__45258),
            .lcout(front_order_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87090),
            .ce(N__45212),
            .sr(N__45166));
    defparam \pid_front.error_p_reg_esr_RNID8VU1_3_LC_10_16_0 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNID8VU1_3_LC_10_16_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNID8VU1_3_LC_10_16_0 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pid_front.error_p_reg_esr_RNID8VU1_3_LC_10_16_0  (
            .in0(N__51623),
            .in1(N__51372),
            .in2(N__45120),
            .in3(N__54683),
            .lcout(\pid_front.error_p_reg_esr_RNID8VU1Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIUAE8_0_4_LC_10_16_1 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIUAE8_0_4_LC_10_16_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIUAE8_0_4_LC_10_16_1 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_front.error_p_reg_esr_RNIUAE8_0_4_LC_10_16_1  (
            .in0(N__45789),
            .in1(N__45771),
            .in2(_gnd_net_),
            .in3(N__49052),
            .lcout(\pid_front.error_p_reg_esr_RNIUAE8_0Z0Z_4 ),
            .ltout(\pid_front.error_p_reg_esr_RNIUAE8_0Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIMI772_3_LC_10_16_2 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIMI772_3_LC_10_16_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIMI772_3_LC_10_16_2 .LUT_INIT=16'b1111101010100000;
    LogicCell40 \pid_front.error_p_reg_esr_RNIMI772_3_LC_10_16_2  (
            .in0(N__51624),
            .in1(N__45801),
            .in2(N__45813),
            .in3(N__54684),
            .lcout(\pid_front.error_p_reg_esr_RNIMI772Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_4_LC_10_16_3 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_4_LC_10_16_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_4_LC_10_16_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_4_LC_10_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49053),
            .lcout(\pid_front.error_d_reg_prevZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87106),
            .ce(N__70482),
            .sr(N__70357));
    defparam \pid_front.error_p_reg_esr_RNIB9N71_0_5_LC_10_16_4 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIB9N71_0_5_LC_10_16_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIB9N71_0_5_LC_10_16_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_front.error_p_reg_esr_RNIB9N71_0_5_LC_10_16_4  (
            .in0(_gnd_net_),
            .in1(N__45743),
            .in2(_gnd_net_),
            .in3(N__55195),
            .lcout(\pid_front.error_p_reg_esr_RNIB9N71_0Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIUAE8_4_LC_10_16_5 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIUAE8_4_LC_10_16_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIUAE8_4_LC_10_16_5 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_front.error_p_reg_esr_RNIUAE8_4_LC_10_16_5  (
            .in0(N__45788),
            .in1(N__45770),
            .in2(_gnd_net_),
            .in3(N__49051),
            .lcout(\pid_front.error_p_reg_esr_RNIUAE8Z0Z_4 ),
            .ltout(\pid_front.error_p_reg_esr_RNIUAE8Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIVOSG_0_5_LC_10_16_6 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIVOSG_0_5_LC_10_16_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIVOSG_0_5_LC_10_16_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \pid_front.error_p_reg_esr_RNIVOSG_0_5_LC_10_16_6  (
            .in0(N__49023),
            .in1(N__45914),
            .in2(N__45762),
            .in3(N__48573),
            .lcout(\pid_front.error_p_reg_esr_RNIVOSG_0Z0Z_5 ),
            .ltout(\pid_front.error_p_reg_esr_RNIVOSG_0Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIB9N71_5_LC_10_16_7 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIB9N71_5_LC_10_16_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIB9N71_5_LC_10_16_7 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \pid_front.error_p_reg_esr_RNIB9N71_5_LC_10_16_7  (
            .in0(N__55196),
            .in1(_gnd_net_),
            .in2(N__45759),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_p_reg_esr_RNIB9N71Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI6B6F_0_6_LC_10_17_0 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI6B6F_0_6_LC_10_17_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI6B6F_0_6_LC_10_17_0 .LUT_INIT=16'b0010110111010010;
    LogicCell40 \pid_front.error_p_reg_esr_RNI6B6F_0_6_LC_10_17_0  (
            .in0(N__48567),
            .in1(N__49020),
            .in2(N__45855),
            .in3(N__45864),
            .lcout(\pid_front.error_p_reg_esr_RNI6B6F_0Z0Z_6 ),
            .ltout(\pid_front.error_p_reg_esr_RNI6B6F_0Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIU9ST_6_LC_10_17_1 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIU9ST_6_LC_10_17_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIU9ST_6_LC_10_17_1 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \pid_front.error_p_reg_esr_RNIU9ST_6_LC_10_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__45747),
            .in3(N__55151),
            .lcout(),
            .ltout(\pid_front.un1_pid_prereg_66_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI8CGM2_5_LC_10_17_2 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI8CGM2_5_LC_10_17_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI8CGM2_5_LC_10_17_2 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \pid_front.error_p_reg_esr_RNI8CGM2_5_LC_10_17_2  (
            .in0(N__55197),
            .in1(N__45744),
            .in2(N__45732),
            .in3(N__45872),
            .lcout(\pid_front.error_p_reg_esr_RNI8CGM2Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIT2PE1_5_LC_10_17_3 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIT2PE1_5_LC_10_17_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIT2PE1_5_LC_10_17_3 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_front.error_p_reg_esr_RNIT2PE1_5_LC_10_17_3  (
            .in0(N__45873),
            .in1(N__45933),
            .in2(_gnd_net_),
            .in3(N__55152),
            .lcout(\pid_front.error_p_reg_esr_RNIT2PE1Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIVOSG_5_LC_10_17_4 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIVOSG_5_LC_10_17_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIVOSG_5_LC_10_17_4 .LUT_INIT=16'b1111011001100000;
    LogicCell40 \pid_front.error_p_reg_esr_RNIVOSG_5_LC_10_17_4  (
            .in0(N__48568),
            .in1(N__49021),
            .in2(N__45918),
            .in3(N__45879),
            .lcout(\pid_front.error_p_reg_esr_RNIVOSGZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNI4SN6_6_LC_10_17_5 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNI4SN6_6_LC_10_17_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNI4SN6_6_LC_10_17_5 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNI4SN6_6_LC_10_17_5  (
            .in0(N__48100),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49778),
            .lcout(\pid_front.N_2155_i ),
            .ltout(\pid_front.N_2155_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI6B6F_6_LC_10_17_6 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI6B6F_6_LC_10_17_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI6B6F_6_LC_10_17_6 .LUT_INIT=16'b1101111100001101;
    LogicCell40 \pid_front.error_p_reg_esr_RNI6B6F_6_LC_10_17_6  (
            .in0(N__48569),
            .in1(N__49022),
            .in2(N__45858),
            .in3(N__45851),
            .lcout(\pid_front.error_p_reg_esr_RNI6B6FZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_6_LC_10_17_7 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_6_LC_10_17_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_6_LC_10_17_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_6_LC_10_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49779),
            .lcout(\pid_front.error_d_reg_prevZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87120),
            .ce(N__70471),
            .sr(N__70355));
    defparam \pid_front.error_d_reg_prev_esr_RNIQK6U_10_LC_10_18_0 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIQK6U_10_LC_10_18_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIQK6U_10_LC_10_18_0 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIQK6U_10_LC_10_18_0  (
            .in0(_gnd_net_),
            .in1(N__46519),
            .in2(_gnd_net_),
            .in3(N__46495),
            .lcout(),
            .ltout(\pid_front.N_2179_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIFM3D1_10_LC_10_18_1 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIFM3D1_10_LC_10_18_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIFM3D1_10_LC_10_18_1 .LUT_INIT=16'b0101101010010110;
    LogicCell40 \pid_front.error_p_reg_esr_RNIFM3D1_10_LC_10_18_1  (
            .in0(N__49515),
            .in1(N__46677),
            .in2(N__45831),
            .in3(N__46701),
            .lcout(\pid_front.error_p_reg_esr_RNIFM3D1Z0Z_10 ),
            .ltout(\pid_front.error_p_reg_esr_RNIFM3D1Z0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIS5CU3_9_LC_10_18_2 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIS5CU3_9_LC_10_18_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIS5CU3_9_LC_10_18_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pid_front.error_p_reg_esr_RNIS5CU3_9_LC_10_18_2  (
            .in0(N__45819),
            .in1(N__46022),
            .in2(N__45828),
            .in3(N__55007),
            .lcout(\pid_front.error_p_reg_esr_RNIS5CU3Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNILQ6F_9_LC_10_18_3 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNILQ6F_9_LC_10_18_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNILQ6F_9_LC_10_18_3 .LUT_INIT=16'b1000111011001111;
    LogicCell40 \pid_front.error_p_reg_esr_RNILQ6F_9_LC_10_18_3  (
            .in0(N__49688),
            .in1(N__46055),
            .in2(N__46647),
            .in3(N__48549),
            .lcout(\pid_front.error_p_reg_esr_RNILQ6FZ0Z_9 ),
            .ltout(\pid_front.error_p_reg_esr_RNILQ6FZ0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIEB5T7_9_LC_10_18_4 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIEB5T7_9_LC_10_18_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIEB5T7_9_LC_10_18_4 .LUT_INIT=16'b1111110011000000;
    LogicCell40 \pid_front.error_p_reg_esr_RNIEB5T7_9_LC_10_18_4  (
            .in0(N__46761),
            .in1(N__46074),
            .in2(N__46068),
            .in3(N__55008),
            .lcout(\pid_front.error_p_reg_esr_RNIEB5T7Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_10_LC_10_18_5 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_10_LC_10_18_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_10_LC_10_18_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_front.error_d_reg_prev_esr_10_LC_10_18_5  (
            .in0(N__46496),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_d_reg_prevZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87135),
            .ce(N__70469),
            .sr(N__70353));
    defparam \pid_front.error_p_reg_esr_RNILQ6F_0_9_LC_10_18_6 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNILQ6F_0_9_LC_10_18_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNILQ6F_0_9_LC_10_18_6 .LUT_INIT=16'b0011110010010110;
    LogicCell40 \pid_front.error_p_reg_esr_RNILQ6F_0_9_LC_10_18_6  (
            .in0(N__48548),
            .in1(N__46643),
            .in2(N__46056),
            .in3(N__49687),
            .lcout(\pid_front.error_p_reg_esr_RNILQ6F_0Z0Z_9 ),
            .ltout(\pid_front.error_p_reg_esr_RNILQ6F_0Z0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI6R6D1_8_LC_10_18_7 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI6R6D1_8_LC_10_18_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI6R6D1_8_LC_10_18_7 .LUT_INIT=16'b1111101010100000;
    LogicCell40 \pid_front.error_p_reg_esr_RNI6R6D1_8_LC_10_18_7  (
            .in0(N__48017),
            .in1(_gnd_net_),
            .in2(N__46026),
            .in3(N__55047),
            .lcout(\pid_front.error_p_reg_esr_RNI6R6D1Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIHDU52_0_22_LC_10_19_0 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIHDU52_0_22_LC_10_19_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIHDU52_0_22_LC_10_19_0 .LUT_INIT=16'b0010010011011011;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIHDU52_0_22_LC_10_19_0  (
            .in0(N__48312),
            .in1(N__46340),
            .in2(N__87429),
            .in3(N__56253),
            .lcout(\pid_front.un1_pid_prereg_0_15 ),
            .ltout(\pid_front.un1_pid_prereg_0_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIBLAI5_22_LC_10_19_1 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIBLAI5_22_LC_10_19_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIBLAI5_22_LC_10_19_1 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIBLAI5_22_LC_10_19_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__46008),
            .in3(N__45947),
            .lcout(\pid_front.error_d_reg_prev_esr_RNIBLAI5Z0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIF7HGD_19_LC_10_19_2 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIF7HGD_19_LC_10_19_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIF7HGD_19_LC_10_19_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_front.error_p_reg_esr_RNIF7HGD_19_LC_10_19_2  (
            .in0(N__45996),
            .in1(N__46121),
            .in2(N__45981),
            .in3(N__48367),
            .lcout(\pid_front.error_p_reg_esr_RNIF7HGDZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIQ7CC3_21_LC_10_19_3 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIQ7CC3_21_LC_10_19_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIQ7CC3_21_LC_10_19_3 .LUT_INIT=16'b1111101010100000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIQ7CC3_21_LC_10_19_3  (
            .in0(N__55695),
            .in1(_gnd_net_),
            .in2(N__48240),
            .in3(N__46131),
            .lcout(\pid_front.un1_pid_prereg_0_14 ),
            .ltout(\pid_front.un1_pid_prereg_0_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIOS1BC_22_LC_10_19_4 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIOS1BC_22_LC_10_19_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIOS1BC_22_LC_10_19_4 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIOS1BC_22_LC_10_19_4  (
            .in0(N__48369),
            .in1(N__46122),
            .in2(N__45936),
            .in3(N__46148),
            .lcout(\pid_front.error_d_reg_prev_esr_RNIOS1BCZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIDVE61_22_LC_10_19_5 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIDVE61_22_LC_10_19_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIDVE61_22_LC_10_19_5 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIDVE61_22_LC_10_19_5  (
            .in0(N__46339),
            .in1(N__87425),
            .in2(_gnd_net_),
            .in3(N__48311),
            .lcout(\pid_front.un1_pid_prereg_370_1 ),
            .ltout(\pid_front.un1_pid_prereg_370_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIQ7CC3_0_21_LC_10_19_6 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIQ7CC3_0_21_LC_10_19_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIQ7CC3_0_21_LC_10_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIQ7CC3_0_21_LC_10_19_6  (
            .in0(_gnd_net_),
            .in1(N__48236),
            .in2(N__46125),
            .in3(N__55694),
            .lcout(\pid_front.un1_pid_prereg_0_13 ),
            .ltout(\pid_front.un1_pid_prereg_0_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNID7NO6_20_LC_10_19_7 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNID7NO6_20_LC_10_19_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNID7NO6_20_LC_10_19_7 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \pid_front.error_p_reg_esr_RNID7NO6_20_LC_10_19_7  (
            .in0(N__48368),
            .in1(_gnd_net_),
            .in2(N__46113),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_p_reg_esr_RNID7NO6Z0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIETB61_3_13_LC_10_20_0 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIETB61_3_13_LC_10_20_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIETB61_3_13_LC_10_20_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_front.error_p_reg_esr_RNIETB61_3_13_LC_10_20_0  (
            .in0(N__48879),
            .in1(N__48820),
            .in2(_gnd_net_),
            .in3(N__48773),
            .lcout(\pid_front.N_4_1_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_fast_esr_RNIOTBC_12_LC_10_20_1 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_fast_esr_RNIOTBC_12_LC_10_20_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_fast_esr_RNIOTBC_12_LC_10_20_1 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \pid_front.error_d_reg_fast_esr_RNIOTBC_12_LC_10_20_1  (
            .in0(_gnd_net_),
            .in1(N__48522),
            .in2(_gnd_net_),
            .in3(N__46587),
            .lcout(),
            .ltout(\pid_front.g1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI6RNI1_13_LC_10_20_2 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI6RNI1_13_LC_10_20_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI6RNI1_13_LC_10_20_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \pid_front.error_p_reg_esr_RNI6RNI1_13_LC_10_20_2  (
            .in0(N__48880),
            .in1(N__48821),
            .in2(N__46101),
            .in3(N__48774),
            .lcout(),
            .ltout(\pid_front.g0_3_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIPCFV3_12_LC_10_20_3 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIPCFV3_12_LC_10_20_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIPCFV3_12_LC_10_20_3 .LUT_INIT=16'b1110000110000111;
    LogicCell40 \pid_front.error_p_reg_esr_RNIPCFV3_12_LC_10_20_3  (
            .in0(N__48968),
            .in1(N__46200),
            .in2(N__46098),
            .in3(N__49074),
            .lcout(\pid_front.g1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIJHNC2_12_LC_10_20_4 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIJHNC2_12_LC_10_20_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIJHNC2_12_LC_10_20_4 .LUT_INIT=16'b1001000011111001;
    LogicCell40 \pid_front.error_p_reg_esr_RNIJHNC2_12_LC_10_20_4  (
            .in0(N__49627),
            .in1(N__48653),
            .in2(N__46095),
            .in3(N__48967),
            .lcout(),
            .ltout(\pid_front.g0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIU52U6_12_LC_10_20_5 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIU52U6_12_LC_10_20_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIU52U6_12_LC_10_20_5 .LUT_INIT=16'b1101010000101011;
    LogicCell40 \pid_front.error_p_reg_esr_RNIU52U6_12_LC_10_20_5  (
            .in0(N__48600),
            .in1(N__46080),
            .in2(N__46218),
            .in3(N__46215),
            .lcout(),
            .ltout(\pid_front.error_p_reg_esr_RNIU52U6Z0Z_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIT79QC_12_LC_10_20_6 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIT79QC_12_LC_10_20_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIT79QC_12_LC_10_20_6 .LUT_INIT=16'b1000111000001100;
    LogicCell40 \pid_front.error_p_reg_esr_RNIT79QC_12_LC_10_20_6  (
            .in0(N__55464),
            .in1(N__55419),
            .in2(N__46209),
            .in3(N__46206),
            .lcout(\pid_front.error_p_reg_esr_RNIT79QCZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIUO6U_1_12_LC_10_20_7 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIUO6U_1_12_LC_10_20_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIUO6U_1_12_LC_10_20_7 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIUO6U_1_12_LC_10_20_7  (
            .in0(N__48652),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49626),
            .lcout(\pid_front.g1_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_5_LC_10_21_0 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_5_LC_10_21_0 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_5_LC_10_21_0 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \pid_front.error_i_reg_5_LC_10_21_0  (
            .in0(N__67533),
            .in1(N__55211),
            .in2(N__75537),
            .in3(N__59513),
            .lcout(\pid_front.error_i_regZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87183),
            .ce(),
            .sr(N__79664));
    defparam \pid_front.error_p_reg_esr_RNI873N_11_LC_10_21_2 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI873N_11_LC_10_21_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI873N_11_LC_10_21_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \pid_front.error_p_reg_esr_RNI873N_11_LC_10_21_2  (
            .in0(_gnd_net_),
            .in1(N__49129),
            .in2(_gnd_net_),
            .in3(N__49203),
            .lcout(\pid_front.un1_pid_prereg_79 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNICU3D1_0_6_LC_10_21_3 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNICU3D1_0_6_LC_10_21_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNICU3D1_0_6_LC_10_21_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_front.error_p_reg_esr_RNICU3D1_0_6_LC_10_21_3  (
            .in0(N__48083),
            .in1(N__46175),
            .in2(_gnd_net_),
            .in3(N__55114),
            .lcout(\pid_front.error_p_reg_esr_RNICU3D1_0Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNICU3D1_6_LC_10_21_4 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNICU3D1_6_LC_10_21_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNICU3D1_6_LC_10_21_4 .LUT_INIT=16'b1111101010100000;
    LogicCell40 \pid_front.error_p_reg_esr_RNICU3D1_6_LC_10_21_4  (
            .in0(N__55115),
            .in1(_gnd_net_),
            .in2(N__46179),
            .in3(N__48084),
            .lcout(\pid_front.error_p_reg_esr_RNICU3D1Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIETB61_0_13_LC_10_21_5 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIETB61_0_13_LC_10_21_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIETB61_0_13_LC_10_21_5 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_front.error_p_reg_esr_RNIETB61_0_13_LC_10_21_5  (
            .in0(N__48882),
            .in1(N__48815),
            .in2(_gnd_net_),
            .in3(N__48770),
            .lcout(\pid_front.N_2198_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIETB61_1_13_LC_10_21_6 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIETB61_1_13_LC_10_21_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIETB61_1_13_LC_10_21_6 .LUT_INIT=16'b1000111010001110;
    LogicCell40 \pid_front.error_p_reg_esr_RNIETB61_1_13_LC_10_21_6  (
            .in0(N__48772),
            .in1(N__48884),
            .in2(N__48822),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_p_reg_esr_RNIETB61_1Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIETB61_2_13_LC_10_21_7 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIETB61_2_13_LC_10_21_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIETB61_2_13_LC_10_21_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_front.error_p_reg_esr_RNIETB61_2_13_LC_10_21_7  (
            .in0(N__48883),
            .in1(N__48816),
            .in2(_gnd_net_),
            .in3(N__48771),
            .lcout(\pid_front.N_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_fast_esr_RNID6KB1_12_LC_10_22_0 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_fast_esr_RNID6KB1_12_LC_10_22_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_fast_esr_RNID6KB1_12_LC_10_22_0 .LUT_INIT=16'b1111011001100000;
    LogicCell40 \pid_front.error_d_reg_fast_esr_RNID6KB1_12_LC_10_22_0  (
            .in0(N__46582),
            .in1(N__48524),
            .in2(N__48972),
            .in3(N__48906),
            .lcout(),
            .ltout(\pid_front.error_d_reg_fast_esr_RNID6KB1Z0Z_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_fast_esr_RNIQSG63_12_LC_10_22_1 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_fast_esr_RNIQSG63_12_LC_10_22_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_fast_esr_RNIQSG63_12_LC_10_22_1 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \pid_front.error_d_reg_fast_esr_RNIQSG63_12_LC_10_22_1  (
            .in0(_gnd_net_),
            .in1(N__46350),
            .in2(N__46446),
            .in3(N__49245),
            .lcout(\pid_front.error_d_reg_fast_esr_RNIQSG63Z0Z_12 ),
            .ltout(\pid_front.error_d_reg_fast_esr_RNIQSG63Z0Z_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI8QSC4_13_LC_10_22_2 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI8QSC4_13_LC_10_22_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI8QSC4_13_LC_10_22_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \pid_front.error_p_reg_esr_RNI8QSC4_13_LC_10_22_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__46443),
            .in3(N__51919),
            .lcout(),
            .ltout(\pid_front.un1_pid_prereg_97_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI8C7GB_13_LC_10_22_3 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI8C7GB_13_LC_10_22_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI8C7GB_13_LC_10_22_3 .LUT_INIT=16'b1110111011101000;
    LogicCell40 \pid_front.error_p_reg_esr_RNI8C7GB_13_LC_10_22_3  (
            .in0(N__54213),
            .in1(N__46440),
            .in2(N__46434),
            .in3(N__46431),
            .lcout(\pid_front.error_p_reg_esr_RNI8C7GBZ0Z_13 ),
            .ltout(\pid_front.error_p_reg_esr_RNI8C7GBZ0Z_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIG7MLR_12_LC_10_22_4 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIG7MLR_12_LC_10_22_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIG7MLR_12_LC_10_22_4 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \pid_front.error_p_reg_esr_RNIG7MLR_12_LC_10_22_4  (
            .in0(_gnd_net_),
            .in1(N__46404),
            .in2(N__46389),
            .in3(N__46379),
            .lcout(\pid_front.error_p_reg_esr_RNIG7MLRZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_fast_esr_RNI5VGK_12_LC_10_22_5 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_fast_esr_RNI5VGK_12_LC_10_22_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_fast_esr_RNI5VGK_12_LC_10_22_5 .LUT_INIT=16'b1101110111101110;
    LogicCell40 \pid_front.error_d_reg_fast_esr_RNI5VGK_12_LC_10_22_5  (
            .in0(N__48523),
            .in1(N__48963),
            .in2(_gnd_net_),
            .in3(N__46581),
            .lcout(\pid_front.error_d_reg_fast_esr_RNI5VGKZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIHDU52_22_LC_10_22_6 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIHDU52_22_LC_10_22_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIHDU52_22_LC_10_22_6 .LUT_INIT=16'b1110111100001000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIHDU52_22_LC_10_22_6  (
            .in0(N__87403),
            .in1(N__48336),
            .in2(N__46344),
            .in3(N__56252),
            .lcout(\pid_front.un1_pid_prereg_0_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNI6J3B5_12_LC_10_22_7 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNI6J3B5_12_LC_10_22_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNI6J3B5_12_LC_10_22_7 .LUT_INIT=16'b1011010001001011;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNI6J3B5_12_LC_10_22_7  (
            .in0(N__49607),
            .in1(N__48657),
            .in2(N__51926),
            .in3(N__48614),
            .lcout(\pid_front.error_d_reg_prev_esr_RNI6J3B5Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_esr_10_LC_10_23_0 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_10_LC_10_23_0 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_10_LC_10_23_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_esr_10_LC_10_23_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46239),
            .lcout(\pid_front.error_d_regZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87215),
            .ce(N__86307),
            .sr(N__86011));
    defparam \pid_front.error_d_reg_esr_11_LC_10_23_1 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_11_LC_10_23_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_11_LC_10_23_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_esr_11_LC_10_23_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46629),
            .lcout(\pid_front.error_d_regZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87215),
            .ce(N__86307),
            .sr(N__86011));
    defparam \pid_front.error_d_reg_esr_9_LC_10_23_2 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_9_LC_10_23_2 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_9_LC_10_23_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_esr_9_LC_10_23_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46608),
            .lcout(\pid_front.error_d_regZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87215),
            .ce(N__86307),
            .sr(N__86011));
    defparam \pid_front.error_d_reg_fast_esr_12_LC_10_23_3 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_fast_esr_12_LC_10_23_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_fast_esr_12_LC_10_23_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_fast_esr_12_LC_10_23_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49656),
            .lcout(\pid_front.error_d_reg_fastZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87215),
            .ce(N__86307),
            .sr(N__86011));
    defparam \pid_front.error_d_reg_esr_13_LC_10_23_4 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_13_LC_10_23_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_13_LC_10_23_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_esr_13_LC_10_23_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46563),
            .lcout(\pid_front.error_d_regZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87215),
            .ce(N__86307),
            .sr(N__86011));
    defparam \pid_front.error_p_reg_esr_RNIKG5U_10_LC_10_24_0 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIKG5U_10_LC_10_24_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIKG5U_10_LC_10_24_0 .LUT_INIT=16'b1111101010110010;
    LogicCell40 \pid_front.error_p_reg_esr_RNIKG5U_10_LC_10_24_0  (
            .in0(N__46484),
            .in1(N__46662),
            .in2(N__49511),
            .in3(N__46694),
            .lcout(\pid_front.error_p_reg_esr_RNIKG5UZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIKG5U_0_10_LC_10_24_1 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIKG5U_0_10_LC_10_24_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIKG5U_0_10_LC_10_24_1 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \pid_front.error_p_reg_esr_RNIKG5U_0_10_LC_10_24_1  (
            .in0(N__46695),
            .in1(N__46485),
            .in2(N__46672),
            .in3(N__49507),
            .lcout(),
            .ltout(\pid_front.error_p_reg_esr_RNIKG5U_0Z0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNI379B2_10_LC_10_24_2 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNI379B2_10_LC_10_24_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNI379B2_10_LC_10_24_2 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNI379B2_10_LC_10_24_2  (
            .in0(_gnd_net_),
            .in1(N__46531),
            .in2(N__46548),
            .in3(N__46545),
            .lcout(\pid_front.error_d_reg_prev_esr_RNI379B2Z0Z_10 ),
            .ltout(\pid_front.error_d_reg_prev_esr_RNI379B2Z0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNI5JRF4_0_10_LC_10_24_3 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNI5JRF4_0_10_LC_10_24_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNI5JRF4_0_10_LC_10_24_3 .LUT_INIT=16'b1101001000101101;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNI5JRF4_0_10_LC_10_24_3  (
            .in0(N__46532),
            .in1(N__46486),
            .in2(N__46464),
            .in3(N__46461),
            .lcout(\pid_front.error_d_reg_prev_esr_RNI5JRF4_0Z0Z_10 ),
            .ltout(\pid_front.error_d_reg_prev_esr_RNI5JRF4_0Z0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIO00C5_0_10_LC_10_24_4 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIO00C5_0_10_LC_10_24_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIO00C5_0_10_LC_10_24_4 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIO00C5_0_10_LC_10_24_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__46764),
            .in3(N__54963),
            .lcout(\pid_front.error_d_reg_prev_esr_RNIO00C5_0Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIO00C5_10_LC_10_24_5 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIO00C5_10_LC_10_24_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIO00C5_10_LC_10_24_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIO00C5_10_LC_10_24_5  (
            .in0(N__54964),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46727),
            .lcout(\pid_front.error_d_reg_prev_esr_RNIO00C5Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_9_LC_10_24_6 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_9_LC_10_24_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_9_LC_10_24_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_9_LC_10_24_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46697),
            .lcout(\pid_front.error_d_reg_prevZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87228),
            .ce(N__70494),
            .sr(N__70347));
    defparam \pid_front.error_d_reg_prev_esr_RNIA2O6_9_LC_10_24_7 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIA2O6_9_LC_10_24_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIA2O6_9_LC_10_24_7 .LUT_INIT=16'b1010010110100101;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIA2O6_9_LC_10_24_7  (
            .in0(N__46696),
            .in1(_gnd_net_),
            .in2(N__46673),
            .in3(_gnd_net_),
            .lcout(\pid_front.N_2173_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_prereg_esr_11_LC_10_25_0 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_11_LC_10_25_0 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_11_LC_10_25_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_11_LC_10_25_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54971),
            .lcout(\pid_front.error_i_acumm_preregZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87242),
            .ce(N__56075),
            .sr(N__79685));
    defparam \pid_front.error_i_acumm_prereg_esr_2_LC_10_25_1 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_2_LC_10_25_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_2_LC_10_25_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_2_LC_10_25_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54761),
            .lcout(\pid_front.error_i_acumm_preregZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87242),
            .ce(N__56075),
            .sr(N__79685));
    defparam \pid_front.error_i_acumm_prereg_esr_4_LC_10_25_2 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_4_LC_10_25_2 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_4_LC_10_25_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_4_LC_10_25_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54682),
            .lcout(\pid_front.error_i_acumm_preregZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87242),
            .ce(N__56075),
            .sr(N__79685));
    defparam \pid_front.error_i_acumm_prereg_esr_5_LC_10_25_3 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_5_LC_10_25_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_5_LC_10_25_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_5_LC_10_25_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55194),
            .lcout(\pid_front.error_i_acumm_preregZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87242),
            .ce(N__56075),
            .sr(N__79685));
    defparam \pid_front.error_i_acumm_prereg_esr_6_LC_10_25_4 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_6_LC_10_25_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_6_LC_10_25_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_6_LC_10_25_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55150),
            .lcout(\pid_front.error_i_acumm_preregZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87242),
            .ce(N__56075),
            .sr(N__79685));
    defparam \pid_front.error_i_acumm_prereg_esr_7_LC_10_25_5 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_7_LC_10_25_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_7_LC_10_25_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_7_LC_10_25_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55116),
            .lcout(\pid_front.error_i_acumm_preregZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87242),
            .ce(N__56075),
            .sr(N__79685));
    defparam \pid_front.error_i_acumm_prereg_esr_10_LC_10_25_7 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_10_LC_10_25_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_10_LC_10_25_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_10_LC_10_25_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55006),
            .lcout(\pid_front.error_i_acumm_preregZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87242),
            .ce(N__56075),
            .sr(N__79685));
    defparam \pid_front.state_RNIPKTD_0_LC_10_27_4 .C_ON=1'b0;
    defparam \pid_front.state_RNIPKTD_0_LC_10_27_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.state_RNIPKTD_0_LC_10_27_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \pid_front.state_RNIPKTD_0_LC_10_27_4  (
            .in0(_gnd_net_),
            .in1(N__60185),
            .in2(_gnd_net_),
            .in3(N__79916),
            .lcout(\pid_front.state_RNIPKTDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIB3GR1_2_LC_11_1_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIB3GR1_2_LC_11_1_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIB3GR1_2_LC_11_1_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIB3GR1_2_LC_11_1_0  (
            .in0(_gnd_net_),
            .in1(N__46818),
            .in2(N__53965),
            .in3(N__57330),
            .lcout(\ppm_encoder_1.N_39_i ),
            .ltout(),
            .carryin(bfn_11_1_0_),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_1_LC_11_1_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_1_LC_11_1_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_1_LC_11_1_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_1_LC_11_1_1  (
            .in0(_gnd_net_),
            .in1(N__49947),
            .in2(_gnd_net_),
            .in3(N__46812),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_1 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_0 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_2_LC_11_1_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_2_LC_11_1_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_2_LC_11_1_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_2_LC_11_1_2  (
            .in0(_gnd_net_),
            .in1(N__57647),
            .in2(N__57285),
            .in3(N__46809),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_2 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_1 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_3_LC_11_1_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_3_LC_11_1_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_3_LC_11_1_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_3_LC_11_1_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__49941),
            .in3(N__46800),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_3 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_2 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_4_LC_11_1_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_4_LC_11_1_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_4_LC_11_1_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_4_LC_11_1_4  (
            .in0(_gnd_net_),
            .in1(N__53004),
            .in2(_gnd_net_),
            .in3(N__46791),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_4 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_3 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_5_LC_11_1_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_5_LC_11_1_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_5_LC_11_1_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_5_LC_11_1_5  (
            .in0(_gnd_net_),
            .in1(N__46788),
            .in2(_gnd_net_),
            .in3(N__46776),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_5 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_4 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_6_LC_11_1_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_6_LC_11_1_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_6_LC_11_1_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_6_LC_11_1_6  (
            .in0(_gnd_net_),
            .in1(N__50240),
            .in2(N__50055),
            .in3(N__46767),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_6 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_5 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_7_LC_11_1_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_7_LC_11_1_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_7_LC_11_1_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_7_LC_11_1_7  (
            .in0(_gnd_net_),
            .in1(N__46923),
            .in2(_gnd_net_),
            .in3(N__46905),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_7 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_6 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_8_LC_11_2_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_8_LC_11_2_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_8_LC_11_2_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_8_LC_11_2_0  (
            .in0(_gnd_net_),
            .in1(N__46902),
            .in2(_gnd_net_),
            .in3(N__46884),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_8 ),
            .ltout(),
            .carryin(bfn_11_2_0_),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_9_LC_11_2_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_9_LC_11_2_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_9_LC_11_2_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_9_LC_11_2_1  (
            .in0(_gnd_net_),
            .in1(N__63282),
            .in2(_gnd_net_),
            .in3(N__46881),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_9 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_8 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_10_LC_11_2_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_10_LC_11_2_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_10_LC_11_2_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_10_LC_11_2_2  (
            .in0(_gnd_net_),
            .in1(N__49932),
            .in2(_gnd_net_),
            .in3(N__46878),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_10 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_9 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_11_LC_11_2_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_11_LC_11_2_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_11_LC_11_2_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_11_LC_11_2_3  (
            .in0(_gnd_net_),
            .in1(N__46875),
            .in2(_gnd_net_),
            .in3(N__46863),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_11 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_10 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_12_LC_11_2_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_12_LC_11_2_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_12_LC_11_2_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_12_LC_11_2_4  (
            .in0(_gnd_net_),
            .in1(N__50046),
            .in2(_gnd_net_),
            .in3(N__46854),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_12 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_11 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_13_LC_11_2_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_13_LC_11_2_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_13_LC_11_2_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_13_LC_11_2_5  (
            .in0(_gnd_net_),
            .in1(N__53437),
            .in2(N__50007),
            .in3(N__46851),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_13 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_12 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_14_LC_11_2_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_14_LC_11_2_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_14_LC_11_2_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_14_LC_11_2_6  (
            .in0(_gnd_net_),
            .in1(N__46848),
            .in2(_gnd_net_),
            .in3(N__46836),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_14 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_13 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_15_LC_11_2_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_15_LC_11_2_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_15_LC_11_2_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_15_LC_11_2_7  (
            .in0(_gnd_net_),
            .in1(N__46953),
            .in2(_gnd_net_),
            .in3(N__46965),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_15 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_14 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_16_LC_11_3_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_16_LC_11_3_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_16_LC_11_3_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_16_LC_11_3_0  (
            .in0(_gnd_net_),
            .in1(N__46947),
            .in2(_gnd_net_),
            .in3(N__46962),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_16 ),
            .ltout(),
            .carryin(bfn_11_3_0_),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_17_LC_11_3_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_17_LC_11_3_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_17_LC_11_3_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_17_LC_11_3_1  (
            .in0(_gnd_net_),
            .in1(N__61080),
            .in2(_gnd_net_),
            .in3(N__46959),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_17 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_16 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_18_LC_11_3_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNO_1_18_LC_11_3_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_18_LC_11_3_2 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_18_LC_11_3_2  (
            .in0(N__60608),
            .in1(N__56948),
            .in2(_gnd_net_),
            .in3(N__46956),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_LC_11_3_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_LC_11_3_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_LC_11_3_3 .LUT_INIT=16'b0011000000010010;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_1_LC_11_3_3  (
            .in0(N__61627),
            .in1(N__79983),
            .in2(N__61396),
            .in3(N__64295),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__86978),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNIV9SJ1_LC_11_3_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNIV9SJ1_LC_11_3_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNIV9SJ1_LC_11_3_4 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_57_c_RNIV9SJ1_LC_11_3_4  (
            .in0(N__64598),
            .in1(N__61105),
            .in2(N__68670),
            .in3(N__61161),
            .lcout(\ppm_encoder_1.counter24_0_I_57_c_RNIV9SJZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIH8MT_0_15_LC_11_3_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIH8MT_0_15_LC_11_3_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIH8MT_0_15_LC_11_3_5 .LUT_INIT=16'b1100110001101100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIH8MT_0_15_LC_11_3_5  (
            .in0(N__64595),
            .in1(N__64654),
            .in2(N__63450),
            .in3(N__64293),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNII9MT_16_LC_11_3_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNII9MT_16_LC_11_3_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNII9MT_16_LC_11_3_7 .LUT_INIT=16'b1111000001111000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNII9MT_16_LC_11_3_7  (
            .in0(N__64596),
            .in1(N__63388),
            .in2(N__63935),
            .in3(N__64294),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_15_LC_11_4_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_15_LC_11_4_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.init_pulses_15_LC_11_4_1 .LUT_INIT=16'b0011000100100000;
    LogicCell40 \ppm_encoder_1.init_pulses_15_LC_11_4_1  (
            .in0(N__55940),
            .in1(N__55774),
            .in2(N__46941),
            .in3(N__46929),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__86984),
            .ce(),
            .sr(N__79562));
    defparam \ppm_encoder_1.init_pulses_16_LC_11_4_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_16_LC_11_4_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.init_pulses_16_LC_11_4_2 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \ppm_encoder_1.init_pulses_16_LC_11_4_2  (
            .in0(N__55775),
            .in1(N__55944),
            .in2(N__47070),
            .in3(N__47061),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__86984),
            .ce(),
            .sr(N__79562));
    defparam \ppm_encoder_1.init_pulses_17_LC_11_4_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_17_LC_11_4_3 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_17_LC_11_4_3 .LUT_INIT=16'b0010001100100000;
    LogicCell40 \ppm_encoder_1.init_pulses_17_LC_11_4_3  (
            .in0(N__47055),
            .in1(N__55776),
            .in2(N__55955),
            .in3(N__47049),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__86984),
            .ce(),
            .sr(N__79562));
    defparam \ppm_encoder_1.init_pulses_18_LC_11_4_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_18_LC_11_4_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.init_pulses_18_LC_11_4_4 .LUT_INIT=16'b0000101100001000;
    LogicCell40 \ppm_encoder_1.init_pulses_18_LC_11_4_4  (
            .in0(N__47043),
            .in1(N__55942),
            .in2(N__55803),
            .in3(N__47037),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__86984),
            .ce(),
            .sr(N__79562));
    defparam \ppm_encoder_1.init_pulses_1_LC_11_4_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_1_LC_11_4_5 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_1_LC_11_4_5 .LUT_INIT=16'b0011001000000010;
    LogicCell40 \ppm_encoder_1.init_pulses_1_LC_11_4_5  (
            .in0(N__47031),
            .in1(N__55780),
            .in2(N__55956),
            .in3(N__47025),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__86984),
            .ce(),
            .sr(N__79562));
    defparam \ppm_encoder_1.init_pulses_10_LC_11_4_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_10_LC_11_4_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.init_pulses_10_LC_11_4_6 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \ppm_encoder_1.init_pulses_10_LC_11_4_6  (
            .in0(N__55773),
            .in1(N__55943),
            .in2(N__47016),
            .in3(N__47004),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__86984),
            .ce(),
            .sr(N__79562));
    defparam \ppm_encoder_1.init_pulses_9_LC_11_4_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_9_LC_11_4_7 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_9_LC_11_4_7 .LUT_INIT=16'b0011000100100000;
    LogicCell40 \ppm_encoder_1.init_pulses_9_LC_11_4_7  (
            .in0(N__55941),
            .in1(N__55781),
            .in2(N__46995),
            .in3(N__46980),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__86984),
            .ce(),
            .sr(N__79562));
    defparam \ppm_encoder_1.init_pulses_RNICIVR4_9_LC_11_5_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNICIVR4_9_LC_11_5_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNICIVR4_9_LC_11_5_0 .LUT_INIT=16'b0101101001101001;
    LogicCell40 \ppm_encoder_1.init_pulses_RNICIVR4_9_LC_11_5_0  (
            .in0(N__56947),
            .in1(N__47100),
            .in2(N__63500),
            .in3(N__50064),
            .lcout(),
            .ltout(\ppm_encoder_1.un1_init_pulses_0_axb_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIEBKU5_9_LC_11_5_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIEBKU5_9_LC_11_5_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIEBKU5_9_LC_11_5_1 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIEBKU5_9_LC_11_5_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__46974),
            .in3(N__47135),
            .lcout(\ppm_encoder_1.init_pulses_RNIEBKU5Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNIGD6O_9_LC_11_5_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNIGD6O_9_LC_11_5_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNIGD6O_9_LC_11_5_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \ppm_encoder_1.elevator_RNIGD6O_9_LC_11_5_2  (
            .in0(N__52909),
            .in1(N__47388),
            .in2(_gnd_net_),
            .in3(N__52792),
            .lcout(\ppm_encoder_1.elevator_RNIGD6OZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNIOEGE_10_LC_11_5_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNIOEGE_10_LC_11_5_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNIOEGE_10_LC_11_5_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \ppm_encoder_1.elevator_RNIOEGE_10_LC_11_5_3  (
            .in0(N__52793),
            .in1(N__56780),
            .in2(_gnd_net_),
            .in3(N__52910),
            .lcout(\ppm_encoder_1.elevator_RNIOEGEZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNI2PK21_9_LC_11_5_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI2PK21_9_LC_11_5_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI2PK21_9_LC_11_5_4 .LUT_INIT=16'b1111000001111000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI2PK21_9_LC_11_5_4  (
            .in0(N__61041),
            .in1(N__60931),
            .in2(N__63499),
            .in3(N__64270),
            .lcout(\ppm_encoder_1.N_265_i_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIRT0E1_9_LC_11_5_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIRT0E1_9_LC_11_5_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIRT0E1_9_LC_11_5_5 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \ppm_encoder_1.throttle_RNIRT0E1_9_LC_11_5_5  (
            .in0(N__47415),
            .in1(N__58004),
            .in2(N__47124),
            .in3(N__57159),
            .lcout(\ppm_encoder_1.un2_throttle_iv_0_1_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_LC_11_5_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_LC_11_5_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_LC_11_5_6 .LUT_INIT=16'b1110111011111100;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_LC_11_5_6  (
            .in0(N__52911),
            .in1(N__79985),
            .in2(N__57453),
            .in3(N__64271),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__86992),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNIB86O_4_LC_11_5_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNIB86O_4_LC_11_5_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNIB86O_4_LC_11_5_7 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \ppm_encoder_1.elevator_RNIB86O_4_LC_11_5_7  (
            .in0(N__52791),
            .in1(N__47094),
            .in2(_gnd_net_),
            .in3(N__52908),
            .lcout(\ppm_encoder_1.elevator_RNIB86OZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m9_0_i_LC_11_6_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m9_0_i_LC_11_6_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m9_0_i_LC_11_6_0 .LUT_INIT=16'b1101110110011001;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m9_0_i_LC_11_6_0  (
            .in0(N__64597),
            .in1(N__63449),
            .in2(_gnd_net_),
            .in3(N__63592),
            .lcout(\ppm_encoder_1.m9_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.rudder_RNIM1KQ_12_LC_11_6_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_RNIM1KQ_12_LC_11_6_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.rudder_RNIM1KQ_12_LC_11_6_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \ppm_encoder_1.rudder_RNIM1KQ_12_LC_11_6_1  (
            .in0(_gnd_net_),
            .in1(N__63779),
            .in2(_gnd_net_),
            .in3(N__50473),
            .lcout(),
            .ltout(\ppm_encoder_1.rudder_RNIM1KQZ0Z_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNIJBB92_12_LC_11_6_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNIJBB92_12_LC_11_6_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNIJBB92_12_LC_11_6_2 .LUT_INIT=16'b1111111111110001;
    LogicCell40 \ppm_encoder_1.elevator_RNIJBB92_12_LC_11_6_2  (
            .in0(N__47286),
            .in1(N__63591),
            .in2(N__47076),
            .in3(N__57067),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_2_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIRE0G4_12_LC_11_6_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIRE0G4_12_LC_11_6_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIRE0G4_12_LC_11_6_3 .LUT_INIT=16'b1001100110010110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIRE0G4_12_LC_11_6_3  (
            .in0(N__50443),
            .in1(N__56940),
            .in2(N__47073),
            .in3(N__47208),
            .lcout(),
            .ltout(\ppm_encoder_1.un1_init_pulses_0_axb_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNI7OHF5_12_LC_11_6_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI7OHF5_12_LC_11_6_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI7OHF5_12_LC_11_6_4 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI7OHF5_12_LC_11_6_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__47319),
            .in3(N__47312),
            .lcout(\ppm_encoder_1.init_pulses_RNI7OHF5Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter_RNIUS1G_4_LC_11_6_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter_RNIUS1G_4_LC_11_6_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter_RNIUS1G_4_LC_11_6_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \ppm_encoder_1.counter_RNIUS1G_4_LC_11_6_5  (
            .in0(N__64923),
            .in1(N__64893),
            .in2(N__64860),
            .in3(N__64953),
            .lcout(\ppm_encoder_1.un1_PPM_STATE_0_sqmuxa_0_i_a2_18_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_12_LC_11_7_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_12_LC_11_7_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_12_LC_11_7_0 .LUT_INIT=16'b0011111100010101;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_12_LC_11_7_0  (
            .in0(N__47284),
            .in1(N__47224),
            .in2(N__68674),
            .in3(N__63593),
            .lcout(\ppm_encoder_1.pulses2count_9_0_3_1_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_12_LC_11_7_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_12_LC_11_7_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_12_LC_11_7_2 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \ppm_encoder_1.throttle_12_LC_11_7_2  (
            .in0(N__47265),
            .in1(N__47241),
            .in2(N__47229),
            .in3(N__65168),
            .lcout(\ppm_encoder_1.throttleZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87006),
            .ce(),
            .sr(N__79577));
    defparam \ppm_encoder_1.throttle_RNIF0NE1_12_LC_11_7_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIF0NE1_12_LC_11_7_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIF0NE1_12_LC_11_7_3 .LUT_INIT=16'b0101110100001100;
    LogicCell40 \ppm_encoder_1.throttle_RNIF0NE1_12_LC_11_7_3  (
            .in0(N__60367),
            .in1(N__58014),
            .in2(N__47228),
            .in3(N__57184),
            .lcout(\ppm_encoder_1.un2_throttle_iv_0_1_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_11_LC_11_7_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_11_LC_11_7_5 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.aileron_11_LC_11_7_5 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.aileron_11_LC_11_7_5  (
            .in0(N__53856),
            .in1(N__47475),
            .in2(N__65264),
            .in3(N__60292),
            .lcout(\ppm_encoder_1.aileronZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87006),
            .ce(),
            .sr(N__79577));
    defparam \ppm_encoder_1.aileron_13_LC_11_7_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_13_LC_11_7_6 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.aileron_13_LC_11_7_6 .LUT_INIT=16'b1001100111110000;
    LogicCell40 \ppm_encoder_1.aileron_13_LC_11_7_6  (
            .in0(N__58314),
            .in1(N__47460),
            .in2(N__61307),
            .in3(N__65167),
            .lcout(\ppm_encoder_1.aileronZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87006),
            .ce(),
            .sr(N__79577));
    defparam \ppm_encoder_1.throttle_7_LC_11_8_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_7_LC_11_8_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_7_LC_11_8_2 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.throttle_7_LC_11_8_2  (
            .in0(N__47202),
            .in1(N__47193),
            .in2(N__65273),
            .in3(N__53647),
            .lcout(\ppm_encoder_1.throttleZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87014),
            .ce(),
            .sr(N__79585));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_8_LC_11_8_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_8_LC_11_8_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_8_LC_11_8_3 .LUT_INIT=16'b0010011100000000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_8_LC_11_8_3  (
            .in0(N__61629),
            .in1(N__47158),
            .in2(N__47441),
            .in3(N__61395),
            .lcout(\ppm_encoder_1.pulses2count_9_i_1_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_8_LC_11_8_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_8_LC_11_8_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.aileron_8_LC_11_8_4 .LUT_INIT=16'b0011101011001010;
    LogicCell40 \ppm_encoder_1.aileron_8_LC_11_8_4  (
            .in0(N__47437),
            .in1(N__53748),
            .in2(N__65272),
            .in3(N__47511),
            .lcout(\ppm_encoder_1.aileronZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87014),
            .ce(),
            .sr(N__79585));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_9_LC_11_8_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_9_LC_11_8_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_9_LC_11_8_6 .LUT_INIT=16'b0000101000100010;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_9_LC_11_8_6  (
            .in0(N__61394),
            .in1(N__47407),
            .in2(N__47387),
            .in3(N__61630),
            .lcout(\ppm_encoder_1.pulses2count_9_i_1_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_0_c_LC_11_9_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_0_c_LC_11_9_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_0_c_LC_11_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_0_c_LC_11_9_0  (
            .in0(_gnd_net_),
            .in1(N__53810),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_9_0_),
            .carryout(\ppm_encoder_1.un1_aileron_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_0_THRU_LUT4_0_LC_11_9_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_0_THRU_LUT4_0_LC_11_9_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_0_THRU_LUT4_0_LC_11_9_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_0_THRU_LUT4_0_LC_11_9_1  (
            .in0(_gnd_net_),
            .in1(N__53828),
            .in2(N__56552),
            .in3(N__47361),
            .lcout(\ppm_encoder_1.un1_aileron_cry_0_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_0 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_1_THRU_LUT4_0_LC_11_9_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_1_THRU_LUT4_0_LC_11_9_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_1_THRU_LUT4_0_LC_11_9_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_1_THRU_LUT4_0_LC_11_9_2  (
            .in0(_gnd_net_),
            .in1(N__58182),
            .in2(_gnd_net_),
            .in3(N__47352),
            .lcout(\ppm_encoder_1.un1_aileron_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_1 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_2_THRU_LUT4_0_LC_11_9_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_2_THRU_LUT4_0_LC_11_9_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_2_THRU_LUT4_0_LC_11_9_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_2_THRU_LUT4_0_LC_11_9_3  (
            .in0(_gnd_net_),
            .in1(N__53871),
            .in2(N__56553),
            .in3(N__47349),
            .lcout(\ppm_encoder_1.un1_aileron_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_2 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_3_THRU_LUT4_0_LC_11_9_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_3_THRU_LUT4_0_LC_11_9_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_3_THRU_LUT4_0_LC_11_9_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_3_THRU_LUT4_0_LC_11_9_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__53769),
            .in3(N__47340),
            .lcout(\ppm_encoder_1.un1_aileron_cry_3_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_3 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_4_THRU_LUT4_0_LC_11_9_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_4_THRU_LUT4_0_LC_11_9_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_4_THRU_LUT4_0_LC_11_9_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_4_THRU_LUT4_0_LC_11_9_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__53534),
            .in3(N__47325),
            .lcout(\ppm_encoder_1.un1_aileron_cry_4_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_4 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_5_THRU_LUT4_0_LC_11_9_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_5_THRU_LUT4_0_LC_11_9_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_5_THRU_LUT4_0_LC_11_9_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_5_THRU_LUT4_0_LC_11_9_6  (
            .in0(_gnd_net_),
            .in1(N__56514),
            .in2(N__58203),
            .in3(N__47322),
            .lcout(\ppm_encoder_1.un1_aileron_cry_5_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_5 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_6_THRU_LUT4_0_LC_11_9_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_6_THRU_LUT4_0_LC_11_9_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_6_THRU_LUT4_0_LC_11_9_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_6_THRU_LUT4_0_LC_11_9_7  (
            .in0(_gnd_net_),
            .in1(N__53511),
            .in2(_gnd_net_),
            .in3(N__47514),
            .lcout(\ppm_encoder_1.un1_aileron_cry_6_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_6 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_7_THRU_LUT4_0_LC_11_10_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_7_THRU_LUT4_0_LC_11_10_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_7_THRU_LUT4_0_LC_11_10_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_7_THRU_LUT4_0_LC_11_10_0  (
            .in0(_gnd_net_),
            .in1(N__53744),
            .in2(_gnd_net_),
            .in3(N__47502),
            .lcout(\ppm_encoder_1.un1_aileron_cry_7_THRU_CO ),
            .ltout(),
            .carryin(bfn_11_10_0_),
            .carryout(\ppm_encoder_1.un1_aileron_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_8_THRU_LUT4_0_LC_11_10_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_8_THRU_LUT4_0_LC_11_10_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_8_THRU_LUT4_0_LC_11_10_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_8_THRU_LUT4_0_LC_11_10_1  (
            .in0(_gnd_net_),
            .in1(N__53726),
            .in2(_gnd_net_),
            .in3(N__47493),
            .lcout(\ppm_encoder_1.un1_aileron_cry_8_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_8 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_9_THRU_LUT4_0_LC_11_10_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_9_THRU_LUT4_0_LC_11_10_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_9_THRU_LUT4_0_LC_11_10_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_9_THRU_LUT4_0_LC_11_10_2  (
            .in0(_gnd_net_),
            .in1(N__53786),
            .in2(_gnd_net_),
            .in3(N__47478),
            .lcout(\ppm_encoder_1.un1_aileron_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_9 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_10_THRU_LUT4_0_LC_11_10_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_10_THRU_LUT4_0_LC_11_10_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_10_THRU_LUT4_0_LC_11_10_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_10_THRU_LUT4_0_LC_11_10_3  (
            .in0(_gnd_net_),
            .in1(N__53855),
            .in2(_gnd_net_),
            .in3(N__47466),
            .lcout(\ppm_encoder_1.un1_aileron_cry_10_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_10 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_11_THRU_LUT4_0_LC_11_10_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_11_THRU_LUT4_0_LC_11_10_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_11_THRU_LUT4_0_LC_11_10_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_11_THRU_LUT4_0_LC_11_10_4  (
            .in0(_gnd_net_),
            .in1(N__58328),
            .in2(_gnd_net_),
            .in3(N__47463),
            .lcout(\ppm_encoder_1.un1_aileron_cry_11_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_11 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_12_THRU_LUT4_0_LC_11_10_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_12_THRU_LUT4_0_LC_11_10_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_12_THRU_LUT4_0_LC_11_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_12_THRU_LUT4_0_LC_11_10_5  (
            .in0(_gnd_net_),
            .in1(N__58310),
            .in2(N__56483),
            .in3(N__47451),
            .lcout(\ppm_encoder_1.un1_aileron_cry_12_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_12 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_esr_14_LC_11_10_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_esr_14_LC_11_10_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.aileron_esr_14_LC_11_10_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.aileron_esr_14_LC_11_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47448),
            .lcout(\ppm_encoder_1.aileronZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87029),
            .ce(N__50154),
            .sr(N__79595));
    defparam \uart_drone.data_Aux_0_LC_11_11_0 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_0_LC_11_11_0 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_Aux_0_LC_11_11_0 .LUT_INIT=16'b1100110011100100;
    LogicCell40 \uart_drone.data_Aux_0_LC_11_11_0  (
            .in0(N__62025),
            .in1(N__47540),
            .in2(N__47996),
            .in3(N__47582),
            .lcout(\uart_drone.data_AuxZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87039),
            .ce(),
            .sr(N__47556));
    defparam \uart_drone.data_Aux_1_LC_11_11_1 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_1_LC_11_11_1 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_Aux_1_LC_11_11_1 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \uart_drone.data_Aux_1_LC_11_11_1  (
            .in0(N__47583),
            .in1(N__47989),
            .in2(N__47529),
            .in3(N__50403),
            .lcout(\uart_drone.data_AuxZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87039),
            .ce(),
            .sr(N__47556));
    defparam \uart_drone.data_Aux_2_LC_11_11_2 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_2_LC_11_11_2 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_Aux_2_LC_11_11_2 .LUT_INIT=16'b1111000010111000;
    LogicCell40 \uart_drone.data_Aux_2_LC_11_11_2  (
            .in0(N__47986),
            .in1(N__50394),
            .in2(N__47718),
            .in3(N__47584),
            .lcout(\uart_drone.data_AuxZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87039),
            .ce(),
            .sr(N__47556));
    defparam \uart_drone.data_Aux_3_LC_11_11_3 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_3_LC_11_11_3 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_Aux_3_LC_11_11_3 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \uart_drone.data_Aux_3_LC_11_11_3  (
            .in0(N__47585),
            .in1(N__47990),
            .in2(N__47703),
            .in3(N__47595),
            .lcout(\uart_drone.data_AuxZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87039),
            .ce(),
            .sr(N__47556));
    defparam \uart_drone.data_Aux_4_LC_11_11_4 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_4_LC_11_11_4 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_Aux_4_LC_11_11_4 .LUT_INIT=16'b1111000010111000;
    LogicCell40 \uart_drone.data_Aux_4_LC_11_11_4  (
            .in0(N__47987),
            .in1(N__50640),
            .in2(N__47688),
            .in3(N__47586),
            .lcout(\uart_drone.data_AuxZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87039),
            .ce(),
            .sr(N__47556));
    defparam \uart_drone.data_Aux_5_LC_11_11_5 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_5_LC_11_11_5 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_Aux_5_LC_11_11_5 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \uart_drone.data_Aux_5_LC_11_11_5  (
            .in0(N__47587),
            .in1(N__47991),
            .in2(N__47673),
            .in3(N__50628),
            .lcout(\uart_drone.data_AuxZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87039),
            .ce(),
            .sr(N__47556));
    defparam \uart_drone.data_Aux_6_LC_11_11_6 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_6_LC_11_11_6 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_Aux_6_LC_11_11_6 .LUT_INIT=16'b1111000010111000;
    LogicCell40 \uart_drone.data_Aux_6_LC_11_11_6  (
            .in0(N__47988),
            .in1(N__50616),
            .in2(N__47658),
            .in3(N__47588),
            .lcout(\uart_drone.data_AuxZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87039),
            .ce(),
            .sr(N__47556));
    defparam \uart_drone.data_Aux_7_LC_11_11_7 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_7_LC_11_11_7 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_Aux_7_LC_11_11_7 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \uart_drone.data_Aux_7_LC_11_11_7  (
            .in0(N__47589),
            .in1(N__47992),
            .in2(N__47643),
            .in3(N__50857),
            .lcout(\uart_drone.data_AuxZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87039),
            .ce(),
            .sr(N__47556));
    defparam \uart_drone.data_esr_0_LC_11_12_0 .C_ON=1'b0;
    defparam \uart_drone.data_esr_0_LC_11_12_0 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_esr_0_LC_11_12_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone.data_esr_0_LC_11_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47541),
            .lcout(uart_drone_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87048),
            .ce(N__47628),
            .sr(N__47616));
    defparam \uart_drone.data_esr_1_LC_11_12_1 .C_ON=1'b0;
    defparam \uart_drone.data_esr_1_LC_11_12_1 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_esr_1_LC_11_12_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone.data_esr_1_LC_11_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47528),
            .lcout(uart_drone_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87048),
            .ce(N__47628),
            .sr(N__47616));
    defparam \uart_drone.data_esr_2_LC_11_12_2 .C_ON=1'b0;
    defparam \uart_drone.data_esr_2_LC_11_12_2 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_esr_2_LC_11_12_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone.data_esr_2_LC_11_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47717),
            .lcout(uart_drone_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87048),
            .ce(N__47628),
            .sr(N__47616));
    defparam \uart_drone.data_esr_3_LC_11_12_3 .C_ON=1'b0;
    defparam \uart_drone.data_esr_3_LC_11_12_3 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_esr_3_LC_11_12_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone.data_esr_3_LC_11_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47702),
            .lcout(uart_drone_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87048),
            .ce(N__47628),
            .sr(N__47616));
    defparam \uart_drone.data_esr_4_LC_11_12_4 .C_ON=1'b0;
    defparam \uart_drone.data_esr_4_LC_11_12_4 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_esr_4_LC_11_12_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone.data_esr_4_LC_11_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47687),
            .lcout(uart_drone_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87048),
            .ce(N__47628),
            .sr(N__47616));
    defparam \uart_drone.data_esr_5_LC_11_12_5 .C_ON=1'b0;
    defparam \uart_drone.data_esr_5_LC_11_12_5 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_esr_5_LC_11_12_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone.data_esr_5_LC_11_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47672),
            .lcout(uart_drone_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87048),
            .ce(N__47628),
            .sr(N__47616));
    defparam \uart_drone.data_esr_6_LC_11_12_6 .C_ON=1'b0;
    defparam \uart_drone.data_esr_6_LC_11_12_6 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_esr_6_LC_11_12_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone.data_esr_6_LC_11_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47657),
            .lcout(uart_drone_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87048),
            .ce(N__47628),
            .sr(N__47616));
    defparam \uart_drone.data_esr_7_LC_11_12_7 .C_ON=1'b0;
    defparam \uart_drone.data_esr_7_LC_11_12_7 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_esr_7_LC_11_12_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone.data_esr_7_LC_11_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47642),
            .lcout(uart_drone_data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87048),
            .ce(N__47628),
            .sr(N__47616));
    defparam \dron_frame_decoder_1.state_ns_0_i_a2_0_5_3_LC_11_13_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_ns_0_i_a2_0_5_3_LC_11_13_0 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_ns_0_i_a2_0_5_3_LC_11_13_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \dron_frame_decoder_1.state_ns_0_i_a2_0_5_3_LC_11_13_0  (
            .in0(N__58790),
            .in1(N__59049),
            .in2(N__58627),
            .in3(N__59274),
            .lcout(\dron_frame_decoder_1.N_230_5 ),
            .ltout(\dron_frame_decoder_1.N_230_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_ns_i_a2_2_0_a2_0_LC_11_13_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_ns_i_a2_2_0_a2_0_LC_11_13_1 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_ns_i_a2_2_0_a2_0_LC_11_13_1 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \dron_frame_decoder_1.state_ns_i_a2_2_0_a2_0_LC_11_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__47601),
            .in3(N__50929),
            .lcout(\dron_frame_decoder_1.N_224 ),
            .ltout(\dron_frame_decoder_1.N_224_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_RNO_0_0_LC_11_13_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNO_0_0_LC_11_13_2 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNO_0_0_LC_11_13_2 .LUT_INIT=16'b1111000010000000;
    LogicCell40 \dron_frame_decoder_1.state_RNO_0_0_LC_11_13_2  (
            .in0(N__47751),
            .in1(N__51000),
            .in2(N__47598),
            .in3(N__47772),
            .lcout(\dron_frame_decoder_1.N_198 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_ns_i_a2_1_1_0_LC_11_13_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_ns_i_a2_1_1_0_LC_11_13_3 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_ns_i_a2_1_1_0_LC_11_13_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \dron_frame_decoder_1.state_ns_i_a2_1_1_0_LC_11_13_3  (
            .in0(_gnd_net_),
            .in1(N__58966),
            .in2(_gnd_net_),
            .in3(N__59147),
            .lcout(),
            .ltout(\dron_frame_decoder_1.state_ns_i_a2_1_1Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_RNIN9KQ1_0_LC_11_13_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNIN9KQ1_0_LC_11_13_4 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNIN9KQ1_0_LC_11_13_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \dron_frame_decoder_1.state_RNIN9KQ1_0_LC_11_13_4  (
            .in0(N__58875),
            .in1(N__58697),
            .in2(N__47775),
            .in3(N__51015),
            .lcout(\dron_frame_decoder_1.N_220 ),
            .ltout(\dron_frame_decoder_1.N_220_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_1_LC_11_13_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_1_LC_11_13_5 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.state_1_LC_11_13_5 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \dron_frame_decoder_1.state_1_LC_11_13_5  (
            .in0(N__51042),
            .in1(N__47766),
            .in2(N__47760),
            .in3(N__51154),
            .lcout(\dron_frame_decoder_1.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87059),
            .ce(),
            .sr(N__79610));
    defparam \dron_frame_decoder_1.state_0_LC_11_13_6 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_0_LC_11_13_6 .SEQ_MODE=4'b1001;
    defparam \dron_frame_decoder_1.state_0_LC_11_13_6 .LUT_INIT=16'b0000000000001101;
    LogicCell40 \dron_frame_decoder_1.state_0_LC_11_13_6  (
            .in0(N__51155),
            .in1(N__51016),
            .in2(N__51027),
            .in3(N__47757),
            .lcout(\dron_frame_decoder_1.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87059),
            .ce(),
            .sr(N__79610));
    defparam \dron_frame_decoder_1.state_RNO_3_0_LC_11_13_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNO_3_0_LC_11_13_7 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNO_3_0_LC_11_13_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \dron_frame_decoder_1.state_RNO_3_0_LC_11_13_7  (
            .in0(N__58698),
            .in1(N__58967),
            .in2(N__59167),
            .in3(N__58876),
            .lcout(\dron_frame_decoder_1.state_ns_i_a2_0_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_RNI0TLI1_4_LC_11_14_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNI0TLI1_4_LC_11_14_0 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNI0TLI1_4_LC_11_14_0 .LUT_INIT=16'b1010101110101010;
    LogicCell40 \dron_frame_decoder_1.state_RNI0TLI1_4_LC_11_14_0  (
            .in0(N__79948),
            .in1(N__47745),
            .in2(N__47862),
            .in3(N__50992),
            .lcout(\dron_frame_decoder_1.N_740_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_RNI7Q6K_5_LC_11_14_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNI7Q6K_5_LC_11_14_1 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNI7Q6K_5_LC_11_14_1 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \dron_frame_decoder_1.state_RNI7Q6K_5_LC_11_14_1  (
            .in0(_gnd_net_),
            .in1(N__50928),
            .in2(_gnd_net_),
            .in3(N__47874),
            .lcout(\dron_frame_decoder_1.un1_sink_data_valid_5_i_0 ),
            .ltout(\dron_frame_decoder_1.un1_sink_data_valid_5_i_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_RNI3T3K1_7_LC_11_14_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNI3T3K1_7_LC_11_14_2 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNI3T3K1_7_LC_11_14_2 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \dron_frame_decoder_1.state_RNI3T3K1_7_LC_11_14_2  (
            .in0(N__51113),
            .in1(N__47850),
            .in2(N__47739),
            .in3(N__50991),
            .lcout(),
            .ltout(\dron_frame_decoder_1.state_RNI3T3K1Z0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_RNI0AAT1_7_LC_11_14_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNI0AAT1_7_LC_11_14_3 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNI0AAT1_7_LC_11_14_3 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \dron_frame_decoder_1.state_RNI0AAT1_7_LC_11_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__47736),
            .in3(N__79949),
            .lcout(\dron_frame_decoder_1.N_732_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_5_LC_11_14_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_5_LC_11_14_4 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.state_5_LC_11_14_4 .LUT_INIT=16'b1111111110100000;
    LogicCell40 \dron_frame_decoder_1.state_5_LC_11_14_4  (
            .in0(N__51168),
            .in1(_gnd_net_),
            .in2(N__47880),
            .in3(N__51183),
            .lcout(\dron_frame_decoder_1.stateZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87066),
            .ce(),
            .sr(N__79617));
    defparam \dron_frame_decoder_1.state_4_LC_11_14_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_4_LC_11_14_5 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.state_4_LC_11_14_5 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \dron_frame_decoder_1.state_4_LC_11_14_5  (
            .in0(N__50945),
            .in1(N__47876),
            .in2(N__47861),
            .in3(N__51167),
            .lcout(\dron_frame_decoder_1.stateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87066),
            .ce(),
            .sr(N__79617));
    defparam \uart_drone.data_rdy_LC_11_14_6 .C_ON=1'b0;
    defparam \uart_drone.data_rdy_LC_11_14_6 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_rdy_LC_11_14_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uart_drone.data_rdy_LC_11_14_6  (
            .in0(_gnd_net_),
            .in1(N__47982),
            .in2(_gnd_net_),
            .in3(N__47901),
            .lcout(uart_drone_data_rdy),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87066),
            .ce(),
            .sr(N__79617));
    defparam \dron_frame_decoder_1.state_RNI1H181_5_LC_11_14_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNI1H181_5_LC_11_14_7 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNI1H181_5_LC_11_14_7 .LUT_INIT=16'b1111111100001000;
    LogicCell40 \dron_frame_decoder_1.state_RNI1H181_5_LC_11_14_7  (
            .in0(N__50944),
            .in1(N__47875),
            .in2(N__47860),
            .in3(N__79950),
            .lcout(\dron_frame_decoder_1.N_716_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_RNI6P6K_4_LC_11_15_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNI6P6K_4_LC_11_15_0 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNI6P6K_4_LC_11_15_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \dron_frame_decoder_1.state_RNI6P6K_4_LC_11_15_0  (
            .in0(_gnd_net_),
            .in1(N__47849),
            .in2(_gnd_net_),
            .in3(N__50947),
            .lcout(\dron_frame_decoder_1.state_RNI6P6KZ0Z_4 ),
            .ltout(\dron_frame_decoder_1.state_RNI6P6KZ0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_RNI36DT_4_LC_11_15_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNI36DT_4_LC_11_15_1 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNI36DT_4_LC_11_15_1 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \dron_frame_decoder_1.state_RNI36DT_4_LC_11_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__47829),
            .in3(N__79936),
            .lcout(\dron_frame_decoder_1.N_724_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNI80O6_8_LC_11_15_3 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNI80O6_8_LC_11_15_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNI80O6_8_LC_11_15_3 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNI80O6_8_LC_11_15_3  (
            .in0(_gnd_net_),
            .in1(N__48547),
            .in2(_gnd_net_),
            .in3(N__49686),
            .lcout(\pid_front.N_2167_i ),
            .ltout(\pid_front.N_2167_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIGL6F_0_8_LC_11_15_4 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIGL6F_0_8_LC_11_15_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIGL6F_0_8_LC_11_15_4 .LUT_INIT=16'b0101101010010110;
    LogicCell40 \pid_front.error_p_reg_esr_RNIGL6F_0_8_LC_11_15_4  (
            .in0(N__48059),
            .in1(N__48041),
            .in2(N__47826),
            .in3(N__49731),
            .lcout(\pid_front.error_p_reg_esr_RNIGL6F_0Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_RNI4N6K_2_LC_11_15_6 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNI4N6K_2_LC_11_15_6 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNI4N6K_2_LC_11_15_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \dron_frame_decoder_1.state_RNI4N6K_2_LC_11_15_6  (
            .in0(_gnd_net_),
            .in1(N__47816),
            .in2(_gnd_net_),
            .in3(N__50946),
            .lcout(\dron_frame_decoder_1.state_RNI4N6KZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIPC5D1_7_LC_11_16_0 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIPC5D1_7_LC_11_16_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIPC5D1_7_LC_11_16_0 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_front.error_p_reg_esr_RNIPC5D1_7_LC_11_16_0  (
            .in0(N__48177),
            .in1(N__48183),
            .in2(_gnd_net_),
            .in3(N__55083),
            .lcout(\pid_front.error_p_reg_esr_RNIPC5D1Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIBG6F_7_LC_11_16_1 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIBG6F_7_LC_11_16_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIBG6F_7_LC_11_16_1 .LUT_INIT=16'b1111010101110001;
    LogicCell40 \pid_front.error_p_reg_esr_RNIBG6F_7_LC_11_16_1  (
            .in0(N__48129),
            .in1(N__48102),
            .in2(N__48123),
            .in3(N__49777),
            .lcout(\pid_front.error_p_reg_esr_RNIBG6FZ0Z_7 ),
            .ltout(\pid_front.error_p_reg_esr_RNIBG6FZ0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI5B9Q2_7_LC_11_16_2 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI5B9Q2_7_LC_11_16_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI5B9Q2_7_LC_11_16_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pid_front.error_p_reg_esr_RNI5B9Q2_7_LC_11_16_2  (
            .in0(N__48176),
            .in1(N__48168),
            .in2(N__48144),
            .in3(N__55082),
            .lcout(\pid_front.error_p_reg_esr_RNI5B9Q2Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNI6UN6_7_LC_11_16_4 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNI6UN6_7_LC_11_16_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNI6UN6_7_LC_11_16_4 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNI6UN6_7_LC_11_16_4  (
            .in0(_gnd_net_),
            .in1(N__48037),
            .in2(_gnd_net_),
            .in3(N__49728),
            .lcout(\pid_front.N_2161_i ),
            .ltout(\pid_front.N_2161_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIBG6F_0_7_LC_11_16_5 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIBG6F_0_7_LC_11_16_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIBG6F_0_7_LC_11_16_5 .LUT_INIT=16'b0101101010010110;
    LogicCell40 \pid_front.error_p_reg_esr_RNIBG6F_0_7_LC_11_16_5  (
            .in0(N__48119),
            .in1(N__48101),
            .in2(N__48087),
            .in3(N__49776),
            .lcout(\pid_front.error_p_reg_esr_RNIBG6F_0Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_7_LC_11_16_6 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_7_LC_11_16_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_7_LC_11_16_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_7_LC_11_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49730),
            .lcout(\pid_front.error_d_reg_prevZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87091),
            .ce(N__70427),
            .sr(N__70356));
    defparam \pid_front.error_p_reg_esr_RNIGL6F_8_LC_11_16_7 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIGL6F_8_LC_11_16_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIGL6F_8_LC_11_16_7 .LUT_INIT=16'b1000110011101111;
    LogicCell40 \pid_front.error_p_reg_esr_RNIGL6F_8_LC_11_16_7  (
            .in0(N__49729),
            .in1(N__48069),
            .in2(N__48042),
            .in3(N__48024),
            .lcout(\pid_front.error_p_reg_esr_RNIGL6FZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_xy_ki_3_rep2_esr_LC_11_17_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_ki_3_rep2_esr_LC_11_17_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_ki_3_rep2_esr_LC_11_17_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_xy_ki_3_rep2_esr_LC_11_17_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84019),
            .lcout(xy_ki_3_rep2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87107),
            .ce(N__78690),
            .sr(N__79641));
    defparam \Commands_frame_decoder.source_xy_ki_fast_esr_3_LC_11_17_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_ki_fast_esr_3_LC_11_17_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_ki_fast_esr_3_LC_11_17_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Commands_frame_decoder.source_xy_ki_fast_esr_3_LC_11_17_1  (
            .in0(N__84021),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(xy_ki_fast_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87107),
            .ce(N__78690),
            .sr(N__79641));
    defparam \Commands_frame_decoder.source_xy_ki_esr_3_LC_11_17_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_ki_esr_3_LC_11_17_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_ki_esr_3_LC_11_17_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_xy_ki_esr_3_LC_11_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84020),
            .lcout(xy_ki_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87107),
            .ce(N__78690),
            .sr(N__79641));
    defparam \Commands_frame_decoder.source_xy_ki_esr_2_LC_11_17_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_ki_esr_2_LC_11_17_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_ki_esr_2_LC_11_17_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_xy_ki_esr_2_LC_11_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__77547),
            .lcout(xy_ki_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87107),
            .ce(N__78690),
            .sr(N__79641));
    defparam \Commands_frame_decoder.source_xy_ki_esr_5_LC_11_17_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_ki_esr_5_LC_11_17_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_ki_esr_5_LC_11_17_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_xy_ki_esr_5_LC_11_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85209),
            .lcout(xy_ki_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87107),
            .ce(N__78690),
            .sr(N__79641));
    defparam \Commands_frame_decoder.source_xy_ki_esr_6_LC_11_17_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_ki_esr_6_LC_11_17_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_ki_esr_6_LC_11_17_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Commands_frame_decoder.source_xy_ki_esr_6_LC_11_17_5  (
            .in0(N__73646),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(xy_ki_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87107),
            .ce(N__78690),
            .sr(N__79641));
    defparam \Commands_frame_decoder.source_xy_ki_esr_7_LC_11_17_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_ki_esr_7_LC_11_17_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_ki_esr_7_LC_11_17_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_xy_ki_esr_7_LC_11_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85374),
            .lcout(xy_ki_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87107),
            .ce(N__78690),
            .sr(N__79641));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_10_LC_11_18_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_10_LC_11_18_0 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_10_LC_11_18_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_10_LC_11_18_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59063),
            .lcout(\dron_frame_decoder_1.drone_H_disp_side_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87121),
            .ce(N__48480),
            .sr(N__79649));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_11_LC_11_18_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_11_LC_11_18_1 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_11_LC_11_18_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_11_LC_11_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58982),
            .lcout(drone_H_disp_side_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87121),
            .ce(N__48480),
            .sr(N__79649));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_12_LC_11_18_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_12_LC_11_18_2 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_12_LC_11_18_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_12_LC_11_18_2  (
            .in0(N__58918),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(drone_H_disp_side_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87121),
            .ce(N__48480),
            .sr(N__79649));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_13_LC_11_18_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_13_LC_11_18_3 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_13_LC_11_18_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_13_LC_11_18_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58825),
            .lcout(drone_H_disp_side_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87121),
            .ce(N__48480),
            .sr(N__79649));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_14_LC_11_18_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_14_LC_11_18_4 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_14_LC_11_18_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_14_LC_11_18_4  (
            .in0(N__58725),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(drone_H_disp_side_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87121),
            .ce(N__48480),
            .sr(N__79649));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_15_LC_11_18_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_15_LC_11_18_5 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_15_LC_11_18_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_15_LC_11_18_5  (
            .in0(N__58634),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(drone_H_disp_side_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87121),
            .ce(N__48480),
            .sr(N__79649));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_8_LC_11_18_6 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_8_LC_11_18_6 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_8_LC_11_18_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_8_LC_11_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59286),
            .lcout(\dron_frame_decoder_1.drone_H_disp_side_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87121),
            .ce(N__48480),
            .sr(N__79649));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_9_LC_11_18_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_9_LC_11_18_7 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_9_LC_11_18_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_9_LC_11_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59182),
            .lcout(\dron_frame_decoder_1.drone_H_disp_side_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87121),
            .ce(N__48480),
            .sr(N__79649));
    defparam \pid_alt.error_i_acumm_5_LC_11_19_0 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_5_LC_11_19_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_5_LC_11_19_0 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \pid_alt.error_i_acumm_5_LC_11_19_0  (
            .in0(N__65396),
            .in1(N__48398),
            .in2(N__48468),
            .in3(N__48435),
            .lcout(\pid_alt.error_i_acummZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87136),
            .ce(),
            .sr(N__49359));
    defparam \pid_front.error_d_reg_prev_esr_RNIBTE61_0_21_LC_11_19_1 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIBTE61_0_21_LC_11_19_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIBTE61_0_21_LC_11_19_1 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIBTE61_0_21_LC_11_19_1  (
            .in0(N__48309),
            .in1(N__48581),
            .in2(_gnd_net_),
            .in3(N__87463),
            .lcout(\pid_front.error_d_reg_prev_esr_RNIBTE61_0Z0Z_21 ),
            .ltout(\pid_front.error_d_reg_prev_esr_RNIBTE61_0Z0Z_21_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIJVAC3_20_LC_11_19_2 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIJVAC3_20_LC_11_19_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIJVAC3_20_LC_11_19_2 .LUT_INIT=16'b1111110011000000;
    LogicCell40 \pid_front.error_p_reg_esr_RNIJVAC3_20_LC_11_19_2  (
            .in0(_gnd_net_),
            .in1(N__48350),
            .in2(N__48372),
            .in3(N__55724),
            .lcout(\pid_front.un1_pid_prereg_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI8QE61_20_LC_11_19_3 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI8QE61_20_LC_11_19_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI8QE61_20_LC_11_19_3 .LUT_INIT=16'b1101110101000100;
    LogicCell40 \pid_front.error_p_reg_esr_RNI8QE61_20_LC_11_19_3  (
            .in0(N__48594),
            .in1(N__48228),
            .in2(_gnd_net_),
            .in3(N__83643),
            .lcout(\pid_front.error_p_reg_esr_RNI8QE61Z0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIBTE61_21_LC_11_19_4 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIBTE61_21_LC_11_19_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIBTE61_21_LC_11_19_4 .LUT_INIT=16'b1010111100001010;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIBTE61_21_LC_11_19_4  (
            .in0(N__87464),
            .in1(_gnd_net_),
            .in2(N__48585),
            .in3(N__48310),
            .lcout(\pid_front.error_d_reg_prev_esr_RNIBTE61Z0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI8QE61_0_20_LC_11_19_5 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI8QE61_0_20_LC_11_19_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI8QE61_0_20_LC_11_19_5 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_front.error_p_reg_esr_RNI8QE61_0_20_LC_11_19_5  (
            .in0(N__48593),
            .in1(N__48227),
            .in2(_gnd_net_),
            .in3(N__83642),
            .lcout(\pid_front.error_p_reg_esr_RNI8QE61_0Z0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIOLN44_12_LC_11_19_6 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIOLN44_12_LC_11_19_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIOLN44_12_LC_11_19_6 .LUT_INIT=16'b0011000011001111;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIOLN44_12_LC_11_19_6  (
            .in0(_gnd_net_),
            .in1(N__49628),
            .in2(N__48672),
            .in3(N__48615),
            .lcout(\pid_front.error_d_reg_prev_esr_RNIOLN44Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIUO6U_0_12_LC_11_19_7 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIUO6U_0_12_LC_11_19_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIUO6U_0_12_LC_11_19_7 .LUT_INIT=16'b1011101110111011;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIUO6U_0_12_LC_11_19_7  (
            .in0(N__49629),
            .in1(N__48667),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.N_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_11_LC_11_20_0 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_11_LC_11_20_0 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_11_LC_11_20_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_front.error_d_reg_prev_esr_11_LC_11_20_0  (
            .in0(N__49181),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_d_reg_prevZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87154),
            .ce(N__70470),
            .sr(N__70351));
    defparam \pid_front.error_d_reg_prev_esr_14_LC_11_20_1 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_14_LC_11_20_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_14_LC_11_20_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_14_LC_11_20_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82775),
            .lcout(\pid_front.error_d_reg_prevZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87154),
            .ce(N__70470),
            .sr(N__70351));
    defparam \pid_front.error_d_reg_prev_esr_19_LC_11_20_2 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_19_LC_11_20_2 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_19_LC_11_20_2 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \pid_front.error_d_reg_prev_esr_19_LC_11_20_2  (
            .in0(_gnd_net_),
            .in1(N__87507),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_d_reg_prevZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87154),
            .ce(N__70470),
            .sr(N__70351));
    defparam \pid_front.error_d_reg_prev_esr_20_LC_11_20_3 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_20_LC_11_20_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_20_LC_11_20_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_20_LC_11_20_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__83641),
            .lcout(\pid_front.error_d_reg_prevZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87154),
            .ce(N__70470),
            .sr(N__70351));
    defparam \pid_front.error_d_reg_prev_esr_21_LC_11_20_4 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_21_LC_11_20_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_21_LC_11_20_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_21_LC_11_20_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__87465),
            .lcout(\pid_front.error_d_reg_prevZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87154),
            .ce(N__70470),
            .sr(N__70351));
    defparam \pid_front.error_d_reg_prev_esr_5_LC_11_20_5 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_5_LC_11_20_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_5_LC_11_20_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_front.error_d_reg_prev_esr_5_LC_11_20_5  (
            .in0(N__49019),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_d_reg_prevZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87154),
            .ce(N__70470),
            .sr(N__70351));
    defparam \pid_front.error_d_reg_prev_esr_8_LC_11_20_6 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_8_LC_11_20_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_8_LC_11_20_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_8_LC_11_20_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49689),
            .lcout(\pid_front.error_d_reg_prevZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87154),
            .ce(N__70470),
            .sr(N__70351));
    defparam \pid_front.error_d_reg_prev_fast_esr_12_LC_11_20_7 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_fast_esr_12_LC_11_20_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_fast_esr_12_LC_11_20_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_prev_fast_esr_12_LC_11_20_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49624),
            .lcout(\pid_front.error_d_reg_prev_fastZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87154),
            .ce(N__70470),
            .sr(N__70351));
    defparam \pid_front.error_d_reg_prev_esr_RNIUO6U_12_LC_11_21_0 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIUO6U_12_LC_11_21_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIUO6U_12_LC_11_21_0 .LUT_INIT=16'b1010111110101111;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIUO6U_12_LC_11_21_0  (
            .in0(N__49622),
            .in1(_gnd_net_),
            .in2(N__48658),
            .in3(_gnd_net_),
            .lcout(\pid_front.N_5_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIUO6U_2_12_LC_11_21_1 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIUO6U_2_12_LC_11_21_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIUO6U_2_12_LC_11_21_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIUO6U_2_12_LC_11_21_1  (
            .in0(_gnd_net_),
            .in1(N__48645),
            .in2(_gnd_net_),
            .in3(N__49621),
            .lcout(),
            .ltout(\pid_front.N_3_i_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIROQ33_12_LC_11_21_2 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIROQ33_12_LC_11_21_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIROQ33_12_LC_11_21_2 .LUT_INIT=16'b0000010100010111;
    LogicCell40 \pid_front.error_p_reg_esr_RNIROQ33_12_LC_11_21_2  (
            .in0(N__48971),
            .in1(N__49246),
            .in2(N__48912),
            .in3(N__48909),
            .lcout(\pid_front.N_3_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIETB61_13_LC_11_21_3 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIETB61_13_LC_11_21_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIETB61_13_LC_11_21_3 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_front.error_p_reg_esr_RNIETB61_13_LC_11_21_3  (
            .in0(N__48881),
            .in1(N__48814),
            .in2(_gnd_net_),
            .in3(N__48769),
            .lcout(),
            .ltout(\pid_front.N_2198_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIVTNC2_14_LC_11_21_4 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIVTNC2_14_LC_11_21_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIVTNC2_14_LC_11_21_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \pid_front.error_p_reg_esr_RNIVTNC2_14_LC_11_21_4  (
            .in0(N__54268),
            .in1(N__54291),
            .in2(N__48735),
            .in3(N__82769),
            .lcout(),
            .ltout(\pid_front.g0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI6D5L7_12_LC_11_21_5 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI6D5L7_12_LC_11_21_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI6D5L7_12_LC_11_21_5 .LUT_INIT=16'b0100101111010010;
    LogicCell40 \pid_front.error_p_reg_esr_RNI6D5L7_12_LC_11_21_5  (
            .in0(N__48732),
            .in1(N__48726),
            .in2(N__48720),
            .in3(N__48717),
            .lcout(),
            .ltout(\pid_front.error_p_reg_esr_RNI6D5L7Z0Z_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIIL0TE_12_LC_11_21_6 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIIL0TE_12_LC_11_21_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIIL0TE_12_LC_11_21_6 .LUT_INIT=16'b1001011001011010;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIIL0TE_12_LC_11_21_6  (
            .in0(N__55414),
            .in1(N__55460),
            .in2(N__48708),
            .in3(N__48705),
            .lcout(\pid_front.un1_pid_prereg_0_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_12_LC_11_21_7 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_12_LC_11_21_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_12_LC_11_21_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_12_LC_11_21_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49623),
            .lcout(\pid_front.error_d_reg_prevZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87169),
            .ce(N__70468),
            .sr(N__70349));
    defparam \pid_alt.error_i_acumm_esr_13_LC_11_22_0 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_esr_13_LC_11_22_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_esr_13_LC_11_22_0 .LUT_INIT=16'b1100110011011101;
    LogicCell40 \pid_alt.error_i_acumm_esr_13_LC_11_22_0  (
            .in0(N__49485),
            .in1(N__49443),
            .in2(_gnd_net_),
            .in3(N__49422),
            .lcout(\pid_alt.error_i_acummZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87184),
            .ce(N__49383),
            .sr(N__49358));
    defparam \pid_front.error_i_acumm_prereg_esr_RNI0V2N_28_LC_11_22_1 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_RNI0V2N_28_LC_11_22_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_acumm_prereg_esr_RNI0V2N_28_LC_11_22_1 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_RNI0V2N_28_LC_11_22_1  (
            .in0(N__60115),
            .in1(N__55497),
            .in2(_gnd_net_),
            .in3(N__79966),
            .lcout(\pid_front.error_i_acumm_3_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI0GC61_0_19_LC_11_22_4 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI0GC61_0_19_LC_11_22_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI0GC61_0_19_LC_11_22_4 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_front.error_p_reg_esr_RNI0GC61_0_19_LC_11_22_4  (
            .in0(N__49286),
            .in1(N__49298),
            .in2(_gnd_net_),
            .in3(N__87502),
            .lcout(\pid_front.error_p_reg_esr_RNI0GC61_0Z0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI0GC61_19_LC_11_22_5 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI0GC61_19_LC_11_22_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI0GC61_19_LC_11_22_5 .LUT_INIT=16'b1010111100001010;
    LogicCell40 \pid_front.error_p_reg_esr_RNI0GC61_19_LC_11_22_5  (
            .in0(N__87503),
            .in1(_gnd_net_),
            .in2(N__49302),
            .in3(N__49287),
            .lcout(\pid_front.error_p_reg_esr_RNI0GC61Z0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI8NB61_0_11_LC_11_22_6 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI8NB61_0_11_LC_11_22_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI8NB61_0_11_LC_11_22_6 .LUT_INIT=16'b1100000011001100;
    LogicCell40 \pid_front.error_p_reg_esr_RNI8NB61_0_11_LC_11_22_6  (
            .in0(_gnd_net_),
            .in1(N__49154),
            .in2(N__49136),
            .in3(N__49215),
            .lcout(\pid_front.un1_pid_prereg_135_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI8NB61_11_LC_11_22_7 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI8NB61_11_LC_11_22_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI8NB61_11_LC_11_22_7 .LUT_INIT=16'b1111010101010000;
    LogicCell40 \pid_front.error_p_reg_esr_RNI8NB61_11_LC_11_22_7  (
            .in0(N__49216),
            .in1(_gnd_net_),
            .in2(N__49167),
            .in3(N__49137),
            .lcout(\pid_front.g0_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_esr_4_LC_11_23_0 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_4_LC_11_23_0 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_4_LC_11_23_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_esr_4_LC_11_23_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49065),
            .lcout(\pid_front.error_d_regZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87197),
            .ce(N__86276),
            .sr(N__86009));
    defparam \pid_front.error_d_reg_esr_5_LC_11_23_1 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_5_LC_11_23_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_5_LC_11_23_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_esr_5_LC_11_23_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49035),
            .lcout(\pid_front.error_d_regZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87197),
            .ce(N__86276),
            .sr(N__86009));
    defparam \pid_front.error_d_reg_esr_6_LC_11_23_2 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_6_LC_11_23_2 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_6_LC_11_23_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_esr_6_LC_11_23_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48993),
            .lcout(\pid_front.error_d_regZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87197),
            .ce(N__86276),
            .sr(N__86009));
    defparam \pid_front.error_d_reg_esr_7_LC_11_23_3 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_7_LC_11_23_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_7_LC_11_23_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_esr_7_LC_11_23_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49752),
            .lcout(\pid_front.error_d_regZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87197),
            .ce(N__86276),
            .sr(N__86009));
    defparam \pid_front.error_d_reg_esr_8_LC_11_23_4 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_8_LC_11_23_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_8_LC_11_23_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_esr_8_LC_11_23_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49710),
            .lcout(\pid_front.error_d_regZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87197),
            .ce(N__86276),
            .sr(N__86009));
    defparam \pid_front.error_d_reg_esr_12_LC_11_23_5 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_12_LC_11_23_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_12_LC_11_23_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_esr_12_LC_11_23_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49652),
            .lcout(\pid_front.error_d_regZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87197),
            .ce(N__86276),
            .sr(N__86009));
    defparam \pid_front.error_p_reg_esr_0_LC_11_23_6 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_0_LC_11_23_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_0_LC_11_23_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_p_reg_esr_0_LC_11_23_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49569),
            .lcout(\pid_front.error_p_regZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87197),
            .ce(N__86276),
            .sr(N__86009));
    defparam \pid_front.error_p_reg_esr_10_LC_11_23_7 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_10_LC_11_23_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_10_LC_11_23_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_p_reg_esr_10_LC_11_23_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49527),
            .lcout(\pid_front.error_p_regZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87197),
            .ce(N__86276),
            .sr(N__86009));
    defparam \pid_front.error_i_acumm_prereg_esr_RNIMNV4_0_LC_11_24_0 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_RNIMNV4_0_LC_11_24_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_acumm_prereg_esr_RNIMNV4_0_LC_11_24_0 .LUT_INIT=16'b1111111000000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_RNIMNV4_0_LC_11_24_0  (
            .in0(N__52214),
            .in1(N__56117),
            .in2(N__52199),
            .in3(N__52181),
            .lcout(\pid_front.un10lt9_1 ),
            .ltout(\pid_front.un10lt9_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_prereg_esr_RNI9SN8_4_LC_11_24_1 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_RNI9SN8_4_LC_11_24_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_acumm_prereg_esr_RNI9SN8_4_LC_11_24_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_RNI9SN8_4_LC_11_24_1  (
            .in0(N__52091),
            .in1(N__52468),
            .in2(N__49491),
            .in3(N__52108),
            .lcout(),
            .ltout(\pid_front.un10lt9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_prereg_esr_RNI5AGC_7_LC_11_24_2 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_RNI5AGC_7_LC_11_24_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_acumm_prereg_esr_RNI5AGC_7_LC_11_24_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_RNI5AGC_7_LC_11_24_2  (
            .in0(N__52046),
            .in1(N__52013),
            .in2(N__49488),
            .in3(N__52523),
            .lcout(\pid_front.un10lt11_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_prereg_esr_RNI9SN8_0_4_LC_11_24_3 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_RNI9SN8_0_4_LC_11_24_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_acumm_prereg_esr_RNI9SN8_0_4_LC_11_24_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_RNI9SN8_0_4_LC_11_24_3  (
            .in0(N__52090),
            .in1(N__52109),
            .in2(N__49863),
            .in3(N__52469),
            .lcout(),
            .ltout(\pid_front.error_i_acumm16lt9_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_prereg_esr_RNIV9S71_12_LC_11_24_4 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_RNIV9S71_12_LC_11_24_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_acumm_prereg_esr_RNIV9S71_12_LC_11_24_4 .LUT_INIT=16'b0010001000101010;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_RNIV9S71_12_LC_11_24_4  (
            .in0(N__52751),
            .in1(N__51093),
            .in2(N__49854),
            .in3(N__49851),
            .lcout(\pid_front.error_i_acumm_prereg_esr_RNIV9S71Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_prereg_esr_RNISDO3_7_LC_11_24_5 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_RNISDO3_7_LC_11_24_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_acumm_prereg_esr_RNISDO3_7_LC_11_24_5 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_RNISDO3_7_LC_11_24_5  (
            .in0(N__52012),
            .in1(N__52522),
            .in2(_gnd_net_),
            .in3(N__52045),
            .lcout(\pid_front.error_i_acumm_prereg_esr_RNISDO3Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_prereg_esr_3_LC_11_24_6 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_3_LC_11_24_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_3_LC_11_24_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_3_LC_11_24_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54717),
            .lcout(\pid_front.error_i_acumm16lto3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87216),
            .ce(N__56081),
            .sr(N__79686));
    defparam \pid_front.error_i_acumm_prereg_esr_1_LC_11_24_7 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_1_LC_11_24_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_1_LC_11_24_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_1_LC_11_24_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54808),
            .lcout(\pid_front.error_i_acumm_preregZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87216),
            .ce(N__56081),
            .sr(N__79686));
    defparam \pid_front.error_p_reg_esr_1_LC_11_25_0 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_1_LC_11_25_0 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_esr_1_LC_11_25_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_p_reg_esr_1_LC_11_25_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49845),
            .lcout(\pid_front.error_p_regZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87229),
            .ce(N__86292),
            .sr(N__86007));
    defparam \pid_front.error_p_reg_esr_RNIL1E8_1_LC_11_25_1 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIL1E8_1_LC_11_25_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIL1E8_1_LC_11_25_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_front.error_p_reg_esr_RNIL1E8_1_LC_11_25_1  (
            .in0(N__52566),
            .in1(N__52279),
            .in2(_gnd_net_),
            .in3(N__52590),
            .lcout(),
            .ltout(\pid_front.un1_pid_prereg_9_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIMRLT_0_LC_11_25_2 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIMRLT_0_LC_11_25_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIMRLT_0_LC_11_25_2 .LUT_INIT=16'b0000111111000011;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIMRLT_0_LC_11_25_2  (
            .in0(N__54809),
            .in1(N__52233),
            .in2(N__49830),
            .in3(N__52254),
            .lcout(\pid_front.error_d_reg_prev_esr_RNIMRLTZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_esr_1_LC_11_25_3 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_1_LC_11_25_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_1_LC_11_25_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_esr_1_LC_11_25_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49812),
            .lcout(\pid_front.error_d_regZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87229),
            .ce(N__86292),
            .sr(N__86007));
    defparam \pid_front.error_d_reg_prev_esr_RNIAHDK_0_LC_11_25_4 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIAHDK_0_LC_11_25_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIAHDK_0_LC_11_25_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIAHDK_0_LC_11_25_4  (
            .in0(N__54845),
            .in1(N__52232),
            .in2(_gnd_net_),
            .in3(N__52253),
            .lcout(\pid_front.error_d_reg_prev_esr_RNIAHDKZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_prereg_esr_RNIRU7I_10_LC_11_25_5 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_RNIRU7I_10_LC_11_25_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_acumm_prereg_esr_RNIRU7I_10_LC_11_25_5 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_RNIRU7I_10_LC_11_25_5  (
            .in0(N__52138),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52447),
            .lcout(),
            .ltout(\pid_front.error_i_acumm_prereg_esr_RNIRU7IZ0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_prereg_esr_RNI0I2H5_12_LC_11_25_6 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_RNI0I2H5_12_LC_11_25_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_acumm_prereg_esr_RNI0I2H5_12_LC_11_25_6 .LUT_INIT=16'b0111011101110011;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_RNI0I2H5_12_LC_11_25_6  (
            .in0(N__52747),
            .in1(N__49869),
            .in2(N__49896),
            .in3(N__49893),
            .lcout(\pid_front.error_i_acumm_prereg_esr_RNI0I2H5Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_esr_0_LC_11_25_7 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_0_LC_11_25_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_0_LC_11_25_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_esr_0_LC_11_25_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49887),
            .lcout(\pid_front.error_d_regZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87229),
            .ce(N__86292),
            .sr(N__86007));
    defparam \pid_front.error_i_acumm_prereg_esr_RNI8II41_18_LC_11_26_0 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_RNI8II41_18_LC_11_26_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_acumm_prereg_esr_RNI8II41_18_LC_11_26_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_RNI8II41_18_LC_11_26_0  (
            .in0(N__52494),
            .in1(N__49991),
            .in2(N__52541),
            .in3(N__49980),
            .lcout(),
            .ltout(\pid_front.un10lto27_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_prereg_esr_RNI18694_0_14_LC_11_26_1 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_RNI18694_0_14_LC_11_26_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_acumm_prereg_esr_RNI18694_0_14_LC_11_26_1 .LUT_INIT=16'b1000000010000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_RNI18694_0_14_LC_11_26_1  (
            .in0(N__52653),
            .in1(N__49998),
            .in2(N__49872),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_i_acumm_prereg_esr_RNI18694_0Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_prereg_esr_18_LC_11_26_3 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_18_LC_11_26_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_18_LC_11_26_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_18_LC_11_26_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55320),
            .lcout(\pid_front.error_i_acumm_preregZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87243),
            .ce(N__56076),
            .sr(N__79692));
    defparam \pid_front.error_i_acumm_prereg_esr_19_LC_11_26_4 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_19_LC_11_26_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_19_LC_11_26_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_19_LC_11_26_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55286),
            .lcout(\pid_front.error_i_acumm_preregZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87243),
            .ce(N__56076),
            .sr(N__79692));
    defparam \pid_front.error_i_acumm_prereg_esr_14_LC_11_26_5 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_14_LC_11_26_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_14_LC_11_26_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_14_LC_11_26_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55418),
            .lcout(\pid_front.error_i_acumm_preregZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87243),
            .ce(N__56076),
            .sr(N__79692));
    defparam \pid_front.error_i_acumm_prereg_esr_15_LC_11_26_7 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_15_LC_11_26_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_15_LC_11_26_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_15_LC_11_26_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55380),
            .lcout(\pid_front.error_i_acumm_preregZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87243),
            .ce(N__56076),
            .sr(N__79692));
    defparam \pid_front.error_i_acumm_prereg_esr_RNIAIG41_14_LC_11_27_0 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_RNIAIG41_14_LC_11_27_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_acumm_prereg_esr_RNIAIG41_14_LC_11_27_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_RNIAIG41_14_LC_11_27_0  (
            .in0(N__52502),
            .in1(N__49955),
            .in2(N__56154),
            .in3(N__49967),
            .lcout(\pid_front.un10lto27_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_prereg_esr_RNI8II41_0_18_LC_11_27_2 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_RNI8II41_0_18_LC_11_27_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_acumm_prereg_esr_RNI8II41_0_18_LC_11_27_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_RNI8II41_0_18_LC_11_27_2  (
            .in0(N__52490),
            .in1(N__49992),
            .in2(N__52542),
            .in3(N__49979),
            .lcout(\pid_front.error_i_acumm16lto27_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_prereg_esr_RNIAIG41_0_14_LC_11_27_5 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_RNIAIG41_0_14_LC_11_27_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_acumm_prereg_esr_RNIAIG41_0_14_LC_11_27_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_RNIAIG41_0_14_LC_11_27_5  (
            .in0(N__49968),
            .in1(N__56153),
            .in2(N__49959),
            .in3(N__52503),
            .lcout(\pid_front.error_i_acumm16lto27_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIQGK21_1_LC_12_1_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIQGK21_1_LC_12_1_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIQGK21_1_LC_12_1_1 .LUT_INIT=16'b1100110001101100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIQGK21_1_LC_12_1_1  (
            .in0(N__60938),
            .in1(N__63682),
            .in2(N__61064),
            .in3(N__64265),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNISIK21_3_LC_12_1_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNISIK21_3_LC_12_1_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNISIK21_3_LC_12_1_3 .LUT_INIT=16'b1100110001101100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNISIK21_3_LC_12_1_3  (
            .in0(N__60939),
            .in1(N__53231),
            .in2(N__61065),
            .in3(N__64266),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIC3MT_10_LC_12_1_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIC3MT_10_LC_12_1_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIC3MT_10_LC_12_1_5 .LUT_INIT=16'b1010101001101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIC3MT_10_LC_12_1_5  (
            .in0(N__60579),
            .in1(N__63381),
            .in2(N__64602),
            .in3(N__64267),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNILU3P_0_LC_12_1_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNILU3P_0_LC_12_1_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNILU3P_0_LC_12_1_7 .LUT_INIT=16'b1111000001111000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNILU3P_0_LC_12_1_7  (
            .in0(N__53586),
            .in1(N__57270),
            .in2(N__63644),
            .in3(N__64264),
            .lcout(\ppm_encoder_1.N_257_i_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_esr_RNI6C0M1_14_LC_12_2_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_esr_RNI6C0M1_14_LC_12_2_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_esr_RNI6C0M1_14_LC_12_2_0 .LUT_INIT=16'b0000110001011101;
    LogicCell40 \ppm_encoder_1.elevator_esr_RNI6C0M1_14_LC_12_2_0  (
            .in0(N__49926),
            .in1(N__63354),
            .in2(N__49914),
            .in3(N__63588),
            .lcout(\ppm_encoder_1.elevator_esr_RNI6C0M1Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m6_i_0_LC_12_2_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m6_i_0_LC_12_2_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m6_i_0_LC_12_2_1 .LUT_INIT=16'b1111101001011010;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m6_i_0_LC_12_2_1  (
            .in0(N__63589),
            .in1(_gnd_net_),
            .in2(N__63404),
            .in3(N__64548),
            .lcout(\ppm_encoder_1.N_56 ),
            .ltout(\ppm_encoder_1.N_56_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_LC_12_2_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_LC_12_2_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_LC_12_2_2 .LUT_INIT=16'b0010001000000011;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_2_LC_12_2_2  (
            .in0(N__63389),
            .in1(N__79984),
            .in2(N__50058),
            .in3(N__64233),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__86972),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIV9203_6_LC_12_2_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIV9203_6_LC_12_2_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIV9203_6_LC_12_2_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIV9203_6_LC_12_2_3  (
            .in0(N__50230),
            .in1(N__56928),
            .in2(N__61690),
            .in3(N__57331),
            .lcout(\ppm_encoder_1.init_pulses_RNIV9203Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNIB7481_3_LC_12_2_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNIB7481_3_LC_12_2_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNIB7481_3_LC_12_2_4 .LUT_INIT=16'b1111111100111001;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_RNIB7481_3_LC_12_2_4  (
            .in0(N__63858),
            .in1(N__63359),
            .in2(N__64585),
            .in3(N__64232),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_RNIB7481Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIE5MT_12_LC_12_2_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIE5MT_12_LC_12_2_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIE5MT_12_LC_12_2_5 .LUT_INIT=16'b1011111101000000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIE5MT_12_LC_12_2_5  (
            .in0(N__64231),
            .in1(N__64547),
            .in2(N__63403),
            .in3(N__50444),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIH8MT_15_LC_12_2_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIH8MT_15_LC_12_2_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIH8MT_15_LC_12_2_6 .LUT_INIT=16'b1111000001111000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIH8MT_15_LC_12_2_6  (
            .in0(N__64546),
            .in1(N__63355),
            .in2(N__64673),
            .in3(N__64230),
            .lcout(\ppm_encoder_1.N_254_i_i ),
            .ltout(\ppm_encoder_1.N_254_i_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNI82G01_15_LC_12_2_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI82G01_15_LC_12_2_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI82G01_15_LC_12_2_7 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI82G01_15_LC_12_2_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__50025),
            .in3(N__64669),
            .lcout(\ppm_encoder_1.init_pulses_RNI82G01Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIDAHV_13_LC_12_3_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIDAHV_13_LC_12_3_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIDAHV_13_LC_12_3_0 .LUT_INIT=16'b1001110011001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIDAHV_13_LC_12_3_0  (
            .in0(N__64147),
            .in1(N__53368),
            .in2(N__61057),
            .in3(N__60908),
            .lcout(\ppm_encoder_1.N_268_i_i ),
            .ltout(\ppm_encoder_1.N_268_i_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNITIRP2_13_LC_12_3_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNITIRP2_13_LC_12_3_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNITIRP2_13_LC_12_3_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNITIRP2_13_LC_12_3_1  (
            .in0(N__56938),
            .in1(N__53372),
            .in2(N__50010),
            .in3(N__57332),
            .lcout(\ppm_encoder_1.init_pulses_RNITIRP2Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNITLK21_6_LC_12_3_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNITLK21_6_LC_12_3_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNITLK21_6_LC_12_3_3 .LUT_INIT=16'b1111000001111000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNITLK21_6_LC_12_3_3  (
            .in0(N__63793),
            .in1(N__57711),
            .in2(N__61694),
            .in3(N__64146),
            .lcout(\ppm_encoder_1.N_262_i_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNILN0E1_6_LC_12_3_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNILN0E1_6_LC_12_3_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNILN0E1_6_LC_12_3_4 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \ppm_encoder_1.throttle_RNILN0E1_6_LC_12_3_4  (
            .in0(N__58005),
            .in1(N__61730),
            .in2(N__61770),
            .in3(N__57182),
            .lcout(\ppm_encoder_1.un2_throttle_iv_0_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.rudder_RNIRRSI2_6_LC_12_3_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_RNIRRSI2_6_LC_12_3_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.rudder_RNIRRSI2_6_LC_12_3_5 .LUT_INIT=16'b1111111111101100;
    LogicCell40 \ppm_encoder_1.rudder_RNIRRSI2_6_LC_12_3_5  (
            .in0(N__63794),
            .in1(N__57758),
            .in2(N__57794),
            .in3(N__57052),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_1_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIS2VR4_6_LC_12_3_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIS2VR4_6_LC_12_3_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIS2VR4_6_LC_12_3_6 .LUT_INIT=16'b0011011011001001;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIS2VR4_6_LC_12_3_6  (
            .in0(N__50253),
            .in1(N__56937),
            .in2(N__50247),
            .in3(N__61689),
            .lcout(),
            .ltout(\ppm_encoder_1.un1_init_pulses_0_axb_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIPOJU5_6_LC_12_3_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIPOJU5_6_LC_12_3_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIPOJU5_6_LC_12_3_7 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIPOJU5_6_LC_12_3_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__50244),
            .in3(N__50229),
            .lcout(\ppm_encoder_1.init_pulses_RNIPOJU5Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.rudder_esr_RNI0Q0I2_4_LC_12_4_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_esr_RNI0Q0I2_4_LC_12_4_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.rudder_esr_RNI0Q0I2_4_LC_12_4_0 .LUT_INIT=16'b1111111111101100;
    LogicCell40 \ppm_encoder_1.rudder_esr_RNI0Q0I2_4_LC_12_4_0  (
            .in0(N__63757),
            .in1(N__50199),
            .in2(N__59753),
            .in3(N__57010),
            .lcout(\ppm_encoder_1.un2_throttle_iv_0_2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.rudder_esr_4_LC_12_4_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_esr_4_LC_12_4_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.rudder_esr_4_LC_12_4_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.rudder_esr_4_LC_12_4_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50184),
            .lcout(\ppm_encoder_1.rudderZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__86979),
            .ce(N__50160),
            .sr(N__79567));
    defparam \ppm_encoder_1.init_pulses_RNIK58G4_10_LC_12_5_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIK58G4_10_LC_12_5_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIK58G4_10_LC_12_5_0 .LUT_INIT=16'b0101101001101001;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIK58G4_10_LC_12_5_0  (
            .in0(N__56939),
            .in1(N__53349),
            .in2(N__60578),
            .in3(N__50376),
            .lcout(),
            .ltout(\ppm_encoder_1.un1_init_pulses_0_axb_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIUCPF5_10_LC_12_5_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIUCPF5_10_LC_12_5_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIUCPF5_10_LC_12_5_1 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIUCPF5_10_LC_12_5_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__50085),
            .in3(N__50360),
            .lcout(\ppm_encoder_1.init_pulses_RNIUCPF5Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.rudder_RNI22TI2_9_LC_12_5_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_RNI22TI2_9_LC_12_5_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.rudder_RNI22TI2_9_LC_12_5_2 .LUT_INIT=16'b1111111111101100;
    LogicCell40 \ppm_encoder_1.rudder_RNI22TI2_9_LC_12_5_2  (
            .in0(N__60881),
            .in1(N__50070),
            .in2(N__61808),
            .in3(N__57026),
            .lcout(\ppm_encoder_1.un2_throttle_iv_0_2_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.rudder_RNII8J92_10_LC_12_5_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_RNII8J92_10_LC_12_5_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.rudder_RNII8J92_10_LC_12_5_3 .LUT_INIT=16'b1111111111101010;
    LogicCell40 \ppm_encoder_1.rudder_RNII8J92_10_LC_12_5_3  (
            .in0(N__57027),
            .in1(N__60879),
            .in2(N__60798),
            .in3(N__50382),
            .lcout(\ppm_encoder_1.un2_throttle_iv_0_2_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIA7HV_10_LC_12_5_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIA7HV_10_LC_12_5_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIA7HV_10_LC_12_5_4 .LUT_INIT=16'b1111000001111000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIA7HV_10_LC_12_5_4  (
            .in0(N__60880),
            .in1(N__60985),
            .in2(N__60577),
            .in3(N__64272),
            .lcout(\ppm_encoder_1.N_255_i_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_LC_12_5_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_LC_12_5_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_LC_12_5_5 .LUT_INIT=16'b1111111111011000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_0_LC_12_5_5  (
            .in0(N__64273),
            .in1(N__61565),
            .in2(N__57449),
            .in3(N__79990),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__86985),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_LC_12_5_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_LC_12_5_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_LC_12_5_6 .LUT_INIT=16'b0000101000000110;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_LC_12_5_6  (
            .in0(N__52795),
            .in1(N__61566),
            .in2(N__80001),
            .in3(N__64274),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__86985),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNIDA6O_6_LC_12_5_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNIDA6O_6_LC_12_5_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNIDA6O_6_LC_12_5_7 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \ppm_encoder_1.elevator_RNIDA6O_6_LC_12_5_7  (
            .in0(N__50555),
            .in1(N__52794),
            .in2(_gnd_net_),
            .in3(N__52912),
            .lcout(\ppm_encoder_1.elevator_RNIDA6OZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_1_LC_12_6_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_1_LC_12_6_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_1_LC_12_6_0 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_1_LC_12_6_0  (
            .in0(N__68887),
            .in1(N__57904),
            .in2(N__53256),
            .in3(N__68660),
            .lcout(\ppm_encoder_1.pulses2count_9_0_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_1_LC_12_6_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_1_LC_12_6_1 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.aileron_1_LC_12_6_1 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \ppm_encoder_1.aileron_1_LC_12_6_1  (
            .in0(N__53255),
            .in1(N__50349),
            .in2(N__65189),
            .in3(N__53832),
            .lcout(\ppm_encoder_1.aileronZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__86993),
            .ce(),
            .sr(N__79578));
    defparam \ppm_encoder_1.throttle_1_LC_12_6_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_1_LC_12_6_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_1_LC_12_6_2 .LUT_INIT=16'b1010010111001100;
    LogicCell40 \ppm_encoder_1.throttle_1_LC_12_6_2  (
            .in0(N__50337),
            .in1(N__57905),
            .in2(N__50325),
            .in3(N__65099),
            .lcout(\ppm_encoder_1.throttleZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__86993),
            .ce(),
            .sr(N__79578));
    defparam \ppm_encoder_1.elevator_7_LC_12_6_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_7_LC_12_6_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.elevator_7_LC_12_6_5 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.elevator_7_LC_12_6_5  (
            .in0(N__50298),
            .in1(N__50283),
            .in2(N__65190),
            .in3(N__50262),
            .lcout(\ppm_encoder_1.elevatorZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__86993),
            .ce(),
            .sr(N__79578));
    defparam \ppm_encoder_1.elevator_RNIEB6O_7_LC_12_6_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNIEB6O_7_LC_12_6_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNIEB6O_7_LC_12_6_6 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \ppm_encoder_1.elevator_RNIEB6O_7_LC_12_6_6  (
            .in0(N__50261),
            .in1(N__52796),
            .in2(_gnd_net_),
            .in3(N__52913),
            .lcout(\ppm_encoder_1.elevator_RNIEB6OZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_11_LC_12_7_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_11_LC_12_7_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_11_LC_12_7_1 .LUT_INIT=16'b0101111100010011;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_11_LC_12_7_1  (
            .in0(N__57377),
            .in1(N__52634),
            .in2(N__68675),
            .in3(N__63584),
            .lcout(),
            .ltout(\ppm_encoder_1.pulses2count_9_0_3_1_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_11_LC_12_7_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_11_LC_12_7_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_11_LC_12_7_2 .LUT_INIT=16'b1110111110101111;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_11_LC_12_7_2  (
            .in0(N__53592),
            .in1(N__64443),
            .in2(N__50505),
            .in3(N__53063),
            .lcout(\ppm_encoder_1.pulses2count_9_0_3_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNIRHGE_13_LC_12_7_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNIRHGE_13_LC_12_7_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNIRHGE_13_LC_12_7_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \ppm_encoder_1.elevator_RNIRHGE_13_LC_12_7_5  (
            .in0(N__50502),
            .in1(N__52817),
            .in2(_gnd_net_),
            .in3(N__52934),
            .lcout(\ppm_encoder_1.elevator_RNIRHGEZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_12_LC_12_7_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_12_LC_12_7_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_12_LC_12_7_6 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_12_LC_12_7_6  (
            .in0(N__60924),
            .in1(N__63864),
            .in2(_gnd_net_),
            .in3(N__50484),
            .lcout(),
            .ltout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_12_LC_12_7_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_12_LC_12_7_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_12_LC_12_7_7 .LUT_INIT=16'b1111101111110011;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_12_LC_12_7_7  (
            .in0(N__64442),
            .in1(N__50457),
            .in2(N__50451),
            .in3(N__50448),
            .lcout(\ppm_encoder_1.pulses2count_9_0_3_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_LC_12_8_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_LC_12_8_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_LC_12_8_0 .LUT_INIT=16'b0000101100000001;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_LC_12_8_0  (
            .in0(N__64292),
            .in1(N__57416),
            .in2(N__79999),
            .in3(N__63756),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87007),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.PPM_STATE_RNISH5F_1_LC_12_8_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_RNISH5F_1_LC_12_8_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.PPM_STATE_RNISH5F_1_LC_12_8_1 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \ppm_encoder_1.PPM_STATE_RNISH5F_1_LC_12_8_1  (
            .in0(_gnd_net_),
            .in1(N__79937),
            .in2(_gnd_net_),
            .in3(N__64291),
            .lcout(\ppm_encoder_1.N_295_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.data_Aux_RNO_0_1_LC_12_8_2 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_RNO_0_1_LC_12_8_2 .SEQ_MODE=4'b0000;
    defparam \uart_drone.data_Aux_RNO_0_1_LC_12_8_2 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \uart_drone.data_Aux_RNO_0_1_LC_12_8_2  (
            .in0(N__62133),
            .in1(N__62190),
            .in2(_gnd_net_),
            .in3(N__62070),
            .lcout(\uart_drone.data_Auxce_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.data_Aux_RNO_0_2_LC_12_8_3 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_RNO_0_2_LC_12_8_3 .SEQ_MODE=4'b0000;
    defparam \uart_drone.data_Aux_RNO_0_2_LC_12_8_3 .LUT_INIT=16'b0000010100000000;
    LogicCell40 \uart_drone.data_Aux_RNO_0_2_LC_12_8_3  (
            .in0(N__62071),
            .in1(_gnd_net_),
            .in2(N__62205),
            .in3(N__62134),
            .lcout(\uart_drone.data_Auxce_0_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.data_Aux_RNO_0_4_LC_12_8_5 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_RNO_0_4_LC_12_8_5 .SEQ_MODE=4'b0000;
    defparam \uart_drone.data_Aux_RNO_0_4_LC_12_8_5 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \uart_drone.data_Aux_RNO_0_4_LC_12_8_5  (
            .in0(N__62072),
            .in1(_gnd_net_),
            .in2(N__62206),
            .in3(N__62135),
            .lcout(\uart_drone.data_Auxce_0_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.data_Aux_RNO_0_5_LC_12_8_6 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_RNO_0_5_LC_12_8_6 .SEQ_MODE=4'b0000;
    defparam \uart_drone.data_Aux_RNO_0_5_LC_12_8_6 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \uart_drone.data_Aux_RNO_0_5_LC_12_8_6  (
            .in0(N__62136),
            .in1(N__62197),
            .in2(_gnd_net_),
            .in3(N__62073),
            .lcout(\uart_drone.data_Auxce_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.data_Aux_RNO_0_6_LC_12_8_7 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_RNO_0_6_LC_12_8_7 .SEQ_MODE=4'b0000;
    defparam \uart_drone.data_Aux_RNO_0_6_LC_12_8_7 .LUT_INIT=16'b0101000000000000;
    LogicCell40 \uart_drone.data_Aux_RNO_0_6_LC_12_8_7  (
            .in0(N__62074),
            .in1(_gnd_net_),
            .in2(N__62207),
            .in3(N__62137),
            .lcout(\uart_drone.data_Auxce_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_3_LC_12_9_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_3_LC_12_9_0 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.aileron_3_LC_12_9_0 .LUT_INIT=16'b1101100001110010;
    LogicCell40 \ppm_encoder_1.aileron_3_LC_12_9_0  (
            .in0(N__65183),
            .in1(N__53870),
            .in2(N__68170),
            .in3(N__50604),
            .lcout(\ppm_encoder_1.aileronZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87015),
            .ce(),
            .sr(N__79596));
    defparam \ppm_encoder_1.aileron_12_LC_12_9_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_12_LC_12_9_3 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.aileron_12_LC_12_9_3 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \ppm_encoder_1.aileron_12_LC_12_9_3  (
            .in0(N__58338),
            .in1(N__50598),
            .in2(N__60371),
            .in3(N__65182),
            .lcout(\ppm_encoder_1.aileronZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87015),
            .ce(),
            .sr(N__79596));
    defparam \ppm_encoder_1.elevator_6_LC_12_9_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_6_LC_12_9_5 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.elevator_6_LC_12_9_5 .LUT_INIT=16'b1001100111110000;
    LogicCell40 \ppm_encoder_1.elevator_6_LC_12_9_5  (
            .in0(N__50592),
            .in1(N__50580),
            .in2(N__50556),
            .in3(N__65188),
            .lcout(\ppm_encoder_1.elevatorZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87015),
            .ce(),
            .sr(N__79596));
    defparam \ppm_encoder_1.aileron_6_LC_12_9_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_6_LC_12_9_6 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.aileron_6_LC_12_9_6 .LUT_INIT=16'b1001111110010000;
    LogicCell40 \ppm_encoder_1.aileron_6_LC_12_9_6  (
            .in0(N__50538),
            .in1(N__58202),
            .in2(N__65271),
            .in3(N__61723),
            .lcout(\ppm_encoder_1.aileronZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87015),
            .ce(),
            .sr(N__79596));
    defparam \ppm_encoder_1.aileron_7_LC_12_9_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_7_LC_12_9_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.aileron_7_LC_12_9_7 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \ppm_encoder_1.aileron_7_LC_12_9_7  (
            .in0(N__50532),
            .in1(N__53510),
            .in2(N__53679),
            .in3(N__65187),
            .lcout(\ppm_encoder_1.aileronZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87015),
            .ce(),
            .sr(N__79596));
    defparam \uart_drone.bit_Count_1_LC_12_10_2 .C_ON=1'b0;
    defparam \uart_drone.bit_Count_1_LC_12_10_2 .SEQ_MODE=4'b1000;
    defparam \uart_drone.bit_Count_1_LC_12_10_2 .LUT_INIT=16'b0001010001010000;
    LogicCell40 \uart_drone.bit_Count_1_LC_12_10_2  (
            .in0(N__50873),
            .in1(N__62084),
            .in2(N__62141),
            .in3(N__50526),
            .lcout(\uart_drone.bit_CountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87021),
            .ce(),
            .sr(N__79602));
    defparam \uart_drone.bit_Count_2_LC_12_10_5 .C_ON=1'b0;
    defparam \uart_drone.bit_Count_2_LC_12_10_5 .SEQ_MODE=4'b1000;
    defparam \uart_drone.bit_Count_2_LC_12_10_5 .LUT_INIT=16'b0000000001101010;
    LogicCell40 \uart_drone.bit_Count_2_LC_12_10_5  (
            .in0(N__62185),
            .in1(N__62130),
            .in2(N__50886),
            .in3(N__50874),
            .lcout(\uart_drone.bit_CountZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87021),
            .ce(),
            .sr(N__79602));
    defparam \uart_drone.timer_Count_RNIU8TV1_3_LC_12_10_7 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_RNIU8TV1_3_LC_12_10_7 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNIU8TV1_3_LC_12_10_7 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uart_drone.timer_Count_RNIU8TV1_3_LC_12_10_7  (
            .in0(N__50858),
            .in1(N__50838),
            .in2(_gnd_net_),
            .in3(N__50787),
            .lcout(\uart_drone.N_144_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_xy_kp_0_e_0_4_LC_12_11_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_kp_0_e_0_4_LC_12_11_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_kp_0_e_0_4_LC_12_11_5 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_xy_kp_0_e_0_4_LC_12_11_5  (
            .in0(_gnd_net_),
            .in1(N__85198),
            .in2(_gnd_net_),
            .in3(N__86173),
            .lcout(xy_kp_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87030),
            .ce(N__82675),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_xy_kp_e_0_5_LC_12_11_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_kp_e_0_5_LC_12_11_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_kp_e_0_5_LC_12_11_6 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Commands_frame_decoder.source_xy_kp_e_0_5_LC_12_11_6  (
            .in0(N__86174),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73650),
            .lcout(xy_kp_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87030),
            .ce(N__82675),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_14_LC_12_12_0 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_14_LC_12_12_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_14_LC_12_12_0 .LUT_INIT=16'b0011101011001010;
    LogicCell40 \pid_side.pid_prereg_14_LC_12_12_0  (
            .in0(N__72685),
            .in1(N__81930),
            .in2(N__59859),
            .in3(N__69459),
            .lcout(\pid_side.pid_preregZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87040),
            .ce(),
            .sr(N__79611));
    defparam \pid_side.state_RNIL5IF_0_LC_12_12_2 .C_ON=1'b0;
    defparam \pid_side.state_RNIL5IF_0_LC_12_12_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.state_RNIL5IF_0_LC_12_12_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \pid_side.state_RNIL5IF_0_LC_12_12_2  (
            .in0(_gnd_net_),
            .in1(N__59835),
            .in2(_gnd_net_),
            .in3(N__79917),
            .lcout(\pid_side.state_RNIL5IFZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.state_1_LC_12_12_3 .C_ON=1'b0;
    defparam \pid_side.state_1_LC_12_12_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.state_1_LC_12_12_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.state_1_LC_12_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59848),
            .lcout(\pid_side.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87040),
            .ce(),
            .sr(N__79611));
    defparam \pid_alt.state_0_LC_12_12_4 .C_ON=1'b0;
    defparam \pid_alt.state_0_LC_12_12_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.state_0_LC_12_12_4 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \pid_alt.state_0_LC_12_12_4  (
            .in0(N__56018),
            .in1(N__59920),
            .in2(_gnd_net_),
            .in3(N__65347),
            .lcout(\pid_alt.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87040),
            .ce(),
            .sr(N__79611));
    defparam \pid_alt.state_1_LC_12_12_5 .C_ON=1'b0;
    defparam \pid_alt.state_1_LC_12_12_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.state_1_LC_12_12_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.state_1_LC_12_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56019),
            .lcout(\pid_alt.N_72_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87040),
            .ce(),
            .sr(N__79611));
    defparam \dron_frame_decoder_1.state_RNO_0_3_LC_12_13_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNO_0_3_LC_12_13_0 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNO_0_3_LC_12_13_0 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \dron_frame_decoder_1.state_RNO_0_3_LC_12_13_0  (
            .in0(N__50942),
            .in1(N__58968),
            .in2(N__58738),
            .in3(N__59166),
            .lcout(),
            .ltout(\dron_frame_decoder_1.state_ns_0_i_a2_0_2_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_3_LC_12_13_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_3_LC_12_13_1 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.state_3_LC_12_13_1 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \dron_frame_decoder_1.state_3_LC_12_13_1  (
            .in0(N__51073),
            .in1(N__51048),
            .in2(N__51081),
            .in3(N__51156),
            .lcout(\dron_frame_decoder_1.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87049),
            .ce(),
            .sr(N__79618));
    defparam \dron_frame_decoder_1.state_RNO_1_3_LC_12_13_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNO_1_3_LC_12_13_2 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNO_1_3_LC_12_13_2 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \dron_frame_decoder_1.state_RNO_1_3_LC_12_13_2  (
            .in0(N__58877),
            .in1(N__51054),
            .in2(_gnd_net_),
            .in3(N__51041),
            .lcout(\dron_frame_decoder_1.state_ns_0_i_a2_0_3_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_6_LC_12_13_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_6_LC_12_13_3 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.state_6_LC_12_13_3 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \dron_frame_decoder_1.state_6_LC_12_13_3  (
            .in0(N__50993),
            .in1(N__50943),
            .in2(N__51117),
            .in3(N__51157),
            .lcout(\dron_frame_decoder_1.stateZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87049),
            .ce(),
            .sr(N__79618));
    defparam \dron_frame_decoder_1.state_RNO_1_0_LC_12_13_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNO_1_0_LC_12_13_4 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNO_1_0_LC_12_13_4 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \dron_frame_decoder_1.state_RNO_1_0_LC_12_13_4  (
            .in0(N__51018),
            .in1(N__51040),
            .in2(N__50994),
            .in3(N__50935),
            .lcout(\dron_frame_decoder_1.N_200 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_RNO_2_0_LC_12_13_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNO_2_0_LC_12_13_5 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNO_2_0_LC_12_13_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \dron_frame_decoder_1.state_RNO_2_0_LC_12_13_5  (
            .in0(_gnd_net_),
            .in1(N__50986),
            .in2(_gnd_net_),
            .in3(N__51017),
            .lcout(\dron_frame_decoder_1.state_ns_i_a2_0_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_data_valid_LC_12_13_6 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_data_valid_LC_12_13_6 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_data_valid_LC_12_13_6 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \dron_frame_decoder_1.source_data_valid_LC_12_13_6  (
            .in0(N__50990),
            .in1(N__50936),
            .in2(_gnd_net_),
            .in3(N__59908),
            .lcout(debug_CH1_0A_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87049),
            .ce(),
            .sr(N__79618));
    defparam \pid_alt.state_RNIFCSD1_0_LC_12_13_7 .C_ON=1'b0;
    defparam \pid_alt.state_RNIFCSD1_0_LC_12_13_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.state_RNIFCSD1_0_LC_12_13_7 .LUT_INIT=16'b1111111100000010;
    LogicCell40 \pid_alt.state_RNIFCSD1_0_LC_12_13_7  (
            .in0(N__59907),
            .in1(N__65340),
            .in2(N__56020),
            .in3(N__79918),
            .lcout(\pid_alt.state_RNIFCSD1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.state_RNIVIRQ_0_LC_12_14_0 .C_ON=1'b0;
    defparam \pid_front.state_RNIVIRQ_0_LC_12_14_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.state_RNIVIRQ_0_LC_12_14_0 .LUT_INIT=16'b1111111100000010;
    LogicCell40 \pid_front.state_RNIVIRQ_0_LC_12_14_0  (
            .in0(N__59916),
            .in1(N__60195),
            .in2(N__60093),
            .in3(N__79919),
            .lcout(\pid_front.state_RNIVIRQZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNID18S_4_LC_12_14_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNID18S_4_LC_12_14_5 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNID18S_4_LC_12_14_5 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \Commands_frame_decoder.state_RNID18S_4_LC_12_14_5  (
            .in0(N__79921),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51339),
            .lcout(\Commands_frame_decoder.source_CH3data_1_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.state_RNI4FBH2_0_LC_12_14_7 .C_ON=1'b0;
    defparam \pid_side.state_RNI4FBH2_0_LC_12_14_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.state_RNI4FBH2_0_LC_12_14_7 .LUT_INIT=16'b1010111011111110;
    LogicCell40 \pid_side.state_RNI4FBH2_0_LC_12_14_7  (
            .in0(N__79920),
            .in1(N__59802),
            .in2(N__72637),
            .in3(N__59844),
            .lcout(\pid_side.error_i_acumm_1_sqmuxa_1_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_xy_kp_e_0_0_LC_12_15_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_kp_e_0_0_LC_12_15_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_kp_e_0_0_LC_12_15_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_xy_kp_e_0_0_LC_12_15_0  (
            .in0(_gnd_net_),
            .in1(N__83807),
            .in2(_gnd_net_),
            .in3(N__86161),
            .lcout(xy_kp_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87067),
            .ce(N__82688),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_xy_kp_e_0_2_LC_12_15_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_kp_e_0_2_LC_12_15_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_kp_e_0_2_LC_12_15_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_xy_kp_e_0_2_LC_12_15_2  (
            .in0(_gnd_net_),
            .in1(N__77585),
            .in2(_gnd_net_),
            .in3(N__86162),
            .lcout(xy_kp_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87067),
            .ce(N__82688),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_xy_kp_e_0_3_LC_12_15_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_kp_e_0_3_LC_12_15_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_kp_e_0_3_LC_12_15_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Commands_frame_decoder.source_xy_kp_e_0_3_LC_12_15_3  (
            .in0(N__86163),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84002),
            .lcout(xy_kp_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87067),
            .ce(N__82688),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_xy_kp_e_0_6_LC_12_15_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_kp_e_0_6_LC_12_15_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_kp_e_0_6_LC_12_15_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_xy_kp_e_0_6_LC_12_15_6  (
            .in0(_gnd_net_),
            .in1(N__85380),
            .in2(_gnd_net_),
            .in3(N__86164),
            .lcout(xy_kp_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87067),
            .ce(N__82688),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_RNI14DT_2_LC_12_15_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNI14DT_2_LC_12_15_7 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNI14DT_2_LC_12_15_7 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \dron_frame_decoder_1.state_RNI14DT_2_LC_12_15_7  (
            .in0(N__51179),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79959),
            .lcout(\dron_frame_decoder_1.N_708_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_7_LC_12_16_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_7_LC_12_16_0 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.state_7_LC_12_16_0 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \dron_frame_decoder_1.state_7_LC_12_16_0  (
            .in0(N__51166),
            .in1(N__51123),
            .in2(_gnd_net_),
            .in3(N__51112),
            .lcout(\dron_frame_decoder_1.stateZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87078),
            .ce(),
            .sr(N__79642));
    defparam \pid_front.error_i_acumm_prereg_esr_RNIRU7I_0_10_LC_12_16_1 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_RNIRU7I_0_10_LC_12_16_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_acumm_prereg_esr_RNIRU7I_0_10_LC_12_16_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_RNIRU7I_0_10_LC_12_16_1  (
            .in0(_gnd_net_),
            .in1(N__52455),
            .in2(_gnd_net_),
            .in3(N__52152),
            .lcout(\pid_front.error_i_acumm_prereg_esr_RNIRU7I_0Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.state_RNIFM151_0_LC_12_16_2 .C_ON=1'b0;
    defparam \pid_front.state_RNIFM151_0_LC_12_16_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.state_RNIFM151_0_LC_12_16_2 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \pid_front.state_RNIFM151_0_LC_12_16_2  (
            .in0(N__56094),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70362),
            .lcout(\pid_front.N_764_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.state_RNIM14N_0_LC_12_16_3 .C_ON=1'b0;
    defparam \pid_front.state_RNIM14N_0_LC_12_16_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.state_RNIM14N_0_LC_12_16_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \pid_front.state_RNIM14N_0_LC_12_16_3  (
            .in0(_gnd_net_),
            .in1(N__86148),
            .in2(_gnd_net_),
            .in3(N__56093),
            .lcout(\pid_front.state_RNIM14NZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.state_RNISV141_0_LC_12_16_4 .C_ON=1'b0;
    defparam \pid_front.state_RNISV141_0_LC_12_16_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.state_RNISV141_0_LC_12_16_4 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \pid_front.state_RNISV141_0_LC_12_16_4  (
            .in0(N__86150),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51405),
            .lcout(\pid_front.N_789_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNITU3P4_10_LC_12_16_5 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNITU3P4_10_LC_12_16_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNITU3P4_10_LC_12_16_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNITU3P4_10_LC_12_16_5  (
            .in0(_gnd_net_),
            .in1(N__78870),
            .in2(_gnd_net_),
            .in3(N__78903),
            .lcout(\pid_side.error_d_reg_prev_esr_RNITU3P4Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIUREI_7_LC_12_16_6 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIUREI_7_LC_12_16_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIUREI_7_LC_12_16_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIUREI_7_LC_12_16_6  (
            .in0(_gnd_net_),
            .in1(N__54027),
            .in2(_gnd_net_),
            .in3(N__81233),
            .lcout(\pid_side.N_2368_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.state_RNIIIOO_0_LC_12_16_7 .C_ON=1'b0;
    defparam \pid_side.state_RNIIIOO_0_LC_12_16_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.state_RNIIIOO_0_LC_12_16_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \pid_side.state_RNIIIOO_0_LC_12_16_7  (
            .in0(N__69908),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__86149),
            .lcout(\pid_side.state_RNIIIOOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI3I672_2_LC_12_17_0 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI3I672_2_LC_12_17_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI3I672_2_LC_12_17_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_front.error_p_reg_esr_RNI3I672_2_LC_12_17_0  (
            .in0(N__51381),
            .in1(N__54715),
            .in2(N__52308),
            .in3(N__51347),
            .lcout(\pid_front.error_p_reg_esr_RNI3I672Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIO4E8_2_LC_12_17_1 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIO4E8_2_LC_12_17_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIO4E8_2_LC_12_17_1 .LUT_INIT=16'b1000100011101110;
    LogicCell40 \pid_front.error_p_reg_esr_RNIO4E8_2_LC_12_17_1  (
            .in0(N__85421),
            .in1(N__51681),
            .in2(_gnd_net_),
            .in3(N__51660),
            .lcout(\pid_front.error_p_reg_esr_RNIO4E8Z0Z_2 ),
            .ltout(\pid_front.error_p_reg_esr_RNIO4E8Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI2VEV_2_LC_12_17_2 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI2VEV_2_LC_12_17_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI2VEV_2_LC_12_17_2 .LUT_INIT=16'b1111110011000000;
    LogicCell40 \pid_front.error_p_reg_esr_RNI2VEV_2_LC_12_17_2  (
            .in0(_gnd_net_),
            .in1(N__51348),
            .in2(N__51375),
            .in3(N__54716),
            .lcout(\pid_front.error_p_reg_esr_RNI2VEVZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIR7E8_0_3_LC_12_17_3 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIR7E8_0_3_LC_12_17_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIR7E8_0_3_LC_12_17_3 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_front.error_p_reg_esr_RNIR7E8_0_3_LC_12_17_3  (
            .in0(N__51650),
            .in1(N__51632),
            .in2(_gnd_net_),
            .in3(N__71218),
            .lcout(\pid_front.error_p_reg_esr_RNIR7E8_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_2_LC_12_17_4 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_2_LC_12_17_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_2_LC_12_17_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_2_LC_12_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85422),
            .lcout(\pid_front.error_d_reg_prevZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87092),
            .ce(N__70428),
            .sr(N__70352));
    defparam \pid_front.error_p_reg_esr_RNIO4E8_0_2_LC_12_17_5 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIO4E8_0_2_LC_12_17_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIO4E8_0_2_LC_12_17_5 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_front.error_p_reg_esr_RNIO4E8_0_2_LC_12_17_5  (
            .in0(N__85420),
            .in1(N__51680),
            .in2(_gnd_net_),
            .in3(N__51659),
            .lcout(\pid_front.error_p_reg_esr_RNIO4E8_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_3_LC_12_17_6 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_3_LC_12_17_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_3_LC_12_17_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_front.error_d_reg_prev_esr_3_LC_12_17_6  (
            .in0(N__71220),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_d_reg_prevZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87092),
            .ce(N__70428),
            .sr(N__70352));
    defparam \pid_front.error_p_reg_esr_RNIR7E8_3_LC_12_17_7 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIR7E8_3_LC_12_17_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIR7E8_3_LC_12_17_7 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_front.error_p_reg_esr_RNIR7E8_3_LC_12_17_7  (
            .in0(N__51651),
            .in1(N__51633),
            .in2(_gnd_net_),
            .in3(N__71219),
            .lcout(\pid_front.error_p_reg_esr_RNIR7E8Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNISPHM_15_LC_12_18_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNISPHM_15_LC_12_18_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNISPHM_15_LC_12_18_0 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNISPHM_15_LC_12_18_0  (
            .in0(N__51609),
            .in1(N__51509),
            .in2(_gnd_net_),
            .in3(N__51554),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNISPHMZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_15_LC_12_18_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_15_LC_12_18_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_15_LC_12_18_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_15_LC_12_18_1  (
            .in0(N__51555),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87108),
            .ce(N__51472),
            .sr(N__79657));
    defparam \pid_front.error_axb_7_LC_12_18_3 .C_ON=1'b0;
    defparam \pid_front.error_axb_7_LC_12_18_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_axb_7_LC_12_18_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_front.error_axb_7_LC_12_18_3  (
            .in0(_gnd_net_),
            .in1(N__54480),
            .in2(_gnd_net_),
            .in3(N__54462),
            .lcout(\pid_front.error_axbZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNI3C23_12_LC_12_18_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNI3C23_12_LC_12_18_4 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNI3C23_12_LC_12_18_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_RNI3C23_12_LC_12_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54506),
            .lcout(drone_H_disp_front_i_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_1_0_c_RNIAGTB1_LC_12_18_6 .C_ON=1'b0;
    defparam \pid_front.error_cry_1_0_c_RNIAGTB1_LC_12_18_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_1_0_c_RNIAGTB1_LC_12_18_6 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \pid_front.error_cry_1_0_c_RNIAGTB1_LC_12_18_6  (
            .in0(N__78213),
            .in1(N__67739),
            .in2(_gnd_net_),
            .in3(N__67669),
            .lcout(\pid_front.N_51_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNI8SE96_12_LC_12_18_7 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNI8SE96_12_LC_12_18_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNI8SE96_12_LC_12_18_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNI8SE96_12_LC_12_18_7  (
            .in0(N__55459),
            .in1(N__51927),
            .in2(_gnd_net_),
            .in3(N__51891),
            .lcout(\pid_front.error_d_reg_prev_esr_RNI8SE96Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNITCC61_0_18_LC_12_19_0 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNITCC61_0_18_LC_12_19_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNITCC61_0_18_LC_12_19_0 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_front.error_p_reg_esr_RNITCC61_0_18_LC_12_19_0  (
            .in0(N__87539),
            .in1(N__70202),
            .in2(_gnd_net_),
            .in3(N__70515),
            .lcout(\pid_front.error_p_reg_esr_RNITCC61_0Z0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_17_LC_12_19_1 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_17_LC_12_19_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_17_LC_12_19_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_17_LC_12_19_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__87579),
            .lcout(\pid_front.error_d_reg_prevZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87122),
            .ce(N__70467),
            .sr(N__70350));
    defparam \pid_front.error_p_reg_esr_RNIQ9C61_17_LC_12_19_2 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIQ9C61_17_LC_12_19_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIQ9C61_17_LC_12_19_2 .LUT_INIT=16'b1010111100001010;
    LogicCell40 \pid_front.error_p_reg_esr_RNIQ9C61_17_LC_12_19_2  (
            .in0(N__87578),
            .in1(_gnd_net_),
            .in2(N__51750),
            .in3(N__51768),
            .lcout(\pid_front.error_p_reg_esr_RNIQ9C61Z0Z_17 ),
            .ltout(\pid_front.error_p_reg_esr_RNIQ9C61Z0Z_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI3F9B3_17_LC_12_19_3 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI3F9B3_17_LC_12_19_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI3F9B3_17_LC_12_19_3 .LUT_INIT=16'b1111101010100000;
    LogicCell40 \pid_front.error_p_reg_esr_RNI3F9B3_17_LC_12_19_3  (
            .in0(N__55319),
            .in1(_gnd_net_),
            .in2(N__51846),
            .in3(N__51836),
            .lcout(\pid_front.un1_pid_prereg_0_6 ),
            .ltout(\pid_front.un1_pid_prereg_0_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNICS5DD_16_LC_12_19_4 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNICS5DD_16_LC_12_19_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNICS5DD_16_LC_12_19_4 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \pid_front.error_p_reg_esr_RNICS5DD_16_LC_12_19_4  (
            .in0(N__51822),
            .in1(N__51801),
            .in2(N__51780),
            .in3(N__51692),
            .lcout(\pid_front.error_p_reg_esr_RNICS5DDZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIQ9C61_0_17_LC_12_19_5 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIQ9C61_0_17_LC_12_19_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIQ9C61_0_17_LC_12_19_5 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_front.error_p_reg_esr_RNIQ9C61_0_17_LC_12_19_5  (
            .in0(N__51767),
            .in1(N__51746),
            .in2(_gnd_net_),
            .in3(N__87577),
            .lcout(\pid_front.error_p_reg_esr_RNIQ9C61_0Z0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIBOAB3_0_18_LC_12_19_6 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIBOAB3_0_18_LC_12_19_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIBOAB3_0_18_LC_12_19_6 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pid_front.error_p_reg_esr_RNIBOAB3_0_18_LC_12_19_6  (
            .in0(N__70535),
            .in1(_gnd_net_),
            .in2(N__51719),
            .in3(N__55282),
            .lcout(\pid_front.un1_pid_prereg_0_7 ),
            .ltout(\pid_front.un1_pid_prereg_0_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIE7KM6_17_LC_12_19_7 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIE7KM6_17_LC_12_19_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIE7KM6_17_LC_12_19_7 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \pid_front.error_p_reg_esr_RNIE7KM6_17_LC_12_19_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__51969),
            .in3(N__51962),
            .lcout(\pid_front.error_p_reg_esr_RNIE7KM6Z0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_CH3data_esr_0_LC_12_20_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH3data_esr_0_LC_12_20_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH3data_esr_0_LC_12_20_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Commands_frame_decoder.source_CH3data_esr_0_LC_12_20_0  (
            .in0(N__83835),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(front_command_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87137),
            .ce(N__51939),
            .sr(N__79672));
    defparam \Commands_frame_decoder.source_CH3data_esr_1_LC_12_20_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH3data_esr_1_LC_12_20_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH3data_esr_1_LC_12_20_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH3data_esr_1_LC_12_20_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84209),
            .lcout(front_command_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87137),
            .ce(N__51939),
            .sr(N__79672));
    defparam \Commands_frame_decoder.source_CH3data_esr_2_LC_12_20_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH3data_esr_2_LC_12_20_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH3data_esr_2_LC_12_20_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH3data_esr_2_LC_12_20_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__77578),
            .lcout(front_command_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87137),
            .ce(N__51939),
            .sr(N__79672));
    defparam \Commands_frame_decoder.source_CH3data_esr_3_LC_12_20_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH3data_esr_3_LC_12_20_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH3data_esr_3_LC_12_20_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH3data_esr_3_LC_12_20_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84029),
            .lcout(front_command_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87137),
            .ce(N__51939),
            .sr(N__79672));
    defparam \Commands_frame_decoder.source_CH3data_esr_4_LC_12_20_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH3data_esr_4_LC_12_20_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH3data_esr_4_LC_12_20_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH3data_esr_4_LC_12_20_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85041),
            .lcout(front_command_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87137),
            .ce(N__51939),
            .sr(N__79672));
    defparam \Commands_frame_decoder.source_CH3data_esr_5_LC_12_20_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH3data_esr_5_LC_12_20_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH3data_esr_5_LC_12_20_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH3data_esr_5_LC_12_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85210),
            .lcout(front_command_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87137),
            .ce(N__51939),
            .sr(N__79672));
    defparam \Commands_frame_decoder.source_CH3data_esr_6_LC_12_20_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH3data_esr_6_LC_12_20_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH3data_esr_6_LC_12_20_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH3data_esr_6_LC_12_20_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73655),
            .lcout(front_command_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87137),
            .ce(N__51939),
            .sr(N__79672));
    defparam \Commands_frame_decoder.source_CH3data_ess_7_LC_12_20_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH3data_ess_7_LC_12_20_7 .SEQ_MODE=4'b1001;
    defparam \Commands_frame_decoder.source_CH3data_ess_7_LC_12_20_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Commands_frame_decoder.source_CH3data_ess_7_LC_12_20_7  (
            .in0(N__85400),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(front_command_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87137),
            .ce(N__51939),
            .sr(N__79672));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_10_LC_12_21_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_10_LC_12_21_0 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_10_LC_12_21_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_10_LC_12_21_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59105),
            .lcout(\dron_frame_decoder_1.drone_H_disp_front_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87155),
            .ce(N__51990),
            .sr(N__79678));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_11_LC_12_21_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_11_LC_12_21_1 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_11_LC_12_21_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_11_LC_12_21_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59024),
            .lcout(drone_H_disp_front_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87155),
            .ce(N__51990),
            .sr(N__79678));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_12_LC_12_21_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_12_LC_12_21_2 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_12_LC_12_21_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_12_LC_12_21_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58928),
            .lcout(drone_H_disp_front_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87155),
            .ce(N__51990),
            .sr(N__79678));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_13_LC_12_21_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_13_LC_12_21_3 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_13_LC_12_21_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_13_LC_12_21_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58842),
            .lcout(drone_H_disp_front_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87155),
            .ce(N__51990),
            .sr(N__79678));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_14_LC_12_21_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_14_LC_12_21_4 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_14_LC_12_21_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_14_LC_12_21_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58752),
            .lcout(drone_H_disp_front_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87155),
            .ce(N__51990),
            .sr(N__79678));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_15_LC_12_21_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_15_LC_12_21_5 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_15_LC_12_21_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_15_LC_12_21_5  (
            .in0(N__58659),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(drone_H_disp_front_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87155),
            .ce(N__51990),
            .sr(N__79678));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_8_LC_12_21_6 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_8_LC_12_21_6 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_8_LC_12_21_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_8_LC_12_21_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59334),
            .lcout(\dron_frame_decoder_1.drone_H_disp_front_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87155),
            .ce(N__51990),
            .sr(N__79678));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_9_LC_12_21_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_9_LC_12_21_7 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_9_LC_12_21_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_9_LC_12_21_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59195),
            .lcout(\dron_frame_decoder_1.drone_H_disp_front_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87155),
            .ce(N__51990),
            .sr(N__79678));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNIOBV3_8_LC_12_22_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNIOBV3_8_LC_12_22_0 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNIOBV3_8_LC_12_22_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_RNIOBV3_8_LC_12_22_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51975),
            .lcout(drone_H_disp_front_i_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.state_RNI26LH_0_LC_12_22_1 .C_ON=1'b0;
    defparam \pid_front.state_RNI26LH_0_LC_12_22_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.state_RNI26LH_0_LC_12_22_1 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \pid_front.state_RNI26LH_0_LC_12_22_1  (
            .in0(N__60081),
            .in1(N__59950),
            .in2(_gnd_net_),
            .in3(N__60197),
            .lcout(\pid_front.state_ns_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNI4D23_13_LC_12_22_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNI4D23_13_LC_12_22_2 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNI4D23_13_LC_12_22_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_RNI4D23_13_LC_12_22_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54893),
            .lcout(drone_H_disp_front_i_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNI1A23_10_LC_12_22_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNI1A23_10_LC_12_22_3 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNI1A23_10_LC_12_22_3 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_RNI1A23_10_LC_12_22_3  (
            .in0(_gnd_net_),
            .in1(N__52071),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(drone_H_disp_front_i_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_0_c_RNIBQAV_LC_12_22_4 .C_ON=1'b0;
    defparam \pid_front.error_cry_0_c_RNIBQAV_LC_12_22_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_0_c_RNIBQAV_LC_12_22_4 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \pid_front.error_cry_0_c_RNIBQAV_LC_12_22_4  (
            .in0(N__78243),
            .in1(N__77166),
            .in2(_gnd_net_),
            .in3(N__77119),
            .lcout(\pid_front.N_3 ),
            .ltout(\pid_front.N_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_0_c_RNIGBBP1_LC_12_22_5 .C_ON=1'b0;
    defparam \pid_front.error_cry_0_c_RNIGBBP1_LC_12_22_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_0_c_RNIGBBP1_LC_12_22_5 .LUT_INIT=16'b0100011100000011;
    LogicCell40 \pid_front.error_cry_0_c_RNIGBBP1_LC_12_22_5  (
            .in0(N__78403),
            .in1(N__77874),
            .in2(N__52065),
            .in3(N__77262),
            .lcout(\pid_front.m2_0_03_3_i_0 ),
            .ltout(\pid_front.m2_0_03_3_i_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_0_6_LC_12_22_6 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_0_6_LC_12_22_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_0_6_LC_12_22_6 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_0_6_LC_12_22_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__52062),
            .in3(N__77386),
            .lcout(\pid_front.N_55_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNIPCV3_9_LC_12_22_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNIPCV3_9_LC_12_22_7 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNIPCV3_9_LC_12_22_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_RNIPCV3_9_LC_12_22_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52059),
            .lcout(drone_H_disp_front_i_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_12_LC_12_23_0 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_12_LC_12_23_0 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_12_LC_12_23_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \pid_front.error_i_acumm_12_LC_12_23_0  (
            .in0(N__52029),
            .in1(N__52392),
            .in2(_gnd_net_),
            .in3(N__52752),
            .lcout(\pid_front.error_i_acummZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87185),
            .ce(N__60006),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_7_LC_12_23_1 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_7_LC_12_23_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_7_LC_12_23_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \pid_front.error_i_acumm_7_LC_12_23_1  (
            .in0(N__52395),
            .in1(N__52030),
            .in2(_gnd_net_),
            .in3(N__52053),
            .lcout(\pid_front.error_i_acummZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87185),
            .ce(N__60006),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_8_LC_12_23_2 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_8_LC_12_23_2 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_8_LC_12_23_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \pid_front.error_i_acumm_8_LC_12_23_2  (
            .in0(N__52031),
            .in1(N__52396),
            .in2(_gnd_net_),
            .in3(N__52524),
            .lcout(\pid_front.error_i_acummZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87185),
            .ce(N__60006),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_9_LC_12_23_3 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_9_LC_12_23_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_9_LC_12_23_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \pid_front.error_i_acumm_9_LC_12_23_3  (
            .in0(N__52397),
            .in1(N__52032),
            .in2(_gnd_net_),
            .in3(N__52017),
            .lcout(\pid_front.error_i_acummZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87185),
            .ce(N__60006),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_1_LC_12_23_4 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_1_LC_12_23_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_1_LC_12_23_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \pid_front.error_i_acumm_1_LC_12_23_4  (
            .in0(_gnd_net_),
            .in1(N__52393),
            .in2(_gnd_net_),
            .in3(N__52215),
            .lcout(\pid_front.error_i_acummZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87185),
            .ce(N__60006),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_2_LC_12_23_5 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_2_LC_12_23_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_2_LC_12_23_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \pid_front.error_i_acumm_2_LC_12_23_5  (
            .in0(N__52394),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52203),
            .lcout(\pid_front.error_i_acummZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87185),
            .ce(N__60006),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_0_LC_12_23_6 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_0_LC_12_23_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_0_LC_12_23_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \pid_front.error_i_acumm_0_LC_12_23_6  (
            .in0(_gnd_net_),
            .in1(N__52391),
            .in2(_gnd_net_),
            .in3(N__56118),
            .lcout(\pid_front.error_i_acummZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87185),
            .ce(N__60006),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_3_LC_12_23_7 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_3_LC_12_23_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_3_LC_12_23_7 .LUT_INIT=16'b1000100011011000;
    LogicCell40 \pid_front.error_i_acumm_3_LC_12_23_7  (
            .in0(N__52398),
            .in1(N__52182),
            .in2(N__60129),
            .in3(N__66045),
            .lcout(\pid_front.error_i_acummZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87185),
            .ce(N__60006),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_prereg_esr_RNI38E36_28_LC_12_24_0 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_RNI38E36_28_LC_12_24_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_acumm_prereg_esr_RNI38E36_28_LC_12_24_0 .LUT_INIT=16'b0000000011110010;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_RNI38E36_28_LC_12_24_0  (
            .in0(N__52704),
            .in1(N__52170),
            .in2(N__55496),
            .in3(N__66039),
            .lcout(\pid_front.error_i_acumm_2_sqmuxa_1 ),
            .ltout(\pid_front.error_i_acumm_2_sqmuxa_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_prereg_esr_RNI6CD2C_28_LC_12_24_1 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_RNI6CD2C_28_LC_12_24_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_acumm_prereg_esr_RNI6CD2C_28_LC_12_24_1 .LUT_INIT=16'b0010000010100000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_RNI6CD2C_28_LC_12_24_1  (
            .in0(N__60116),
            .in1(N__55492),
            .in2(N__52164),
            .in3(N__52161),
            .lcout(\pid_front.error_i_acumm_2_sqmuxa ),
            .ltout(\pid_front.error_i_acumm_2_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_10_LC_12_24_2 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_10_LC_12_24_2 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_10_LC_12_24_2 .LUT_INIT=16'b1111100000001000;
    LogicCell40 \pid_front.error_i_acumm_10_LC_12_24_2  (
            .in0(N__52414),
            .in1(N__60119),
            .in2(N__52155),
            .in3(N__52148),
            .lcout(\pid_front.error_i_acummZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87198),
            .ce(N__60005),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_4_LC_12_24_3 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_4_LC_12_24_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_4_LC_12_24_3 .LUT_INIT=16'b1111000010001000;
    LogicCell40 \pid_front.error_i_acumm_4_LC_12_24_3  (
            .in0(N__60117),
            .in1(N__52416),
            .in2(N__52119),
            .in3(N__52388),
            .lcout(\pid_front.error_i_acummZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87198),
            .ce(N__60005),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_5_LC_12_24_4 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_5_LC_12_24_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_5_LC_12_24_4 .LUT_INIT=16'b1110101001000000;
    LogicCell40 \pid_front.error_i_acumm_5_LC_12_24_4  (
            .in0(N__52389),
            .in1(N__60121),
            .in2(N__52425),
            .in3(N__52095),
            .lcout(\pid_front.error_i_acummZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87198),
            .ce(N__60005),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_6_LC_12_24_5 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_6_LC_12_24_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_6_LC_12_24_5 .LUT_INIT=16'b1111000010001000;
    LogicCell40 \pid_front.error_i_acumm_6_LC_12_24_5  (
            .in0(N__60118),
            .in1(N__52417),
            .in2(N__52479),
            .in3(N__52390),
            .lcout(\pid_front.error_i_acummZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87198),
            .ce(N__60005),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_13_LC_12_24_6 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_13_LC_12_24_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_13_LC_12_24_6 .LUT_INIT=16'b1110101001000000;
    LogicCell40 \pid_front.error_i_acumm_13_LC_12_24_6  (
            .in0(N__52387),
            .in1(N__60120),
            .in2(N__52424),
            .in3(N__52674),
            .lcout(\pid_front.error_i_acummZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87198),
            .ce(N__60005),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_11_LC_12_24_7 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_11_LC_12_24_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_11_LC_12_24_7 .LUT_INIT=16'b1010101011000000;
    LogicCell40 \pid_front.error_i_acumm_11_LC_12_24_7  (
            .in0(N__52451),
            .in1(N__52415),
            .in2(N__60128),
            .in3(N__52386),
            .lcout(\pid_front.error_i_acummZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87198),
            .ce(N__60005),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI2BC9_0_1_LC_12_25_0 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI2BC9_0_1_LC_12_25_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI2BC9_0_1_LC_12_25_0 .LUT_INIT=16'b1111001101110001;
    LogicCell40 \pid_front.error_p_reg_esr_RNI2BC9_0_1_LC_12_25_0  (
            .in0(N__52231),
            .in1(N__52586),
            .in2(N__52281),
            .in3(N__52251),
            .lcout(),
            .ltout(\pid_front.error_p_reg_esr_RNI2BC9_0Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNIFSHO_1_LC_12_25_1 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIFSHO_1_LC_12_25_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIFSHO_1_LC_12_25_1 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIFSHO_1_LC_12_25_1  (
            .in0(N__52558),
            .in1(_gnd_net_),
            .in2(N__52353),
            .in3(N__52260),
            .lcout(\pid_front.error_d_reg_prev_esr_RNIFSHOZ0Z_1 ),
            .ltout(\pid_front.error_d_reg_prev_esr_RNIFSHOZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNID19M1_1_LC_12_25_2 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNID19M1_1_LC_12_25_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNID19M1_1_LC_12_25_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNID19M1_1_LC_12_25_2  (
            .in0(N__54757),
            .in1(N__52331),
            .in2(N__52350),
            .in3(N__52596),
            .lcout(\pid_front.error_d_reg_prev_esr_RNID19M1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_RNI1JN71_1_LC_12_25_3 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNI1JN71_1_LC_12_25_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNI1JN71_1_LC_12_25_3 .LUT_INIT=16'b1110111110001100;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNI1JN71_1_LC_12_25_3  (
            .in0(N__52588),
            .in1(N__52332),
            .in2(N__52565),
            .in3(N__52314),
            .lcout(\pid_front.error_d_reg_prev_esr_RNI1JN71Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNI2BC9_1_LC_12_25_4 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNI2BC9_1_LC_12_25_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNI2BC9_1_LC_12_25_4 .LUT_INIT=16'b1111110011010100;
    LogicCell40 \pid_front.error_p_reg_esr_RNI2BC9_1_LC_12_25_4  (
            .in0(N__52230),
            .in1(N__52585),
            .in2(N__52280),
            .in3(N__52250),
            .lcout(\pid_front.error_p_reg_esr_RNI2BC9Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_0_LC_12_25_5 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_0_LC_12_25_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_0_LC_12_25_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_front.error_d_reg_prev_esr_0_LC_12_25_5  (
            .in0(N__52252),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_d_reg_prevZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87217),
            .ce(N__70453),
            .sr(N__70346));
    defparam \pid_front.error_d_reg_prev_esr_RNIQHN6_1_LC_12_25_6 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_RNIQHN6_1_LC_12_25_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_d_reg_prev_esr_RNIQHN6_1_LC_12_25_6 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \pid_front.error_d_reg_prev_esr_RNIQHN6_1_LC_12_25_6  (
            .in0(_gnd_net_),
            .in1(N__52557),
            .in2(_gnd_net_),
            .in3(N__52587),
            .lcout(\pid_front.error_d_reg_prev_esr_RNIQHN6Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_1_LC_12_25_7 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_1_LC_12_25_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_1_LC_12_25_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_front.error_d_reg_prev_esr_1_LC_12_25_7  (
            .in0(N__52589),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_d_reg_prevZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87217),
            .ce(N__70453),
            .sr(N__70346));
    defparam \pid_front.error_i_acumm_prereg_esr_21_LC_12_26_0 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_21_LC_12_26_0 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_21_LC_12_26_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_21_LC_12_26_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55712),
            .lcout(\pid_front.error_i_acumm_preregZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87230),
            .ce(N__56079),
            .sr(N__79694));
    defparam \pid_front.error_i_acumm_prereg_esr_13_LC_12_26_1 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_13_LC_12_26_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_13_LC_12_26_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_13_LC_12_26_1  (
            .in0(N__55458),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_i_acumm_preregZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87230),
            .ce(N__56079),
            .sr(N__79694));
    defparam \pid_front.error_i_acumm_prereg_esr_22_LC_12_26_2 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_22_LC_12_26_2 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_22_LC_12_26_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_22_LC_12_26_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55685),
            .lcout(\pid_front.error_i_acumm_preregZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87230),
            .ce(N__56079),
            .sr(N__79694));
    defparam \pid_front.error_i_acumm_prereg_esr_8_LC_12_26_3 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_8_LC_12_26_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_8_LC_12_26_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_8_LC_12_26_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55076),
            .lcout(\pid_front.error_i_acumm_preregZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87230),
            .ce(N__56079),
            .sr(N__79694));
    defparam \pid_front.error_i_acumm_prereg_esr_24_LC_12_26_4 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_24_LC_12_26_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_24_LC_12_26_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_24_LC_12_26_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55655),
            .lcout(\pid_front.error_i_acumm_preregZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87230),
            .ce(N__56079),
            .sr(N__79694));
    defparam \pid_front.error_i_acumm_prereg_esr_16_LC_12_26_5 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_16_LC_12_26_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_16_LC_12_26_5 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_16_LC_12_26_5  (
            .in0(_gnd_net_),
            .in1(N__55345),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_i_acumm_preregZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87230),
            .ce(N__56079),
            .sr(N__79694));
    defparam \pid_front.error_i_acumm_prereg_esr_20_LC_12_26_6 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_20_LC_12_26_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_20_LC_12_26_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_20_LC_12_26_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55241),
            .lcout(\pid_front.error_i_acumm_preregZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87230),
            .ce(N__56079),
            .sr(N__79694));
    defparam \pid_front.error_i_acumm_prereg_esr_12_LC_12_26_7 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_12_LC_12_26_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_12_LC_12_26_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_12_LC_12_26_7  (
            .in0(N__54931),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.un10lto12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87230),
            .ce(N__56079),
            .sr(N__79694));
    defparam \pid_front.error_i_acumm_prereg_esr_RNI6IK41_0_22_LC_12_27_0 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_RNI6IK41_0_22_LC_12_27_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_acumm_prereg_esr_RNI6IK41_0_22_LC_12_27_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_RNI6IK41_0_22_LC_12_27_0  (
            .in0(N__56220),
            .in1(N__56264),
            .in2(N__52686),
            .in3(N__52695),
            .lcout(\pid_front.error_i_acumm16lto27_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_prereg_esr_RNI9HER_26_LC_12_27_1 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_RNI9HER_26_LC_12_27_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_acumm_prereg_esr_RNI9HER_26_LC_12_27_1 .LUT_INIT=16'b0000000000000101;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_RNI9HER_26_LC_12_27_1  (
            .in0(N__52670),
            .in1(_gnd_net_),
            .in2(N__52647),
            .in3(N__56184),
            .lcout(),
            .ltout(\pid_front.error_i_acumm16lto27_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_prereg_esr_RNI18694_14_LC_12_27_2 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_RNI18694_14_LC_12_27_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_acumm_prereg_esr_RNI18694_14_LC_12_27_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_RNI18694_14_LC_12_27_2  (
            .in0(N__52728),
            .in1(N__52722),
            .in2(N__52713),
            .in3(N__52710),
            .lcout(\pid_front.error_i_acumm16lto27_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_prereg_esr_RNI6IK41_22_LC_12_27_5 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_RNI6IK41_22_LC_12_27_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_acumm_prereg_esr_RNI6IK41_22_LC_12_27_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_RNI6IK41_22_LC_12_27_5  (
            .in0(N__52694),
            .in1(N__52682),
            .in2(N__56265),
            .in3(N__56219),
            .lcout(),
            .ltout(\pid_front.un10lto27_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_prereg_esr_RNIF3302_26_LC_12_27_6 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_RNIF3302_26_LC_12_27_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_acumm_prereg_esr_RNIF3302_26_LC_12_27_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_RNIF3302_26_LC_12_27_6  (
            .in0(N__56183),
            .in1(N__52669),
            .in2(N__52656),
            .in3(N__52643),
            .lcout(\pid_front.un10lto27_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_prereg_esr_26_LC_12_27_7 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_26_LC_12_27_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_26_LC_12_27_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_26_LC_12_27_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55625),
            .lcout(\pid_front.error_i_acumm_preregZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87244),
            .ce(N__56077),
            .sr(N__79700));
    defparam \ppm_encoder_1.elevator_RNIPFGE_11_LC_13_1_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNIPFGE_11_LC_13_1_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNIPFGE_11_LC_13_1_0 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \ppm_encoder_1.elevator_RNIPFGE_11_LC_13_1_0  (
            .in0(N__52635),
            .in1(N__52828),
            .in2(_gnd_net_),
            .in3(N__52945),
            .lcout(),
            .ltout(\ppm_encoder_1.elevator_RNIPFGEZ0Z_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.rudder_RNIKAJ92_11_LC_13_1_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_RNIKAJ92_11_LC_13_1_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.rudder_RNIKAJ92_11_LC_13_1_1 .LUT_INIT=16'b1111111111110100;
    LogicCell40 \ppm_encoder_1.rudder_RNIKAJ92_11_LC_13_1_1  (
            .in0(N__53618),
            .in1(N__60907),
            .in2(N__52599),
            .in3(N__57066),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_2_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIPA8G4_11_LC_13_1_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIPA8G4_11_LC_13_1_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIPA8G4_11_LC_13_1_2 .LUT_INIT=16'b1010100101010110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIPA8G4_11_LC_13_1_2  (
            .in0(N__53062),
            .in1(N__57345),
            .in2(N__53082),
            .in3(N__56944),
            .lcout(),
            .ltout(\ppm_encoder_1.un1_init_pulses_0_axb_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNI4JPF5_11_LC_13_1_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI4JPF5_11_LC_13_1_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI4JPF5_11_LC_13_1_3 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI4JPF5_11_LC_13_1_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__53079),
            .in3(N__53015),
            .lcout(\ppm_encoder_1.init_pulses_RNI4JPF5Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIB8HV_11_LC_13_1_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIB8HV_11_LC_13_1_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIB8HV_11_LC_13_1_4 .LUT_INIT=16'b1111000001111000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIB8HV_11_LC_13_1_4  (
            .in0(N__60905),
            .in1(N__61019),
            .in2(N__53064),
            .in3(N__64269),
            .lcout(\ppm_encoder_1.N_266_i_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_2_LC_13_1_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_2_LC_13_1_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_2_LC_13_1_5 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_2_LC_13_1_5  (
            .in0(_gnd_net_),
            .in1(N__68625),
            .in2(_gnd_net_),
            .in3(N__53343),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNITJK21_4_LC_13_1_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNITJK21_4_LC_13_1_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNITJK21_4_LC_13_1_7 .LUT_INIT=16'b1001110011001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNITJK21_4_LC_13_1_7  (
            .in0(N__64268),
            .in1(N__59716),
            .in2(N__61043),
            .in3(N__60906),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_13_LC_13_2_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_13_LC_13_2_0 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_13_LC_13_2_0 .LUT_INIT=16'b0010001100100000;
    LogicCell40 \ppm_encoder_1.init_pulses_13_LC_13_2_0  (
            .in0(N__52995),
            .in1(N__55822),
            .in2(N__55908),
            .in3(N__52986),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__86969),
            .ce(),
            .sr(N__79563));
    defparam \ppm_encoder_1.init_pulses_2_LC_13_2_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_2_LC_13_2_2 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_2_LC_13_2_2 .LUT_INIT=16'b0000000011011000;
    LogicCell40 \ppm_encoder_1.init_pulses_2_LC_13_2_2  (
            .in0(N__55876),
            .in1(N__52974),
            .in2(N__52962),
            .in3(N__55823),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__86969),
            .ce(),
            .sr(N__79563));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNIUTMR_LC_13_2_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNIUTMR_LC_13_2_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNIUTMR_LC_13_2_3 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNIUTMR_LC_13_2_3  (
            .in0(N__63803),
            .in1(N__52829),
            .in2(_gnd_net_),
            .in3(N__52946),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNIUTMRZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_3_LC_13_2_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_3_LC_13_2_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_3_LC_13_2_6 .LUT_INIT=16'b1000010110000000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_3_LC_13_2_6  (
            .in0(N__52947),
            .in1(N__52866),
            .in2(N__52833),
            .in3(N__63804),
            .lcout(),
            .ltout(\ppm_encoder_1.pulses2count_9_0_0_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_3_LC_13_2_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_3_LC_13_2_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_3_LC_13_2_7 .LUT_INIT=16'b1111110011110000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_3_LC_13_2_7  (
            .in0(_gnd_net_),
            .in1(N__64398),
            .in2(N__53235),
            .in3(N__53226),
            .lcout(\ppm_encoder_1.pulses2count_9_0_0_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNI9B0E1_0_LC_13_3_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNI9B0E1_0_LC_13_3_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNI9B0E1_0_LC_13_3_0 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \ppm_encoder_1.throttle_RNI9B0E1_0_LC_13_3_0  (
            .in0(N__53137),
            .in1(N__58010),
            .in2(N__53126),
            .in3(N__57166),
            .lcout(\ppm_encoder_1.un2_throttle_iv_0_0_0 ),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNI25564_0_LC_13_3_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNI25564_0_LC_13_3_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNI25564_0_LC_13_3_1 .LUT_INIT=16'b1111111111111010;
    LogicCell40 \ppm_encoder_1.throttle_RNI25564_0_LC_13_3_1  (
            .in0(N__53181),
            .in1(N__53964),
            .in2(N__53193),
            .in3(N__57057),
            .lcout(\ppm_encoder_1.throttle_RNI25564Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNIV0IU_0_LC_13_3_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNIV0IU_0_LC_13_3_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNIV0IU_0_LC_13_3_2 .LUT_INIT=16'b1110101010101010;
    LogicCell40 \ppm_encoder_1.elevator_RNIV0IU_0_LC_13_3_2  (
            .in0(N__57261),
            .in1(N__57606),
            .in2(N__63617),
            .in3(N__57212),
            .lcout(\ppm_encoder_1.un2_throttle_iv_0_1_0 ),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_0_LC_13_3_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNO_0_0_LC_13_3_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_0_LC_13_3_3 .LUT_INIT=16'b0011001100110110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_0_LC_13_3_3  (
            .in0(N__53175),
            .in1(N__53963),
            .in2(N__53169),
            .in3(N__57058),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_0_LC_13_3_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_0_LC_13_3_4 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.aileron_0_LC_13_3_4 .LUT_INIT=16'b0010001011101110;
    LogicCell40 \ppm_encoder_1.aileron_0_LC_13_3_4  (
            .in0(N__53139),
            .in1(N__65243),
            .in2(_gnd_net_),
            .in3(N__53811),
            .lcout(\ppm_encoder_1.aileronZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__86971),
            .ce(),
            .sr(N__79568));
    defparam \ppm_encoder_1.throttle_0_LC_13_3_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_0_LC_13_3_5 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.throttle_0_LC_13_3_5 .LUT_INIT=16'b0111011100100010;
    LogicCell40 \ppm_encoder_1.throttle_0_LC_13_3_5  (
            .in0(N__65247),
            .in1(N__53166),
            .in2(_gnd_net_),
            .in3(N__53125),
            .lcout(\ppm_encoder_1.throttleZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__86971),
            .ce(),
            .sr(N__79568));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_0_LC_13_3_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_0_LC_13_3_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_0_LC_13_3_6 .LUT_INIT=16'b0011000010001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_0_LC_13_3_6  (
            .in0(N__53138),
            .in1(N__61417),
            .in2(N__53127),
            .in3(N__61631),
            .lcout(\ppm_encoder_1.pulses2count_9_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_0_LC_13_3_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_0_LC_13_3_7 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.elevator_0_LC_13_3_7 .LUT_INIT=16'b0101111101010000;
    LogicCell40 \ppm_encoder_1.elevator_0_LC_13_3_7  (
            .in0(N__53109),
            .in1(_gnd_net_),
            .in2(N__65295),
            .in3(N__63613),
            .lcout(\ppm_encoder_1.elevatorZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__86971),
            .ce(),
            .sr(N__79568));
    defparam \ppm_encoder_1.aileron_esr_RNI5B2L1_14_LC_13_4_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_esr_RNI5B2L1_14_LC_13_4_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.aileron_esr_RNI5B2L1_14_LC_13_4_0 .LUT_INIT=16'b0101110100001100;
    LogicCell40 \ppm_encoder_1.aileron_esr_RNI5B2L1_14_LC_13_4_0  (
            .in0(N__57536),
            .in1(N__57990),
            .in2(N__57573),
            .in3(N__57155),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_i_i_0_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIVCA75_14_LC_13_4_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIVCA75_14_LC_13_4_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIVCA75_14_LC_13_4_1 .LUT_INIT=16'b0011001100110110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIVCA75_14_LC_13_4_1  (
            .in0(N__57470),
            .in1(N__53274),
            .in2(N__53310),
            .in3(N__57056),
            .lcout(),
            .ltout(\ppm_encoder_1.un1_init_pulses_0_axb_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIE8336_14_LC_13_4_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIE8336_14_LC_13_4_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIE8336_14_LC_13_4_2 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIE8336_14_LC_13_4_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__53307),
            .in3(N__53285),
            .lcout(\ppm_encoder_1.init_pulses_RNIE8336Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.PPM_STATE_RNIV4V5_1_LC_13_4_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_RNIV4V5_1_LC_13_4_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.PPM_STATE_RNIV4V5_1_LC_13_4_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \ppm_encoder_1.PPM_STATE_RNIV4V5_1_LC_13_4_3  (
            .in0(_gnd_net_),
            .in1(N__61202),
            .in2(_gnd_net_),
            .in3(N__61135),
            .lcout(\ppm_encoder_1.PPM_STATE_RNIV4V5Z0Z_1 ),
            .ltout(\ppm_encoder_1.PPM_STATE_RNIV4V5Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIFROR_14_LC_13_4_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIFROR_14_LC_13_4_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIFROR_14_LC_13_4_4 .LUT_INIT=16'b1100011011001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIFROR_14_LC_13_4_4  (
            .in0(N__61053),
            .in1(N__57505),
            .in2(N__53295),
            .in3(N__63391),
            .lcout(\ppm_encoder_1.N_269_i_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIFROR_0_14_LC_13_4_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIFROR_0_14_LC_13_4_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIFROR_0_14_LC_13_4_5 .LUT_INIT=16'b0000111110000111;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIFROR_0_14_LC_13_4_5  (
            .in0(N__63390),
            .in1(N__61052),
            .in2(N__57509),
            .in3(N__64239),
            .lcout(\ppm_encoder_1.N_269_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.PPM_STATE_1_LC_13_4_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_1_LC_13_4_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.PPM_STATE_1_LC_13_4_6 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \ppm_encoder_1.PPM_STATE_1_LC_13_4_6  (
            .in0(N__61136),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61178),
            .lcout(\ppm_encoder_1.PPM_STATEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__86973),
            .ce(),
            .sr(N__79571));
    defparam \ppm_encoder_1.PPM_STATE_0_LC_13_4_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_0_LC_13_4_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.PPM_STATE_0_LC_13_4_7 .LUT_INIT=16'b1010101010111011;
    LogicCell40 \ppm_encoder_1.PPM_STATE_0_LC_13_4_7  (
            .in0(N__61179),
            .in1(N__53268),
            .in2(_gnd_net_),
            .in3(N__61203),
            .lcout(\ppm_encoder_1.PPM_STATEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__86973),
            .ce(),
            .sr(N__79571));
    defparam \ppm_encoder_1.aileron_RNIFUAP_1_LC_13_5_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_RNIFUAP_1_LC_13_5_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.aileron_RNIFUAP_1_LC_13_5_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \ppm_encoder_1.aileron_RNIFUAP_1_LC_13_5_0  (
            .in0(_gnd_net_),
            .in1(N__53251),
            .in2(_gnd_net_),
            .in3(N__57122),
            .lcout(\ppm_encoder_1.aileron_RNIFUAPZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m9_0_i_o2_LC_13_5_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m9_0_i_o2_LC_13_5_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m9_0_i_o2_LC_13_5_1 .LUT_INIT=16'b0000111111111111;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m9_0_i_o2_LC_13_5_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__57602),
            .in3(N__57209),
            .lcout(\ppm_encoder_1.m9_0_i_o2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIHO7D_0_LC_13_5_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIHO7D_0_LC_13_5_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIHO7D_0_LC_13_5_2 .LUT_INIT=16'b1110111011101110;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIHO7D_0_LC_13_5_2  (
            .in0(N__57210),
            .in1(N__57597),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIHO7DZ0Z_0 ),
            .ltout(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIHO7DZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI5QE01_3_LC_13_5_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI5QE01_3_LC_13_5_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI5QE01_3_LC_13_5_3 .LUT_INIT=16'b1111111111101101;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI5QE01_3_LC_13_5_3  (
            .in0(N__57256),
            .in1(N__53579),
            .in2(N__53352),
            .in3(N__64101),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI5QE01Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un11lto30_i_a2_2_c_RNO_LC_13_5_4 .C_ON=1'b0;
    defparam \pid_side.un11lto30_i_a2_2_c_RNO_LC_13_5_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.un11lto30_i_a2_2_c_RNO_LC_13_5_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_side.un11lto30_i_a2_2_c_RNO_LC_13_5_4  (
            .in0(N__71670),
            .in1(N__71838),
            .in2(N__71772),
            .in3(N__71631),
            .lcout(\pid_side.N_11_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIBSME1_10_LC_13_5_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIBSME1_10_LC_13_5_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIBSME1_10_LC_13_5_5 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \ppm_encoder_1.throttle_RNIBSME1_10_LC_13_5_5  (
            .in0(N__57124),
            .in1(N__60759),
            .in2(N__56816),
            .in3(N__57982),
            .lcout(\ppm_encoder_1.un2_throttle_iv_0_1_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIJQ7D_1_LC_13_5_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIJQ7D_1_LC_13_5_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIJQ7D_1_LC_13_5_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIJQ7D_1_LC_13_5_6  (
            .in0(_gnd_net_),
            .in1(N__57255),
            .in2(_gnd_net_),
            .in3(N__57593),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIJQ7DZ0Z_1 ),
            .ltout(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIJQ7DZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIDF0E1_2_LC_13_5_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIDF0E1_2_LC_13_5_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIDF0E1_2_LC_13_5_7 .LUT_INIT=16'b0011000010111010;
    LogicCell40 \ppm_encoder_1.throttle_RNIDF0E1_2_LC_13_5_7  (
            .in0(N__57123),
            .in1(N__53339),
            .in2(N__53313),
            .in3(N__68843),
            .lcout(\ppm_encoder_1.un2_throttle_iv_0_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep2_LC_13_6_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep2_LC_13_6_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep2_LC_13_6_1 .LUT_INIT=16'b0100010000000101;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_2_rep2_LC_13_6_1  (
            .in0(N__79981),
            .in1(N__60897),
            .in2(N__57417),
            .in3(N__64302),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__86983),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNINP0E1_7_LC_13_6_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNINP0E1_7_LC_13_6_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNINP0E1_7_LC_13_6_2 .LUT_INIT=16'b0101110100001100;
    LogicCell40 \ppm_encoder_1.throttle_RNINP0E1_7_LC_13_6_2  (
            .in0(N__53678),
            .in1(N__57978),
            .in2(N__53652),
            .in3(N__57144),
            .lcout(\ppm_encoder_1.un2_throttle_iv_0_0_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.rudder_RNIUTSI2_7_LC_13_6_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_RNIUTSI2_7_LC_13_6_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.rudder_RNIUTSI2_7_LC_13_6_3 .LUT_INIT=16'b1111111111001110;
    LogicCell40 \ppm_encoder_1.rudder_RNIUTSI2_7_LC_13_6_3  (
            .in0(N__60859),
            .in1(N__57824),
            .in2(N__57869),
            .in3(N__57025),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_0_1_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNI28VR4_7_LC_13_6_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI28VR4_7_LC_13_6_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI28VR4_7_LC_13_6_4 .LUT_INIT=16'b1001100110010110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI28VR4_7_LC_13_6_4  (
            .in0(N__56719),
            .in1(N__56924),
            .in2(N__53496),
            .in3(N__53493),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNI0NK21_7_LC_13_6_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI0NK21_7_LC_13_6_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI0NK21_7_LC_13_6_5 .LUT_INIT=16'b1111011100001000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI0NK21_7_LC_13_6_5  (
            .in0(N__60860),
            .in1(N__60986),
            .in2(N__64304),
            .in3(N__56720),
            .lcout(\ppm_encoder_1.N_263_i_i ),
            .ltout(\ppm_encoder_1.N_263_i_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNI2VJU5_7_LC_13_6_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI2VJU5_7_LC_13_6_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI2VJU5_7_LC_13_6_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI2VJU5_7_LC_13_6_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__53472),
            .in3(N__53469),
            .lcout(\ppm_encoder_1.init_pulses_RNI2VJU5Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_3_rep2_LC_13_6_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_3_rep2_LC_13_6_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_3_rep2_LC_13_6_7 .LUT_INIT=16'b0100010000000101;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_3_rep2_LC_13_6_7  (
            .in0(N__79982),
            .in1(N__60987),
            .in2(N__63903),
            .in3(N__64303),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_3_repZ0Z2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__86983),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNI2L8G4_13_LC_13_7_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI2L8G4_13_LC_13_7_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI2L8G4_13_LC_13_7_0 .LUT_INIT=16'b0101101001101001;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI2L8G4_13_LC_13_7_0  (
            .in0(N__56945),
            .in1(N__53397),
            .in2(N__53382),
            .in3(N__53403),
            .lcout(),
            .ltout(\ppm_encoder_1.un1_init_pulses_0_axb_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIFVPF5_13_LC_13_7_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIFVPF5_13_LC_13_7_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIFVPF5_13_LC_13_7_1 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIFVPF5_13_LC_13_7_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__53451),
            .in3(N__53444),
            .lcout(\ppm_encoder_1.init_pulses_RNIFVPF5Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNINEJ92_13_LC_13_7_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNINEJ92_13_LC_13_7_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNINEJ92_13_LC_13_7_2 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \ppm_encoder_1.elevator_RNINEJ92_13_LC_13_7_2  (
            .in0(N__53543),
            .in1(N__53390),
            .in2(_gnd_net_),
            .in3(N__57051),
            .lcout(\ppm_encoder_1.un2_throttle_iv_0_1_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIH2NE1_13_LC_13_7_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIH2NE1_13_LC_13_7_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIH2NE1_13_LC_13_7_3 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \ppm_encoder_1.throttle_RNIH2NE1_13_LC_13_7_3  (
            .in0(N__61303),
            .in1(N__58009),
            .in2(N__61487),
            .in3(N__57183),
            .lcout(\ppm_encoder_1.un2_throttle_iv_0_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_13_LC_13_7_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_13_LC_13_7_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_13_LC_13_7_5 .LUT_INIT=16'b1111111111101010;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_13_LC_13_7_5  (
            .in0(N__53391),
            .in1(N__53381),
            .in2(N__64449),
            .in3(N__53544),
            .lcout(\ppm_encoder_1.pulses2count_9_0_2_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.rudder_13_LC_13_7_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_13_LC_13_7_7 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.rudder_13_LC_13_7_7 .LUT_INIT=16'b1001100111110000;
    LogicCell40 \ppm_encoder_1.rudder_13_LC_13_7_7  (
            .in0(N__53712),
            .in1(N__53691),
            .in2(N__53559),
            .in3(N__65081),
            .lcout(\ppm_encoder_1.rudderZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__86991),
            .ce(),
            .sr(N__79591));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_7_LC_13_8_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_7_LC_13_8_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_7_LC_13_8_0 .LUT_INIT=16'b0001000100001010;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_7_LC_13_8_0  (
            .in0(N__61604),
            .in1(N__53671),
            .in2(N__53651),
            .in3(N__61458),
            .lcout(\ppm_encoder_1.pulses2count_9_i_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_11_LC_13_8_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_11_LC_13_8_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_11_LC_13_8_3 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_11_LC_13_8_3  (
            .in0(N__53622),
            .in1(N__60923),
            .in2(_gnd_net_),
            .in3(N__63857),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.source_data_valid_esr_RNO_LC_13_8_4 .C_ON=1'b0;
    defparam \pid_alt.source_data_valid_esr_RNO_LC_13_8_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.source_data_valid_esr_RNO_LC_13_8_4 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \pid_alt.source_data_valid_esr_RNO_LC_13_8_4  (
            .in0(_gnd_net_),
            .in1(N__56030),
            .in2(_gnd_net_),
            .in3(N__79963),
            .lcout(\pid_alt.state_1_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_3_LC_13_8_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_3_LC_13_8_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_3_LC_13_8_6 .LUT_INIT=16'b0000000011000101;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_3_LC_13_8_6  (
            .in0(N__63907),
            .in1(N__53578),
            .in2(N__64305),
            .in3(N__79964),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__86999),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.rudder_RNIN2KQ_13_LC_13_8_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_RNIN2KQ_13_LC_13_8_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.rudder_RNIN2KQ_13_LC_13_8_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ppm_encoder_1.rudder_RNIN2KQ_13_LC_13_8_7  (
            .in0(_gnd_net_),
            .in1(N__63741),
            .in2(_gnd_net_),
            .in3(N__53555),
            .lcout(\ppm_encoder_1.rudder_RNIN2KQZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.source_pid_1_esr_5_LC_13_9_0 .C_ON=1'b0;
    defparam \pid_side.source_pid_1_esr_5_LC_13_9_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.source_pid_1_esr_5_LC_13_9_0 .LUT_INIT=16'b1101110000000000;
    LogicCell40 \pid_side.source_pid_1_esr_5_LC_13_9_0  (
            .in0(N__71595),
            .in1(N__69999),
            .in2(N__58120),
            .in3(N__69375),
            .lcout(side_order_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87004),
            .ce(N__58281),
            .sr(N__58251));
    defparam \pid_side.source_pid_1_esr_7_LC_13_9_1 .C_ON=1'b0;
    defparam \pid_side.source_pid_1_esr_7_LC_13_9_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.source_pid_1_esr_7_LC_13_9_1 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \pid_side.source_pid_1_esr_7_LC_13_9_1  (
            .in0(N__69993),
            .in1(N__58107),
            .in2(_gnd_net_),
            .in3(N__71805),
            .lcout(side_order_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87004),
            .ce(N__58281),
            .sr(N__58251));
    defparam \pid_side.source_pid_1_esr_3_LC_13_9_2 .C_ON=1'b0;
    defparam \pid_side.source_pid_1_esr_3_LC_13_9_2 .SEQ_MODE=4'b1000;
    defparam \pid_side.source_pid_1_esr_3_LC_13_9_2 .LUT_INIT=16'b0000000011100000;
    LogicCell40 \pid_side.source_pid_1_esr_3_LC_13_9_2  (
            .in0(N__58110),
            .in1(N__69998),
            .in2(N__69090),
            .in3(N__58152),
            .lcout(side_order_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87004),
            .ce(N__58281),
            .sr(N__58251));
    defparam \pid_side.source_pid_1_esr_11_LC_13_9_3 .C_ON=1'b0;
    defparam \pid_side.source_pid_1_esr_11_LC_13_9_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.source_pid_1_esr_11_LC_13_9_3 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \pid_side.source_pid_1_esr_11_LC_13_9_3  (
            .in0(N__69992),
            .in1(N__58103),
            .in2(_gnd_net_),
            .in3(N__71771),
            .lcout(side_order_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87004),
            .ce(N__58281),
            .sr(N__58251));
    defparam \pid_side.source_pid_1_esr_1_LC_13_9_4 .C_ON=1'b0;
    defparam \pid_side.source_pid_1_esr_1_LC_13_9_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.source_pid_1_esr_1_LC_13_9_4 .LUT_INIT=16'b0000000011100000;
    LogicCell40 \pid_side.source_pid_1_esr_1_LC_13_9_4  (
            .in0(N__58109),
            .in1(N__69997),
            .in2(N__69153),
            .in3(N__58151),
            .lcout(side_order_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87004),
            .ce(N__58281),
            .sr(N__58251));
    defparam \pid_side.source_pid_1_esr_0_LC_13_9_5 .C_ON=1'b0;
    defparam \pid_side.source_pid_1_esr_0_LC_13_9_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.source_pid_1_esr_0_LC_13_9_5 .LUT_INIT=16'b0000111000000000;
    LogicCell40 \pid_side.source_pid_1_esr_0_LC_13_9_5  (
            .in0(N__69994),
            .in1(N__58108),
            .in2(N__58157),
            .in3(N__69195),
            .lcout(side_order_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87004),
            .ce(N__58281),
            .sr(N__58251));
    defparam \pid_side.source_pid_1_esr_10_LC_13_9_6 .C_ON=1'b0;
    defparam \pid_side.source_pid_1_esr_10_LC_13_9_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.source_pid_1_esr_10_LC_13_9_6 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \pid_side.source_pid_1_esr_10_LC_13_9_6  (
            .in0(N__58102),
            .in1(N__69996),
            .in2(_gnd_net_),
            .in3(N__71837),
            .lcout(side_order_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87004),
            .ce(N__58281),
            .sr(N__58251));
    defparam \pid_side.source_pid_1_esr_4_LC_13_9_7 .C_ON=1'b0;
    defparam \pid_side.source_pid_1_esr_4_LC_13_9_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.source_pid_1_esr_4_LC_13_9_7 .LUT_INIT=16'b1111111111110001;
    LogicCell40 \pid_side.source_pid_1_esr_4_LC_13_9_7  (
            .in0(N__69995),
            .in1(N__58111),
            .in2(N__58158),
            .in3(N__69416),
            .lcout(side_order_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87004),
            .ce(N__58281),
            .sr(N__58251));
    defparam \pid_side.pid_prereg_esr_RNII463_20_LC_13_10_0 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_esr_RNII463_20_LC_13_10_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_esr_RNII463_20_LC_13_10_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_side.pid_prereg_esr_RNII463_20_LC_13_10_0  (
            .in0(N__69747),
            .in1(N__69762),
            .in2(N__69717),
            .in3(N__69432),
            .lcout(\pid_side.un11lto30_i_a2_4_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.source_pid_1_esr_8_LC_13_10_6 .C_ON=1'b0;
    defparam \pid_side.source_pid_1_esr_8_LC_13_10_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.source_pid_1_esr_8_LC_13_10_6 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \pid_side.source_pid_1_esr_8_LC_13_10_6  (
            .in0(N__58118),
            .in1(N__70006),
            .in2(_gnd_net_),
            .in3(N__71630),
            .lcout(side_order_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87012),
            .ce(N__58292),
            .sr(N__58246));
    defparam \pid_side.source_pid_1_esr_9_LC_13_10_7 .C_ON=1'b0;
    defparam \pid_side.source_pid_1_esr_9_LC_13_10_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.source_pid_1_esr_9_LC_13_10_7 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \pid_side.source_pid_1_esr_9_LC_13_10_7  (
            .in0(N__70005),
            .in1(N__58119),
            .in2(_gnd_net_),
            .in3(N__71669),
            .lcout(side_order_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87012),
            .ce(N__58292),
            .sr(N__58246));
    defparam \pid_side.state_RNI7OA81_0_LC_13_11_0 .C_ON=1'b0;
    defparam \pid_side.state_RNI7OA81_0_LC_13_11_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.state_RNI7OA81_0_LC_13_11_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \pid_side.state_RNI7OA81_0_LC_13_11_0  (
            .in0(_gnd_net_),
            .in1(N__69909),
            .in2(_gnd_net_),
            .in3(N__83177),
            .lcout(\pid_side.N_838_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_2_LC_13_11_1 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_2_LC_13_11_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_2_LC_13_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_2_LC_13_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82449),
            .lcout(\pid_side.error_d_reg_prevZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87019),
            .ce(N__83329),
            .sr(N__83218));
    defparam \pid_side.error_d_reg_prev_esr_4_LC_13_11_2 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_4_LC_13_11_2 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_4_LC_13_11_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_4_LC_13_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81531),
            .lcout(\pid_side.error_d_reg_prevZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87019),
            .ce(N__83329),
            .sr(N__83218));
    defparam \pid_side.error_d_reg_prev_esr_7_LC_13_11_3 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_7_LC_13_11_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_7_LC_13_11_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_7_LC_13_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81234),
            .lcout(\pid_side.error_d_reg_prevZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87019),
            .ce(N__83329),
            .sr(N__83218));
    defparam \pid_side.error_d_reg_prev_esr_5_LC_13_11_4 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_5_LC_13_11_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_5_LC_13_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_5_LC_13_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81381),
            .lcout(\pid_side.error_d_reg_prevZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87019),
            .ce(N__83329),
            .sr(N__83218));
    defparam \ppm_encoder_1.counter_RNI5K08_0_LC_13_11_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter_RNI5K08_0_LC_13_11_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter_RNI5K08_0_LC_13_11_5 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \ppm_encoder_1.counter_RNI5K08_0_LC_13_11_5  (
            .in0(_gnd_net_),
            .in1(N__63999),
            .in2(_gnd_net_),
            .in3(N__64026),
            .lcout(\ppm_encoder_1.N_486_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_0_LC_13_11_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNO_1_0_LC_13_11_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_0_LC_13_11_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_0_LC_13_11_6  (
            .in0(_gnd_net_),
            .in1(N__53982),
            .in2(_gnd_net_),
            .in3(N__57333),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.N_2725_i_l_ofx_LC_13_11_7 .C_ON=1'b0;
    defparam \scaler_4.N_2725_i_l_ofx_LC_13_11_7 .SEQ_MODE=4'b0000;
    defparam \scaler_4.N_2725_i_l_ofx_LC_13_11_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \scaler_4.N_2725_i_l_ofx_LC_13_11_7  (
            .in0(_gnd_net_),
            .in1(N__53934),
            .in2(_gnd_net_),
            .in3(N__53910),
            .lcout(\scaler_4.N_2725_i_l_ofxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNISPTC1_8_LC_13_12_0 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNISPTC1_8_LC_13_12_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNISPTC1_8_LC_13_12_0 .LUT_INIT=16'b1000110011101111;
    LogicCell40 \pid_side.error_p_reg_esr_RNISPTC1_8_LC_13_12_0  (
            .in0(N__81229),
            .in1(N__84384),
            .in2(N__54026),
            .in3(N__54033),
            .lcout(\pid_side.error_p_reg_esr_RNISPTC1Z0Z_8 ),
            .ltout(\pid_side.error_p_reg_esr_RNISPTC1Z0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNIECBV6_8_LC_13_12_1 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIECBV6_8_LC_13_12_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIECBV6_8_LC_13_12_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pid_side.error_p_reg_esr_RNIECBV6_8_LC_13_12_1  (
            .in0(N__54041),
            .in1(N__69285),
            .in2(N__53874),
            .in3(N__66425),
            .lcout(\pid_side.error_p_reg_esr_RNIECBV6Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNIIAPH3_8_LC_13_12_2 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIIAPH3_8_LC_13_12_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIIAPH3_8_LC_13_12_2 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_side.error_p_reg_esr_RNIIAPH3_8_LC_13_12_2  (
            .in0(N__66426),
            .in1(N__54048),
            .in2(_gnd_net_),
            .in3(N__54042),
            .lcout(\pid_side.error_p_reg_esr_RNIIAPH3Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNI1VTC1_0_9_LC_13_12_3 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNI1VTC1_0_9_LC_13_12_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNI1VTC1_0_9_LC_13_12_3 .LUT_INIT=16'b0110100101100110;
    LogicCell40 \pid_side.error_p_reg_esr_RNI1VTC1_0_9_LC_13_12_3  (
            .in0(N__73013),
            .in1(N__80156),
            .in2(N__81170),
            .in3(N__53999),
            .lcout(\pid_side.error_p_reg_esr_RNI1VTC1_0Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI0UEI_8_LC_13_12_4 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI0UEI_8_LC_13_12_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI0UEI_8_LC_13_12_4 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI0UEI_8_LC_13_12_4  (
            .in0(_gnd_net_),
            .in1(N__53998),
            .in2(_gnd_net_),
            .in3(N__81162),
            .lcout(\pid_side.N_2374_i ),
            .ltout(\pid_side.N_2374_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNISPTC1_0_8_LC_13_12_5 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNISPTC1_0_8_LC_13_12_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNISPTC1_0_8_LC_13_12_5 .LUT_INIT=16'b0101101010010110;
    LogicCell40 \pid_side.error_p_reg_esr_RNISPTC1_0_8_LC_13_12_5  (
            .in0(N__84383),
            .in1(N__54019),
            .in2(N__54003),
            .in3(N__81228),
            .lcout(\pid_side.error_p_reg_esr_RNISPTC1_0Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_8_LC_13_12_6 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_8_LC_13_12_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_8_LC_13_12_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_8_LC_13_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81169),
            .lcout(\pid_side.error_d_reg_prevZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87027),
            .ce(N__83385),
            .sr(N__83183));
    defparam \pid_side.error_p_reg_esr_RNI1VTC1_9_LC_13_12_7 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNI1VTC1_9_LC_13_12_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNI1VTC1_9_LC_13_12_7 .LUT_INIT=16'b1101010011011101;
    LogicCell40 \pid_side.error_p_reg_esr_RNI1VTC1_9_LC_13_12_7  (
            .in0(N__73014),
            .in1(N__80157),
            .in2(N__81171),
            .in3(N__54000),
            .lcout(\pid_side.error_p_reg_esr_RNI1VTC1Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.state_0_LC_13_13_2 .C_ON=1'b0;
    defparam \pid_side.state_0_LC_13_13_2 .SEQ_MODE=4'b1000;
    defparam \pid_side.state_0_LC_13_13_2 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \pid_side.state_0_LC_13_13_2  (
            .in0(N__72587),
            .in1(N__59921),
            .in2(_gnd_net_),
            .in3(N__59849),
            .lcout(\pid_side.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87037),
            .ce(),
            .sr(N__79626));
    defparam \pid_side.error_cry_7_c_RNIRFCV2_LC_13_14_0 .C_ON=1'b0;
    defparam \pid_side.error_cry_7_c_RNIRFCV2_LC_13_14_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_7_c_RNIRFCV2_LC_13_14_0 .LUT_INIT=16'b0001010110110101;
    LogicCell40 \pid_side.error_cry_7_c_RNIRFCV2_LC_13_14_0  (
            .in0(N__80787),
            .in1(N__74072),
            .in2(N__80931),
            .in3(N__74188),
            .lcout(\pid_side.m36_1_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_0_22_LC_13_14_1 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_0_22_LC_13_14_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_0_22_LC_13_14_1 .LUT_INIT=16'b0010101011101010;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_0_22_LC_13_14_1  (
            .in0(N__74928),
            .in1(N__75704),
            .in2(N__71531),
            .in3(N__58428),
            .lcout(),
            .ltout(\pid_side.error_i_reg_esr_RNO_0Z0Z_22_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_22_LC_13_14_2 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_22_LC_13_14_2 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_esr_22_LC_13_14_2 .LUT_INIT=16'b1100100001000000;
    LogicCell40 \pid_side.error_i_reg_esr_22_LC_13_14_2  (
            .in0(N__76789),
            .in1(N__76639),
            .in2(N__53985),
            .in3(N__58434),
            .lcout(\pid_side.error_i_regZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87047),
            .ce(N__75305),
            .sr(N__79634));
    defparam \pid_side.error_cry_8_c_RNIVDRT4_LC_13_14_3 .C_ON=1'b0;
    defparam \pid_side.error_cry_8_c_RNIVDRT4_LC_13_14_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_8_c_RNIVDRT4_LC_13_14_3 .LUT_INIT=16'b1000100111001101;
    LogicCell40 \pid_side.error_cry_8_c_RNIVDRT4_LC_13_14_3  (
            .in0(N__72045),
            .in1(N__54075),
            .in2(N__74514),
            .in3(N__74420),
            .lcout(\pid_side.N_37_1 ),
            .ltout(\pid_side.N_37_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_8_c_RNIDO1S8_LC_13_14_4 .C_ON=1'b0;
    defparam \pid_side.error_cry_8_c_RNIDO1S8_LC_13_14_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_8_c_RNIDO1S8_LC_13_14_4 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \pid_side.error_cry_8_c_RNIDO1S8_LC_13_14_4  (
            .in0(_gnd_net_),
            .in1(N__71480),
            .in2(N__54069),
            .in3(N__62534),
            .lcout(\pid_side.N_39_1 ),
            .ltout(\pid_side.N_39_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_10_LC_13_14_5 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_10_LC_13_14_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_esr_10_LC_13_14_5 .LUT_INIT=16'b1000101000000010;
    LogicCell40 \pid_side.error_i_reg_esr_10_LC_13_14_5  (
            .in0(N__75508),
            .in1(N__75705),
            .in2(N__54066),
            .in3(N__54057),
            .lcout(\pid_side.error_i_regZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87047),
            .ce(N__75305),
            .sr(N__79634));
    defparam \pid_side.error_i_reg_esr_RNO_4_21_LC_13_14_6 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_4_21_LC_13_14_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_4_21_LC_13_14_6 .LUT_INIT=16'b0100000001111111;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_4_21_LC_13_14_6  (
            .in0(N__74421),
            .in1(N__72046),
            .in2(N__80796),
            .in3(N__74927),
            .lcout(),
            .ltout(\pid_side.N_126_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_0_21_LC_13_14_7 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_0_21_LC_13_14_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_0_21_LC_13_14_7 .LUT_INIT=16'b1100110111101111;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_0_21_LC_13_14_7  (
            .in0(N__71481),
            .in1(N__76788),
            .in2(N__54063),
            .in3(N__58557),
            .lcout(\pid_side.g1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_0_c_RNI5A3A1_LC_13_15_0 .C_ON=1'b0;
    defparam \pid_side.error_cry_0_c_RNI5A3A1_LC_13_15_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_0_c_RNI5A3A1_LC_13_15_0 .LUT_INIT=16'b0100010001000100;
    LogicCell40 \pid_side.error_cry_0_c_RNI5A3A1_LC_13_15_0  (
            .in0(N__80520),
            .in1(N__62307),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.N_55_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_0_c_RNI0KQ11_LC_13_15_1 .C_ON=1'b0;
    defparam \pid_side.error_cry_0_c_RNI0KQ11_LC_13_15_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_0_c_RNI0KQ11_LC_13_15_1 .LUT_INIT=16'b0100000001110011;
    LogicCell40 \pid_side.error_cry_0_c_RNI0KQ11_LC_13_15_1  (
            .in0(N__80786),
            .in1(N__80976),
            .in2(N__81067),
            .in3(N__62495),
            .lcout(\pid_side.m2_0_03_3_i_0 ),
            .ltout(\pid_side.m2_0_03_3_i_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_0_c_RNIN9TO4_LC_13_15_2 .C_ON=1'b0;
    defparam \pid_side.error_cry_0_c_RNIN9TO4_LC_13_15_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_0_c_RNIN9TO4_LC_13_15_2 .LUT_INIT=16'b1010000011110101;
    LogicCell40 \pid_side.error_cry_0_c_RNIN9TO4_LC_13_15_2  (
            .in0(N__80521),
            .in1(_gnd_net_),
            .in2(N__54060),
            .in3(N__62567),
            .lcout(\pid_side.N_41_0 ),
            .ltout(\pid_side.N_41_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_0_26_LC_13_15_3 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_0_26_LC_13_15_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_0_26_LC_13_15_3 .LUT_INIT=16'b1110001000000000;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_0_26_LC_13_15_3  (
            .in0(N__74924),
            .in1(N__76868),
            .in2(N__54051),
            .in3(N__76617),
            .lcout(),
            .ltout(\pid_side.error_i_reg_9_rn_0_26_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_26_LC_13_15_4 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_26_LC_13_15_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_esr_26_LC_13_15_4 .LUT_INIT=16'b0011000011111100;
    LogicCell40 \pid_side.error_i_reg_esr_26_LC_13_15_4  (
            .in0(_gnd_net_),
            .in1(N__68295),
            .in2(N__54099),
            .in3(N__54092),
            .lcout(\pid_side.error_i_regZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87057),
            .ce(N__75372),
            .sr(N__79643));
    defparam \pid_side.error_i_reg_esr_RNO_1_18_LC_13_15_5 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_1_18_LC_13_15_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_1_18_LC_13_15_5 .LUT_INIT=16'b0000000011010001;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_1_18_LC_13_15_5  (
            .in0(N__62568),
            .in1(N__80522),
            .in2(N__62317),
            .in3(N__80394),
            .lcout(),
            .ltout(\pid_side.m6_2_03_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_0_18_LC_13_15_6 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_0_18_LC_13_15_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_0_18_LC_13_15_6 .LUT_INIT=16'b1010001010000000;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_0_18_LC_13_15_6  (
            .in0(N__76616),
            .in1(N__76869),
            .in2(N__54096),
            .in3(N__74925),
            .lcout(),
            .ltout(\pid_side.error_i_reg_9_rn_0_18_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_18_LC_13_15_7 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_18_LC_13_15_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_esr_18_LC_13_15_7 .LUT_INIT=16'b0101010111110000;
    LogicCell40 \pid_side.error_i_reg_esr_18_LC_13_15_7  (
            .in0(N__54093),
            .in1(_gnd_net_),
            .in2(N__54084),
            .in3(N__71282),
            .lcout(\pid_side.error_i_regZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87057),
            .ce(N__75372),
            .sr(N__79643));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_5_LC_13_16_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_5_LC_13_16_0 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_5_LC_13_16_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_5_LC_13_16_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58829),
            .lcout(\dron_frame_decoder_1.drone_H_disp_side_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87064),
            .ce(N__54194),
            .sr(N__79650));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_6_LC_13_16_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_6_LC_13_16_1 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_6_LC_13_16_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_6_LC_13_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58742),
            .lcout(\dron_frame_decoder_1.drone_H_disp_side_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87064),
            .ce(N__54194),
            .sr(N__79650));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_7_LC_13_16_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_7_LC_13_16_2 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_7_LC_13_16_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_7_LC_13_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58651),
            .lcout(\dron_frame_decoder_1.drone_H_disp_side_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87064),
            .ce(N__54194),
            .sr(N__79650));
    defparam \pid_side.error_axb_2_LC_13_17_0 .C_ON=1'b0;
    defparam \pid_side.error_axb_2_LC_13_17_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_axb_2_LC_13_17_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_side.error_axb_2_LC_13_17_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54081),
            .lcout(\pid_side.error_axbZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_2_LC_13_17_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_2_LC_13_17_1 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_2_LC_13_17_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_2_LC_13_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59094),
            .lcout(drone_H_disp_side_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87076),
            .ce(N__54195),
            .sr(N__79658));
    defparam \pid_side.error_axb_3_LC_13_17_2 .C_ON=1'b0;
    defparam \pid_side.error_axb_3_LC_13_17_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_axb_3_LC_13_17_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_side.error_axb_3_LC_13_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54201),
            .lcout(\pid_side.error_axbZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_3_LC_13_17_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_3_LC_13_17_3 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_3_LC_13_17_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_3_LC_13_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59016),
            .lcout(drone_H_disp_side_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87076),
            .ce(N__54195),
            .sr(N__79658));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_0_LC_13_17_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_0_LC_13_17_4 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_0_LC_13_17_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_0_LC_13_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59318),
            .lcout(drone_H_disp_side_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87076),
            .ce(N__54195),
            .sr(N__79658));
    defparam \dron_frame_decoder_1.source_H_disp_side_fast_esr_0_LC_13_17_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_fast_esr_0_LC_13_17_5 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_fast_esr_0_LC_13_17_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_fast_esr_0_LC_13_17_5  (
            .in0(N__59319),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(dron_frame_decoder_1_source_H_disp_side_fast_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87076),
            .ce(N__54195),
            .sr(N__79658));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_1_LC_13_17_6 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_1_LC_13_17_6 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_1_LC_13_17_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_1_LC_13_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59197),
            .lcout(drone_H_disp_side_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87076),
            .ce(N__54195),
            .sr(N__79658));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_4_LC_13_17_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_4_LC_13_17_7 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_4_LC_13_17_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_4_LC_13_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58934),
            .lcout(\dron_frame_decoder_1.drone_H_disp_side_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87076),
            .ce(N__54195),
            .sr(N__79658));
    defparam \pid_alt.error_axb_2_LC_13_18_0 .C_ON=1'b0;
    defparam \pid_alt.error_axb_2_LC_13_18_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_axb_2_LC_13_18_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_alt.error_axb_2_LC_13_18_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54153),
            .lcout(\pid_alt.error_axbZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_2_LC_13_18_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_2_LC_13_18_1 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_2_LC_13_18_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_2_LC_13_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59093),
            .lcout(drone_altitude_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87089),
            .ce(N__54125),
            .sr(N__79665));
    defparam \pid_alt.error_axb_3_LC_13_18_2 .C_ON=1'b0;
    defparam \pid_alt.error_axb_3_LC_13_18_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_axb_3_LC_13_18_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_alt.error_axb_3_LC_13_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54135),
            .lcout(\pid_alt.error_axbZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_3_LC_13_18_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_3_LC_13_18_3 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_3_LC_13_18_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_3_LC_13_18_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59012),
            .lcout(drone_altitude_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87089),
            .ce(N__54125),
            .sr(N__79665));
    defparam \pid_front.error_axb_1_LC_13_18_4 .C_ON=1'b0;
    defparam \pid_front.error_axb_1_LC_13_18_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_axb_1_LC_13_18_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_front.error_axb_1_LC_13_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59112),
            .lcout(\pid_front.error_axbZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_axb_2_LC_13_18_5 .C_ON=1'b0;
    defparam \pid_front.error_axb_2_LC_13_18_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_axb_2_LC_13_18_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_front.error_axb_2_LC_13_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59031),
            .lcout(\pid_front.error_axbZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_axb_3_LC_13_18_6 .C_ON=1'b0;
    defparam \pid_front.error_axb_3_LC_13_18_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_axb_3_LC_13_18_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_front.error_axb_3_LC_13_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58941),
            .lcout(\pid_front.error_axbZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_axb_1_LC_13_18_7 .C_ON=1'b0;
    defparam \pid_side.error_axb_1_LC_13_18_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_axb_1_LC_13_18_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_side.error_axb_1_LC_13_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54384),
            .lcout(\pid_side.error_axbZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_xy_kd_2_LC_13_19_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_kd_2_LC_13_19_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_kd_2_LC_13_19_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_xy_kd_2_LC_13_19_2  (
            .in0(_gnd_net_),
            .in1(N__77573),
            .in2(_gnd_net_),
            .in3(N__86158),
            .lcout(xy_kd_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87105),
            .ce(N__84830),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_xy_kd_6_LC_13_19_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_kd_6_LC_13_19_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_kd_6_LC_13_19_5 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Commands_frame_decoder.source_xy_kd_6_LC_13_19_5  (
            .in0(N__86159),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73651),
            .lcout(xy_kd_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87105),
            .ce(N__84830),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIVIR9_11_LC_13_19_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIVIR9_11_LC_13_19_7 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIVIR9_11_LC_13_19_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_RNIVIR9_11_LC_13_19_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54324),
            .lcout(drone_altitude_i_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_esr_RNIH0C61_0_14_LC_13_20_2 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNIH0C61_0_14_LC_13_20_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNIH0C61_0_14_LC_13_20_2 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_front.error_p_reg_esr_RNIH0C61_0_14_LC_13_20_2  (
            .in0(N__54301),
            .in1(N__54270),
            .in2(_gnd_net_),
            .in3(N__82771),
            .lcout(\pid_front.error_p_reg_esr_RNIH0C61_0Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNIK7V3_4_LC_13_20_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNIK7V3_4_LC_13_20_3 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNIK7V3_4_LC_13_20_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_RNIK7V3_4_LC_13_20_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58848),
            .lcout(drone_H_disp_front_i_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNIL8V3_5_LC_13_20_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNIL8V3_5_LC_13_20_4 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNIL8V3_5_LC_13_20_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_RNIL8V3_5_LC_13_20_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58764),
            .lcout(drone_H_disp_front_i_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNIM9V3_6_LC_13_20_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNIM9V3_6_LC_13_20_5 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNIM9V3_6_LC_13_20_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_RNIM9V3_6_LC_13_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58665),
            .lcout(drone_H_disp_front_i_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNINAV3_7_LC_13_20_6 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNINAV3_7_LC_13_20_6 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNINAV3_7_LC_13_20_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_RNINAV3_7_LC_13_20_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58584),
            .lcout(drone_H_disp_front_i_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_axb_8_l_ofx_LC_13_20_7 .C_ON=1'b0;
    defparam \pid_front.error_axb_8_l_ofx_LC_13_20_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_axb_8_l_ofx_LC_13_20_7 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \pid_front.error_axb_8_l_ofx_LC_13_20_7  (
            .in0(N__54505),
            .in1(N__54476),
            .in2(_gnd_net_),
            .in3(N__54461),
            .lcout(\pid_front.error_axb_8_l_ofx_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_0_c_inv_LC_13_21_0 .C_ON=1'b1;
    defparam \pid_front.error_cry_0_c_inv_LC_13_21_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_0_c_inv_LC_13_21_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_front.error_cry_0_c_inv_LC_13_21_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__54447),
            .in3(N__59256),
            .lcout(\pid_front.error_axb_0 ),
            .ltout(),
            .carryin(bfn_13_21_0_),
            .carryout(\pid_front.error_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_0_c_RNIC7KB_LC_13_21_1 .C_ON=1'b1;
    defparam \pid_front.error_cry_0_c_RNIC7KB_LC_13_21_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_0_c_RNIC7KB_LC_13_21_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_front.error_cry_0_c_RNIC7KB_LC_13_21_1  (
            .in0(_gnd_net_),
            .in1(N__54438),
            .in2(_gnd_net_),
            .in3(N__54429),
            .lcout(\pid_front.error_1 ),
            .ltout(),
            .carryin(\pid_front.error_cry_0 ),
            .carryout(\pid_front.error_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_1_c_RNIEALB_LC_13_21_2 .C_ON=1'b1;
    defparam \pid_front.error_cry_1_c_RNIEALB_LC_13_21_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_1_c_RNIEALB_LC_13_21_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_front.error_cry_1_c_RNIEALB_LC_13_21_2  (
            .in0(_gnd_net_),
            .in1(N__54426),
            .in2(_gnd_net_),
            .in3(N__54417),
            .lcout(\pid_front.error_2 ),
            .ltout(),
            .carryin(\pid_front.error_cry_1 ),
            .carryout(\pid_front.error_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_2_c_RNIGDMB_LC_13_21_3 .C_ON=1'b1;
    defparam \pid_front.error_cry_2_c_RNIGDMB_LC_13_21_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_2_c_RNIGDMB_LC_13_21_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_front.error_cry_2_c_RNIGDMB_LC_13_21_3  (
            .in0(_gnd_net_),
            .in1(N__54414),
            .in2(_gnd_net_),
            .in3(N__54405),
            .lcout(\pid_front.error_3 ),
            .ltout(),
            .carryin(\pid_front.error_cry_2 ),
            .carryout(\pid_front.error_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_3_c_RNIABAG_LC_13_21_4 .C_ON=1'b1;
    defparam \pid_front.error_cry_3_c_RNIABAG_LC_13_21_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_3_c_RNIABAG_LC_13_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_cry_3_c_RNIABAG_LC_13_21_4  (
            .in0(_gnd_net_),
            .in1(N__54402),
            .in2(N__54396),
            .in3(N__54387),
            .lcout(\pid_front.error_4 ),
            .ltout(),
            .carryin(\pid_front.error_cry_3 ),
            .carryout(\pid_front.error_cry_0_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_0_0_c_RNIOQKB_LC_13_21_5 .C_ON=1'b1;
    defparam \pid_front.error_cry_0_0_c_RNIOQKB_LC_13_21_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_0_0_c_RNIOQKB_LC_13_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_cry_0_0_c_RNIOQKB_LC_13_21_5  (
            .in0(_gnd_net_),
            .in1(N__54651),
            .in2(N__54645),
            .in3(N__54636),
            .lcout(\pid_front.error_5 ),
            .ltout(),
            .carryin(\pid_front.error_cry_0_0 ),
            .carryout(\pid_front.error_cry_1_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_1_0_c_RNIR0RF_LC_13_21_6 .C_ON=1'b1;
    defparam \pid_front.error_cry_1_0_c_RNIR0RF_LC_13_21_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_1_0_c_RNIR0RF_LC_13_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_cry_1_0_c_RNIR0RF_LC_13_21_6  (
            .in0(_gnd_net_),
            .in1(N__54633),
            .in2(N__54627),
            .in3(N__54618),
            .lcout(\pid_front.error_6 ),
            .ltout(),
            .carryin(\pid_front.error_cry_1_0 ),
            .carryout(\pid_front.error_cry_2_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_2_0_c_RNIU61K_LC_13_21_7 .C_ON=1'b1;
    defparam \pid_front.error_cry_2_0_c_RNIU61K_LC_13_21_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_2_0_c_RNIU61K_LC_13_21_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_cry_2_0_c_RNIU61K_LC_13_21_7  (
            .in0(_gnd_net_),
            .in1(N__54615),
            .in2(N__54609),
            .in3(N__54600),
            .lcout(\pid_front.error_7 ),
            .ltout(),
            .carryin(\pid_front.error_cry_2_0 ),
            .carryout(\pid_front.error_cry_3_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_3_0_c_RNI1D7O_LC_13_22_0 .C_ON=1'b1;
    defparam \pid_front.error_cry_3_0_c_RNI1D7O_LC_13_22_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_3_0_c_RNI1D7O_LC_13_22_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_cry_3_0_c_RNI1D7O_LC_13_22_0  (
            .in0(_gnd_net_),
            .in1(N__54597),
            .in2(N__54591),
            .in3(N__54579),
            .lcout(\pid_front.error_8 ),
            .ltout(),
            .carryin(bfn_13_22_0_),
            .carryout(\pid_front.error_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_4_c_RNILNBG_LC_13_22_1 .C_ON=1'b1;
    defparam \pid_front.error_cry_4_c_RNILNBG_LC_13_22_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_4_c_RNILNBG_LC_13_22_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_cry_4_c_RNILNBG_LC_13_22_1  (
            .in0(_gnd_net_),
            .in1(N__54576),
            .in2(N__54570),
            .in3(N__54555),
            .lcout(\pid_front.error_9 ),
            .ltout(),
            .carryin(\pid_front.error_cry_4 ),
            .carryout(\pid_front.error_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_5_c_RNIVNFF_LC_13_22_2 .C_ON=1'b1;
    defparam \pid_front.error_cry_5_c_RNIVNFF_LC_13_22_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_5_c_RNIVNFF_LC_13_22_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_cry_5_c_RNIVNFF_LC_13_22_2  (
            .in0(_gnd_net_),
            .in1(N__54552),
            .in2(N__54543),
            .in3(N__54534),
            .lcout(\pid_front.error_10 ),
            .ltout(),
            .carryin(\pid_front.error_cry_5 ),
            .carryout(\pid_front.error_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_6_c_RNI3VJG_LC_13_22_3 .C_ON=1'b1;
    defparam \pid_front.error_cry_6_c_RNI3VJG_LC_13_22_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_6_c_RNI3VJG_LC_13_22_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_front.error_cry_6_c_RNI3VJG_LC_13_22_3  (
            .in0(_gnd_net_),
            .in1(N__54531),
            .in2(_gnd_net_),
            .in3(N__54519),
            .lcout(\pid_front.error_11 ),
            .ltout(),
            .carryin(\pid_front.error_cry_6 ),
            .carryout(\pid_front.error_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_7_c_RNIAPPM_LC_13_22_4 .C_ON=1'b1;
    defparam \pid_front.error_cry_7_c_RNIAPPM_LC_13_22_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_7_c_RNIAPPM_LC_13_22_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_cry_7_c_RNIAPPM_LC_13_22_4  (
            .in0(_gnd_net_),
            .in1(N__54516),
            .in2(N__54507),
            .in3(N__54483),
            .lcout(\pid_front.error_12 ),
            .ltout(),
            .carryin(\pid_front.error_cry_7 ),
            .carryout(\pid_front.error_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_8_c_RNIAC2E_LC_13_22_5 .C_ON=1'b1;
    defparam \pid_front.error_cry_8_c_RNIAC2E_LC_13_22_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_8_c_RNIAC2E_LC_13_22_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_cry_8_c_RNIAC2E_LC_13_22_5  (
            .in0(_gnd_net_),
            .in1(N__54909),
            .in2(N__54897),
            .in3(N__54882),
            .lcout(\pid_front.error_13 ),
            .ltout(),
            .carryin(\pid_front.error_cry_8 ),
            .carryout(\pid_front.error_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_9_c_RNIDG3E_LC_13_22_6 .C_ON=1'b1;
    defparam \pid_front.error_cry_9_c_RNIDG3E_LC_13_22_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_9_c_RNIDG3E_LC_13_22_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_cry_9_c_RNIDG3E_LC_13_22_6  (
            .in0(_gnd_net_),
            .in1(N__54879),
            .in2(N__54864),
            .in3(N__54873),
            .lcout(\pid_front.error_14 ),
            .ltout(),
            .carryin(\pid_front.error_cry_9 ),
            .carryout(\pid_front.error_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_10_c_RNINTDI_LC_13_22_7 .C_ON=1'b0;
    defparam \pid_front.error_cry_10_c_RNINTDI_LC_13_22_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_10_c_RNINTDI_LC_13_22_7 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_front.error_cry_10_c_RNINTDI_LC_13_22_7  (
            .in0(N__54870),
            .in1(N__54863),
            .in2(_gnd_net_),
            .in3(N__54852),
            .lcout(\pid_front.error_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNII1MD_0_LC_13_23_0 .C_ON=1'b1;
    defparam \pid_front.error_i_reg_esr_RNII1MD_0_LC_13_23_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNII1MD_0_LC_13_23_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \pid_front.error_i_reg_esr_RNII1MD_0_LC_13_23_0  (
            .in0(_gnd_net_),
            .in1(N__56129),
            .in2(N__62879),
            .in3(_gnd_net_),
            .lcout(\pid_front.un1_pid_prereg_0 ),
            .ltout(),
            .carryin(bfn_13_23_0_),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_0_c_RNI9AGE_LC_13_23_1 .C_ON=1'b1;
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_0_c_RNI9AGE_LC_13_23_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_0_c_RNI9AGE_LC_13_23_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_0_c_RNI9AGE_LC_13_23_1  (
            .in0(_gnd_net_),
            .in1(N__54819),
            .in2(N__70836),
            .in3(N__54774),
            .lcout(\pid_front.un1_error_i_acumm_prereg_cry_0_c_RNI9AGE ),
            .ltout(),
            .carryin(\pid_front.un1_error_i_acumm_prereg_cry_0 ),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_1_c_RNICEHE_LC_13_23_2 .C_ON=1'b1;
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_1_c_RNICEHE_LC_13_23_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_1_c_RNICEHE_LC_13_23_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_1_c_RNICEHE_LC_13_23_2  (
            .in0(_gnd_net_),
            .in1(N__54771),
            .in2(N__62742),
            .in3(N__54726),
            .lcout(\pid_front.un1_error_i_acumm_prereg_cry_1_c_RNICEHE ),
            .ltout(),
            .carryin(\pid_front.un1_error_i_acumm_prereg_cry_1 ),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_2_c_RNIFIIE_LC_13_23_3 .C_ON=1'b1;
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_2_c_RNIFIIE_LC_13_23_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_2_c_RNIFIIE_LC_13_23_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_2_c_RNIFIIE_LC_13_23_3  (
            .in0(_gnd_net_),
            .in1(N__54723),
            .in2(N__62727),
            .in3(N__54693),
            .lcout(\pid_front.un1_error_i_acumm_prereg_cry_2_c_RNIFIIE ),
            .ltout(),
            .carryin(\pid_front.un1_error_i_acumm_prereg_cry_2 ),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_3_c_RNIIMJE_LC_13_23_4 .C_ON=1'b1;
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_3_c_RNIIMJE_LC_13_23_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_3_c_RNIIMJE_LC_13_23_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_3_c_RNIIMJE_LC_13_23_4  (
            .in0(_gnd_net_),
            .in1(N__54690),
            .in2(N__68217),
            .in3(N__54654),
            .lcout(\pid_front.un1_error_i_acumm_prereg_cry_3_c_RNIIMJE ),
            .ltout(),
            .carryin(\pid_front.un1_error_i_acumm_prereg_cry_3 ),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_4_c_RNICGQM_LC_13_23_5 .C_ON=1'b1;
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_4_c_RNICGQM_LC_13_23_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_4_c_RNICGQM_LC_13_23_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_4_c_RNICGQM_LC_13_23_5  (
            .in0(_gnd_net_),
            .in1(N__55224),
            .in2(N__55218),
            .in3(N__55161),
            .lcout(\pid_front.un1_error_i_acumm_prereg_cry_4_c_RNICGQM ),
            .ltout(),
            .carryin(\pid_front.un1_error_i_acumm_prereg_cry_4 ),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_5_c_RNIOULE_LC_13_23_6 .C_ON=1'b1;
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_5_c_RNIOULE_LC_13_23_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_5_c_RNIOULE_LC_13_23_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_5_c_RNIOULE_LC_13_23_6  (
            .in0(_gnd_net_),
            .in1(N__55158),
            .in2(N__67917),
            .in3(N__55125),
            .lcout(\pid_front.un1_error_i_acumm_prereg_cry_5_c_RNIOULE ),
            .ltout(),
            .carryin(\pid_front.un1_error_i_acumm_prereg_cry_5 ),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_6_c_RNIR2NE_LC_13_23_7 .C_ON=1'b1;
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_6_c_RNIR2NE_LC_13_23_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_6_c_RNIR2NE_LC_13_23_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_6_c_RNIR2NE_LC_13_23_7  (
            .in0(_gnd_net_),
            .in1(N__55122),
            .in2(N__67896),
            .in3(N__55092),
            .lcout(\pid_front.un1_error_i_acumm_prereg_cry_6_c_RNIR2NE ),
            .ltout(),
            .carryin(\pid_front.un1_error_i_acumm_prereg_cry_6 ),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_7_c_RNIU6OE_LC_13_24_0 .C_ON=1'b1;
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_7_c_RNIU6OE_LC_13_24_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_7_c_RNIU6OE_LC_13_24_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_7_c_RNIU6OE_LC_13_24_0  (
            .in0(_gnd_net_),
            .in1(N__55089),
            .in2(N__68052),
            .in3(N__55056),
            .lcout(\pid_front.un1_error_i_acumm_prereg_cry_7_c_RNIU6OE ),
            .ltout(),
            .carryin(bfn_13_24_0_),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_8_c_RNI1BPE_LC_13_24_1 .C_ON=1'b1;
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_8_c_RNI1BPE_LC_13_24_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_8_c_RNI1BPE_LC_13_24_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_8_c_RNI1BPE_LC_13_24_1  (
            .in0(_gnd_net_),
            .in1(N__55053),
            .in2(N__68127),
            .in3(N__55017),
            .lcout(\pid_front.un1_error_i_acumm_prereg_cry_8_c_RNI1BPE ),
            .ltout(),
            .carryin(\pid_front.un1_error_i_acumm_prereg_cry_8 ),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_9_c_RNIIPQK_LC_13_24_2 .C_ON=1'b1;
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_9_c_RNIIPQK_LC_13_24_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_9_c_RNIIPQK_LC_13_24_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_9_c_RNIIPQK_LC_13_24_2  (
            .in0(_gnd_net_),
            .in1(N__55014),
            .in2(N__59601),
            .in3(N__54981),
            .lcout(\pid_front.un1_error_i_acumm_prereg_cry_9_c_RNIIPQK ),
            .ltout(),
            .carryin(\pid_front.un1_error_i_acumm_prereg_cry_9 ),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_10_c_RNIJD4S_LC_13_24_3 .C_ON=1'b1;
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_10_c_RNIJD4S_LC_13_24_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_10_c_RNIJD4S_LC_13_24_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_10_c_RNIJD4S_LC_13_24_3  (
            .in0(_gnd_net_),
            .in1(N__54978),
            .in2(N__67494),
            .in3(N__54942),
            .lcout(\pid_front.un1_error_i_acumm_prereg_cry_10_c_RNIJD4S ),
            .ltout(),
            .carryin(\pid_front.un1_error_i_acumm_prereg_cry_10 ),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNIV4AU_12_LC_13_24_4 .C_ON=1'b1;
    defparam \pid_front.error_i_reg_esr_RNIV4AU_12_LC_13_24_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNIV4AU_12_LC_13_24_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_i_reg_esr_RNIV4AU_12_LC_13_24_4  (
            .in0(_gnd_net_),
            .in1(N__54939),
            .in2(N__59490),
            .in3(N__54912),
            .lcout(\pid_front.error_i_reg_esr_RNIV4AUZ0Z_12 ),
            .ltout(),
            .carryin(\pid_front.un1_error_i_acumm_prereg_cry_11 ),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNI29BU_13_LC_13_24_5 .C_ON=1'b1;
    defparam \pid_front.error_i_reg_esr_RNI29BU_13_LC_13_24_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNI29BU_13_LC_13_24_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_i_reg_esr_RNI29BU_13_LC_13_24_5  (
            .in0(_gnd_net_),
            .in1(N__55558),
            .in2(N__68001),
            .in3(N__55422),
            .lcout(\pid_front.error_i_reg_esr_RNI29BUZ0Z_13 ),
            .ltout(),
            .carryin(\pid_front.un1_error_i_acumm_prereg_cry_12 ),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNI4CCU_14_LC_13_24_6 .C_ON=1'b1;
    defparam \pid_front.error_i_reg_esr_RNI4CCU_14_LC_13_24_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNI4CCU_14_LC_13_24_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_i_reg_esr_RNI4CCU_14_LC_13_24_6  (
            .in0(_gnd_net_),
            .in1(N__59565),
            .in2(N__55590),
            .in3(N__55383),
            .lcout(\pid_front.error_i_reg_esr_RNI4CCUZ0Z_14 ),
            .ltout(),
            .carryin(\pid_front.un1_error_i_acumm_prereg_cry_13 ),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNI6FDU_15_LC_13_24_7 .C_ON=1'b1;
    defparam \pid_front.error_i_reg_esr_RNI6FDU_15_LC_13_24_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNI6FDU_15_LC_13_24_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_i_reg_esr_RNI6FDU_15_LC_13_24_7  (
            .in0(_gnd_net_),
            .in1(N__55562),
            .in2(N__70794),
            .in3(N__55353),
            .lcout(\pid_front.error_i_reg_esr_RNI6FDUZ0Z_15 ),
            .ltout(),
            .carryin(\pid_front.un1_error_i_acumm_prereg_cry_14 ),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNI8IEU_16_LC_13_25_0 .C_ON=1'b1;
    defparam \pid_front.error_i_reg_esr_RNI8IEU_16_LC_13_25_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNI8IEU_16_LC_13_25_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_i_reg_esr_RNI8IEU_16_LC_13_25_0  (
            .in0(_gnd_net_),
            .in1(N__55563),
            .in2(N__59352),
            .in3(N__55326),
            .lcout(\pid_front.error_i_reg_esr_RNI8IEUZ0Z_16 ),
            .ltout(),
            .carryin(bfn_13_25_0_),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNIALFU_17_LC_13_25_1 .C_ON=1'b1;
    defparam \pid_front.error_i_reg_esr_RNIALFU_17_LC_13_25_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNIALFU_17_LC_13_25_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_i_reg_esr_RNIALFU_17_LC_13_25_1  (
            .in0(_gnd_net_),
            .in1(N__72435),
            .in2(N__55591),
            .in3(N__55323),
            .lcout(\pid_front.error_i_reg_esr_RNIALFUZ0Z_17 ),
            .ltout(),
            .carryin(\pid_front.un1_error_i_acumm_prereg_cry_16 ),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNICOGU_18_LC_13_25_2 .C_ON=1'b1;
    defparam \pid_front.error_i_reg_esr_RNICOGU_18_LC_13_25_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNICOGU_18_LC_13_25_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_i_reg_esr_RNICOGU_18_LC_13_25_2  (
            .in0(_gnd_net_),
            .in1(N__55567),
            .in2(N__59481),
            .in3(N__55290),
            .lcout(\pid_front.error_i_reg_esr_RNICOGUZ0Z_18 ),
            .ltout(),
            .carryin(\pid_front.un1_error_i_acumm_prereg_cry_17 ),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNIERHU_19_LC_13_25_3 .C_ON=1'b1;
    defparam \pid_front.error_i_reg_esr_RNIERHU_19_LC_13_25_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNIERHU_19_LC_13_25_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_i_reg_esr_RNIERHU_19_LC_13_25_3  (
            .in0(_gnd_net_),
            .in1(N__67968),
            .in2(N__55592),
            .in3(N__55254),
            .lcout(\pid_front.error_i_reg_esr_RNIERHUZ0Z_19 ),
            .ltout(),
            .carryin(\pid_front.un1_error_i_acumm_prereg_cry_18 ),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNI7MJU_20_LC_13_25_4 .C_ON=1'b1;
    defparam \pid_front.error_i_reg_esr_RNI7MJU_20_LC_13_25_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNI7MJU_20_LC_13_25_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_i_reg_esr_RNI7MJU_20_LC_13_25_4  (
            .in0(_gnd_net_),
            .in1(N__55571),
            .in2(N__63036),
            .in3(N__55227),
            .lcout(\pid_front.error_i_reg_esr_RNI7MJUZ0Z_20 ),
            .ltout(),
            .carryin(\pid_front.un1_error_i_acumm_prereg_cry_19 ),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNI08DV_21_LC_13_25_5 .C_ON=1'b1;
    defparam \pid_front.error_i_reg_esr_RNI08DV_21_LC_13_25_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNI08DV_21_LC_13_25_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_i_reg_esr_RNI08DV_21_LC_13_25_5  (
            .in0(_gnd_net_),
            .in1(N__59496),
            .in2(N__55593),
            .in3(N__55698),
            .lcout(\pid_front.error_i_reg_esr_RNI08DVZ0Z_21 ),
            .ltout(),
            .carryin(\pid_front.un1_error_i_acumm_prereg_cry_20 ),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNI2BEV_22_LC_13_25_6 .C_ON=1'b1;
    defparam \pid_front.error_i_reg_esr_RNI2BEV_22_LC_13_25_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNI2BEV_22_LC_13_25_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_i_reg_esr_RNI2BEV_22_LC_13_25_6  (
            .in0(_gnd_net_),
            .in1(N__55575),
            .in2(N__59544),
            .in3(N__55671),
            .lcout(\pid_front.error_i_reg_esr_RNI2BEVZ0Z_22 ),
            .ltout(),
            .carryin(\pid_front.un1_error_i_acumm_prereg_cry_21 ),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNI4EFV_23_LC_13_25_7 .C_ON=1'b1;
    defparam \pid_front.error_i_reg_esr_RNI4EFV_23_LC_13_25_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNI4EFV_23_LC_13_25_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_i_reg_esr_RNI4EFV_23_LC_13_25_7  (
            .in0(_gnd_net_),
            .in1(N__71328),
            .in2(N__55594),
            .in3(N__55668),
            .lcout(\pid_front.error_i_reg_esr_RNI4EFVZ0Z_23 ),
            .ltout(),
            .carryin(\pid_front.un1_error_i_acumm_prereg_cry_22 ),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNI6HGV_24_LC_13_26_0 .C_ON=1'b1;
    defparam \pid_front.error_i_reg_esr_RNI6HGV_24_LC_13_26_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNI6HGV_24_LC_13_26_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_i_reg_esr_RNI6HGV_24_LC_13_26_0  (
            .in0(_gnd_net_),
            .in1(N__55595),
            .in2(N__63192),
            .in3(N__55641),
            .lcout(\pid_front.error_i_reg_esr_RNI6HGVZ0Z_24 ),
            .ltout(),
            .carryin(bfn_13_26_0_),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNI8KHV_25_LC_13_26_1 .C_ON=1'b1;
    defparam \pid_front.error_i_reg_esr_RNI8KHV_25_LC_13_26_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNI8KHV_25_LC_13_26_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_i_reg_esr_RNI8KHV_25_LC_13_26_1  (
            .in0(_gnd_net_),
            .in1(N__68082),
            .in2(N__55604),
            .in3(N__55638),
            .lcout(\pid_front.error_i_reg_esr_RNI8KHVZ0Z_25 ),
            .ltout(),
            .carryin(\pid_front.un1_error_i_acumm_prereg_cry_24 ),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNIANIV_26_LC_13_26_2 .C_ON=1'b1;
    defparam \pid_front.error_i_reg_esr_RNIANIV_26_LC_13_26_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNIANIV_26_LC_13_26_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_i_reg_esr_RNIANIV_26_LC_13_26_2  (
            .in0(_gnd_net_),
            .in1(N__55599),
            .in2(N__63957),
            .in3(N__55611),
            .lcout(\pid_front.error_i_reg_esr_RNIANIVZ0Z_26 ),
            .ltout(),
            .carryin(\pid_front.un1_error_i_acumm_prereg_cry_25 ),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_26_c_RNICQJV_LC_13_26_3 .C_ON=1'b1;
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_26_c_RNICQJV_LC_13_26_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_26_c_RNICQJV_LC_13_26_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_26_c_RNICQJV_LC_13_26_3  (
            .in0(_gnd_net_),
            .in1(N__67988),
            .in2(N__55605),
            .in3(N__55608),
            .lcout(\pid_front.un1_error_i_acumm_prereg_cry_26_c_RNICQJV ),
            .ltout(),
            .carryin(\pid_front.un1_error_i_acumm_prereg_cry_26 ),
            .carryout(\pid_front.un1_error_i_acumm_prereg_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_27_c_RNIDSKV_LC_13_26_4 .C_ON=1'b0;
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_27_c_RNIDSKV_LC_13_26_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_27_c_RNIDSKV_LC_13_26_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_front.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_27_c_RNIDSKV_LC_13_26_4  (
            .in0(N__67989),
            .in1(N__55603),
            .in2(_gnd_net_),
            .in3(N__55524),
            .lcout(\pid_front.un1_error_i_acumm_prereg_cry_27_c_RNIDSKV ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_acumm_prereg_esr_28_LC_13_26_5 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_28_LC_13_26_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_28_LC_13_26_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_28_LC_13_26_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55511),
            .lcout(\pid_front.error_i_acumm_preregZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87214),
            .ce(N__56082),
            .sr(N__79701));
    defparam \pid_front.error_i_acumm_prereg_esr_25_LC_13_27_0 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_25_LC_13_27_0 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_25_LC_13_27_0 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_25_LC_13_27_0  (
            .in0(_gnd_net_),
            .in1(N__56279),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_i_acumm_preregZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87227),
            .ce(N__56080),
            .sr(N__79705));
    defparam \pid_front.error_i_acumm_prereg_esr_23_LC_13_27_3 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_23_LC_13_27_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_23_LC_13_27_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_23_LC_13_27_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56251),
            .lcout(\pid_front.error_i_acumm_preregZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87227),
            .ce(N__56080),
            .sr(N__79705));
    defparam \pid_front.error_i_acumm_prereg_esr_27_LC_13_27_4 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_27_LC_13_27_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_27_LC_13_27_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_27_LC_13_27_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56198),
            .lcout(\pid_front.error_i_acumm_preregZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87227),
            .ce(N__56080),
            .sr(N__79705));
    defparam \pid_front.error_i_acumm_prereg_esr_17_LC_13_27_5 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_17_LC_13_27_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_17_LC_13_27_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_17_LC_13_27_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56175),
            .lcout(\pid_front.error_i_acumm_preregZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87227),
            .ce(N__56080),
            .sr(N__79705));
    defparam \pid_front.error_i_acumm_prereg_esr_0_LC_13_28_4 .C_ON=1'b0;
    defparam \pid_front.error_i_acumm_prereg_esr_0_LC_13_28_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_acumm_prereg_esr_0_LC_13_28_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_front.error_i_acumm_prereg_esr_0_LC_13_28_4  (
            .in0(_gnd_net_),
            .in1(N__62883),
            .in2(_gnd_net_),
            .in3(N__56139),
            .lcout(\pid_front.error_i_acumm_preregZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87241),
            .ce(N__56078),
            .sr(N__79710));
    defparam \pid_alt.state_RNIH1EN_0_LC_13_29_6 .C_ON=1'b0;
    defparam \pid_alt.state_RNIH1EN_0_LC_13_29_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.state_RNIH1EN_0_LC_13_29_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \pid_alt.state_RNIH1EN_0_LC_13_29_6  (
            .in0(_gnd_net_),
            .in1(N__56037),
            .in2(_gnd_net_),
            .in3(N__79934),
            .lcout(\pid_alt.state_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_0_LC_14_1_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_0_LC_14_1_5 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_0_LC_14_1_5 .LUT_INIT=16'b0000000010101100;
    LogicCell40 \ppm_encoder_1.init_pulses_0_LC_14_1_5  (
            .in0(N__55980),
            .in1(N__55965),
            .in2(N__55954),
            .in3(N__55827),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__86970),
            .ce(),
            .sr(N__79564));
    defparam \ppm_encoder_1.counter24_0_I_1_c_LC_14_2_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_1_c_LC_14_2_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_1_c_LC_14_2_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_1_c_LC_14_2_0  (
            .in0(_gnd_net_),
            .in1(N__64731),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_2_0_),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_9_c_LC_14_2_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_9_c_LC_14_2_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_9_c_LC_14_2_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_9_c_LC_14_2_1  (
            .in0(_gnd_net_),
            .in1(N__60276),
            .in2(N__56635),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ppm_encoder_1.counter24_0_data_tmp_0 ),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_15_c_LC_14_2_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_15_c_LC_14_2_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_15_c_LC_14_2_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_15_c_LC_14_2_2  (
            .in0(_gnd_net_),
            .in1(N__56595),
            .in2(N__59784),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ppm_encoder_1.counter24_0_data_tmp_1 ),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_21_c_LC_14_2_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_21_c_LC_14_2_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_21_c_LC_14_2_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_21_c_LC_14_2_3  (
            .in0(_gnd_net_),
            .in1(N__57879),
            .in2(N__56632),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ppm_encoder_1.counter24_0_data_tmp_2 ),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_27_c_LC_14_2_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_27_c_LC_14_2_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_27_c_LC_14_2_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_27_c_LC_14_2_4  (
            .in0(_gnd_net_),
            .in1(N__60270),
            .in2(N__56636),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ppm_encoder_1.counter24_0_data_tmp_3 ),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_33_c_LC_14_2_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_33_c_LC_14_2_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_33_c_LC_14_2_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_33_c_LC_14_2_5  (
            .in0(_gnd_net_),
            .in1(N__60525),
            .in2(N__56633),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ppm_encoder_1.counter24_0_data_tmp_4 ),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_39_c_LC_14_2_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_39_c_LC_14_2_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_39_c_LC_14_2_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_39_c_LC_14_2_6  (
            .in0(_gnd_net_),
            .in1(N__60384),
            .in2(N__56637),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ppm_encoder_1.counter24_0_data_tmp_5 ),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_45_c_LC_14_2_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_45_c_LC_14_2_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_45_c_LC_14_2_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_45_c_LC_14_2_7  (
            .in0(_gnd_net_),
            .in1(N__68493),
            .in2(N__56634),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ppm_encoder_1.counter24_0_data_tmp_6 ),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_51_c_LC_14_3_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_51_c_LC_14_3_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_51_c_LC_14_3_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_51_c_LC_14_3_0  (
            .in0(_gnd_net_),
            .in1(N__64314),
            .in2(N__56631),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_3_0_),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_57_c_LC_14_3_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_57_c_LC_14_3_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_57_c_LC_14_3_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_57_c_LC_14_3_1  (
            .in0(_gnd_net_),
            .in1(N__56594),
            .in2(N__56754),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ppm_encoder_1.counter24_0_data_tmp_8 ),
            .carryout(\ppm_encoder_1.counter24_0_N_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_N_2_THRU_LUT4_0_LC_14_3_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_N_2_THRU_LUT4_0_LC_14_3_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_N_2_THRU_LUT4_0_LC_14_3_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.counter24_0_N_2_THRU_LUT4_0_LC_14_3_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56820),
            .lcout(\ppm_encoder_1.counter24_0_N_2_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_10_LC_14_3_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_10_LC_14_3_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_10_LC_14_3_3 .LUT_INIT=16'b0001000010110000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_10_LC_14_3_3  (
            .in0(N__61638),
            .in1(N__56817),
            .in2(N__61447),
            .in3(N__56787),
            .lcout(\ppm_encoder_1.pulses2count_9_i_0_1_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNO_LC_14_3_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNO_LC_14_3_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNO_LC_14_3_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ppm_encoder_1.counter24_0_I_57_c_RNO_LC_14_3_4  (
            .in0(_gnd_net_),
            .in1(N__60585),
            .in2(_gnd_net_),
            .in3(N__65514),
            .lcout(\ppm_encoder_1.counter24_0_I_57_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNI7A1R_1_LC_14_3_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI7A1R_1_LC_14_3_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI7A1R_1_LC_14_3_5 .LUT_INIT=16'b1111000001111000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI7A1R_1_LC_14_3_5  (
            .in0(N__57681),
            .in1(N__57262),
            .in2(N__63690),
            .in3(N__64148),
            .lcout(\ppm_encoder_1.N_258_i_i ),
            .ltout(\ppm_encoder_1.N_258_i_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNI40GS4_1_LC_14_3_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI40GS4_1_LC_14_3_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI40GS4_1_LC_14_3_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI40GS4_1_LC_14_3_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__56733),
            .in3(N__56673),
            .lcout(\ppm_encoder_1.init_pulses_RNI40GS4Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_7_LC_14_3_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_7_LC_14_3_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_7_LC_14_3_7 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_7_LC_14_3_7  (
            .in0(_gnd_net_),
            .in1(N__64444),
            .in2(_gnd_net_),
            .in3(N__56721),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_2Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.PPM_STATE_RNI5C4L_1_LC_14_4_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_RNI5C4L_1_LC_14_4_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.PPM_STATE_RNI5C4L_1_LC_14_4_0 .LUT_INIT=16'b1111111111011111;
    LogicCell40 \ppm_encoder_1.PPM_STATE_RNI5C4L_1_LC_14_4_0  (
            .in0(N__57257),
            .in1(N__61204),
            .in2(N__57689),
            .in3(N__61137),
            .lcout(\ppm_encoder_1.PPM_STATE_RNI5C4LZ0Z_1 ),
            .ltout(\ppm_encoder_1.PPM_STATE_RNI5C4LZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNI7A1R_0_1_LC_14_4_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI7A1R_0_1_LC_14_4_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI7A1R_0_1_LC_14_4_1 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI7A1R_0_1_LC_14_4_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__56685),
            .in3(N__63675),
            .lcout(),
            .ltout(\ppm_encoder_1.init_pulses_RNI7A1R_0Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNITLE14_1_LC_14_4_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNITLE14_1_LC_14_4_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNITLE14_1_LC_14_4_2 .LUT_INIT=16'b0000111100011110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNITLE14_1_LC_14_4_2  (
            .in0(N__57888),
            .in1(N__56682),
            .in2(N__56676),
            .in3(N__57039),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_axb_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_2_LC_14_4_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_2_LC_14_4_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_2_LC_14_4_4 .LUT_INIT=16'b0000000010110001;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_2_LC_14_4_4  (
            .in0(N__64165),
            .in1(N__57406),
            .in2(N__57266),
            .in3(N__79980),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__86980),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIDUME1_11_LC_14_4_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIDUME1_11_LC_14_4_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIDUME1_11_LC_14_4_5 .LUT_INIT=16'b0011101100001010;
    LogicCell40 \ppm_encoder_1.throttle_RNIDUME1_11_LC_14_4_5  (
            .in0(N__57983),
            .in1(N__60299),
            .in2(N__57378),
            .in3(N__57151),
            .lcout(\ppm_encoder_1.un2_throttle_iv_0_1_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_3_rep1_LC_14_4_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_3_rep1_LC_14_4_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_3_rep1_LC_14_4_6 .LUT_INIT=16'b0000000010110001;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_3_rep1_LC_14_4_6  (
            .in0(N__64164),
            .in1(N__63908),
            .in2(N__57690),
            .in3(N__79979),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_3_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__86980),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_0_LC_14_4_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_0_LC_14_4_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_0_LC_14_4_7 .LUT_INIT=16'b1111101011101110;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_0_LC_14_4_7  (
            .in0(N__79978),
            .in1(N__57436),
            .in2(N__57216),
            .in3(N__64166),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__86980),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIM4C21_2_LC_14_5_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIM4C21_2_LC_14_5_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIM4C21_2_LC_14_5_0 .LUT_INIT=16'b1111111110011101;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIM4C21_2_LC_14_5_0  (
            .in0(N__57679),
            .in1(N__57254),
            .in2(N__63847),
            .in3(N__64102),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIM4C21Z0Z_2 ),
            .ltout(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIM4C21Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIN1203_2_LC_14_5_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIN1203_2_LC_14_5_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIN1203_2_LC_14_5_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIN1203_2_LC_14_5_1  (
            .in0(N__56864),
            .in1(N__63231),
            .in2(N__57288),
            .in3(N__57625),
            .lcout(\ppm_encoder_1.init_pulses_RNIN1203Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIIP7D_0_LC_14_5_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIIP7D_0_LC_14_5_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIIP7D_0_LC_14_5_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIIP7D_0_LC_14_5_2  (
            .in0(_gnd_net_),
            .in1(N__57253),
            .in2(_gnd_net_),
            .in3(N__57211),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIIP7DZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNIN3K62_2_LC_14_5_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNIN3K62_2_LC_14_5_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNIN3K62_2_LC_14_5_3 .LUT_INIT=16'b1111111110101011;
    LogicCell40 \ppm_encoder_1.elevator_RNIN3K62_2_LC_14_5_3  (
            .in0(N__63789),
            .in1(N__63555),
            .in2(N__58067),
            .in3(N__57009),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_2_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNICULF4_2_LC_14_5_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNICULF4_2_LC_14_5_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNICULF4_2_LC_14_5_4 .LUT_INIT=16'b1100100100110110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNICULF4_2_LC_14_5_4  (
            .in0(N__56958),
            .in1(N__63240),
            .in2(N__56952),
            .in3(N__56863),
            .lcout(),
            .ltout(\ppm_encoder_1.un1_init_pulses_0_axb_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNI5GAI5_2_LC_14_5_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI5GAI5_2_LC_14_5_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI5GAI5_2_LC_14_5_5 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI5GAI5_2_LC_14_5_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__57726),
            .in3(N__57624),
            .lcout(\ppm_encoder_1.init_pulses_RNI5GAI5Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIPHK21_2_LC_14_5_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIPHK21_2_LC_14_5_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIPHK21_2_LC_14_5_6 .LUT_INIT=16'b1111000001111000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIPHK21_2_LC_14_5_6  (
            .in0(N__57680),
            .in1(N__63788),
            .in2(N__63236),
            .in3(N__64103),
            .lcout(\ppm_encoder_1.N_259_i_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_1_LC_14_5_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_1_LC_14_5_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_1_LC_14_5_7 .LUT_INIT=16'b0010001100010000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_1_LC_14_5_7  (
            .in0(N__64104),
            .in1(N__79986),
            .in2(N__61628),
            .in3(N__57601),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__86986),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_14_LC_14_6_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_14_LC_14_6_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_14_LC_14_6_0 .LUT_INIT=16'b0000001001010010;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_14_LC_14_6_0  (
            .in0(N__61637),
            .in1(N__57572),
            .in2(N__61457),
            .in3(N__57540),
            .lcout(),
            .ltout(\ppm_encoder_1.pulses2count_9_i_0_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_14_LC_14_6_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_14_LC_14_6_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_14_LC_14_6_1 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_14_LC_14_6_1  (
            .in0(N__61840),
            .in1(_gnd_net_),
            .in2(N__57513),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\ppm_encoder_1.pulses2count_9_i_1_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_14_LC_14_6_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_14_LC_14_6_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_14_LC_14_6_2 .LUT_INIT=16'b0000000000001101;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_14_LC_14_6_2  (
            .in0(N__64441),
            .in1(N__57510),
            .in2(N__57477),
            .in3(N__57474),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__86994),
            .ce(N__68751),
            .sr(N__79592));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_1_LC_14_6_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_1_LC_14_6_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_1_LC_14_6_3 .LUT_INIT=16'b1010000000001100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_1_LC_14_6_3  (
            .in0(N__58035),
            .in1(N__63460),
            .in2(N__61641),
            .in3(N__61443),
            .lcout(\ppm_encoder_1.pulses2count_9_0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m2_0_a2_0_a2_LC_14_6_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m2_0_a2_0_a2_LC_14_6_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m2_0_a2_0_a2_LC_14_6_4 .LUT_INIT=16'b0001000100110011;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m2_0_a2_0_a2_LC_14_6_4  (
            .in0(N__63459),
            .in1(N__61633),
            .in2(_gnd_net_),
            .in3(N__64600),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_ns_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNIC2521_3_LC_14_6_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNIC2521_3_LC_14_6_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_RNIC2521_3_LC_14_6_5 .LUT_INIT=16'b1010101011101110;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_RNIC2521_3_LC_14_6_5  (
            .in0(N__64599),
            .in1(N__63458),
            .in2(_gnd_net_),
            .in3(N__63545),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_RNIC2521Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_2_LC_14_6_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_2_LC_14_6_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_2_LC_14_6_6 .LUT_INIT=16'b0100001101000000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_2_LC_14_6_6  (
            .in0(N__58068),
            .in1(N__61632),
            .in2(N__61456),
            .in3(N__60904),
            .lcout(\ppm_encoder_1.pulses2count_9_i_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNI2JJC1_1_LC_14_6_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNI2JJC1_1_LC_14_6_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNI2JJC1_1_LC_14_6_7 .LUT_INIT=16'b0000110001011101;
    LogicCell40 \ppm_encoder_1.throttle_RNI2JJC1_1_LC_14_6_7  (
            .in0(N__58034),
            .in1(N__57963),
            .in2(N__57909),
            .in3(N__63544),
            .lcout(\ppm_encoder_1.throttle_RNI2JJC1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_21_c_RNO_LC_14_7_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_21_c_RNO_LC_14_7_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_21_c_RNO_LC_14_7_0 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_21_c_RNO_LC_14_7_0  (
            .in0(N__64850),
            .in1(N__57738),
            .in2(N__57804),
            .in3(N__64889),
            .lcout(\ppm_encoder_1.counter24_0_I_21_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_7_LC_14_7_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_7_LC_14_7_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_7_LC_14_7_1 .LUT_INIT=16'b1111111111011100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_7_LC_14_7_1  (
            .in0(N__57870),
            .in1(N__57843),
            .in2(N__63465),
            .in3(N__57831),
            .lcout(),
            .ltout(\ppm_encoder_1.pulses2count_9_i_2_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_7_LC_14_7_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_7_LC_14_7_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_7_LC_14_7_2 .LUT_INIT=16'b0000000000000011;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_7_LC_14_7_2  (
            .in0(_gnd_net_),
            .in1(N__57813),
            .in2(N__57807),
            .in3(N__61850),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87000),
            .ce(N__68744),
            .sr(N__79597));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_6_LC_14_7_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_6_LC_14_7_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_6_LC_14_7_3 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_6_LC_14_7_3  (
            .in0(N__63461),
            .in1(N__57795),
            .in2(N__61650),
            .in3(N__57762),
            .lcout(),
            .ltout(\ppm_encoder_1.pulses2count_9_0_2_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_6_LC_14_7_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_6_LC_14_7_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_6_LC_14_7_4 .LUT_INIT=16'b1111111111111100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_6_LC_14_7_4  (
            .in0(_gnd_net_),
            .in1(N__61701),
            .in2(N__57741),
            .in3(N__61849),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87000),
            .ce(N__68744),
            .sr(N__79597));
    defparam \ppm_encoder_1.pulses2count_esr_13_LC_14_7_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_13_LC_14_7_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_13_LC_14_7_7 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_13_LC_14_7_7  (
            .in0(N__61848),
            .in1(N__61281),
            .in2(_gnd_net_),
            .in3(N__57732),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87000),
            .ce(N__68744),
            .sr(N__79597));
    defparam \pid_side.un11lto30_i_a2_0_c_RNO_LC_14_8_1 .C_ON=1'b0;
    defparam \pid_side.un11lto30_i_a2_0_c_RNO_LC_14_8_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.un11lto30_i_a2_0_c_RNO_LC_14_8_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_side.un11lto30_i_a2_0_c_RNO_LC_14_8_1  (
            .in0(N__69116),
            .in1(N__69146),
            .in2(N__69089),
            .in3(N__69184),
            .lcout(\pid_side.source_pid10lt4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un11lto30_i_a2_1_c_RNO_LC_14_8_2 .C_ON=1'b0;
    defparam \pid_side.un11lto30_i_a2_1_c_RNO_LC_14_8_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.un11lto30_i_a2_1_c_RNO_LC_14_8_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_side.un11lto30_i_a2_1_c_RNO_LC_14_8_2  (
            .in0(N__69366),
            .in1(N__71732),
            .in2(N__71804),
            .in3(N__69411),
            .lcout(\pid_side.un11lto30_i_a2_0_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.source_pid_1_esr_6_LC_14_8_3 .C_ON=1'b0;
    defparam \pid_side.source_pid_1_esr_6_LC_14_8_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.source_pid_1_esr_6_LC_14_8_3 .LUT_INIT=16'b1010101010101111;
    LogicCell40 \pid_side.source_pid_1_esr_6_LC_14_8_3  (
            .in0(N__71733),
            .in1(_gnd_net_),
            .in2(N__58121),
            .in3(N__69990),
            .lcout(side_order_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87008),
            .ce(N__58293),
            .sr(N__58245));
    defparam \pid_side.source_pid_1_esr_2_LC_14_8_7 .C_ON=1'b0;
    defparam \pid_side.source_pid_1_esr_2_LC_14_8_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.source_pid_1_esr_2_LC_14_8_7 .LUT_INIT=16'b0010001000100000;
    LogicCell40 \pid_side.source_pid_1_esr_2_LC_14_8_7  (
            .in0(N__69117),
            .in1(N__58156),
            .in2(N__58122),
            .in3(N__69991),
            .lcout(side_order_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87008),
            .ce(N__58293),
            .sr(N__58245));
    defparam \pid_side.state_RNIH98N9_1_LC_14_9_0 .C_ON=1'b0;
    defparam \pid_side.state_RNIH98N9_1_LC_14_9_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.state_RNIH98N9_1_LC_14_9_0 .LUT_INIT=16'b1111101111110000;
    LogicCell40 \pid_side.state_RNIH98N9_1_LC_14_9_0  (
            .in0(N__61953),
            .in1(N__58128),
            .in2(N__66044),
            .in3(N__72618),
            .lcout(\pid_side.un1_reset_0_i ),
            .ltout(\pid_side.un1_reset_0_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.state_RNIA3KT9_1_LC_14_9_1 .C_ON=1'b0;
    defparam \pid_side.state_RNIA3KT9_1_LC_14_9_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.state_RNIA3KT9_1_LC_14_9_1 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \pid_side.state_RNIA3KT9_1_LC_14_9_1  (
            .in0(N__72619),
            .in1(_gnd_net_),
            .in2(N__58161),
            .in3(_gnd_net_),
            .lcout(\pid_side.state_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_esr_RNIRALN2_4_LC_14_9_3 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_esr_RNIRALN2_4_LC_14_9_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_esr_RNIRALN2_4_LC_14_9_3 .LUT_INIT=16'b0101010000000000;
    LogicCell40 \pid_side.pid_prereg_esr_RNIRALN2_4_LC_14_9_3  (
            .in0(N__69988),
            .in1(N__69374),
            .in2(N__69417),
            .in3(N__71590),
            .lcout(\pid_side.N_75 ),
            .ltout(\pid_side.N_75_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_esr_RNIDHBS3_30_LC_14_9_4 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_esr_RNIDHBS3_30_LC_14_9_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_esr_RNIDHBS3_30_LC_14_9_4 .LUT_INIT=16'b1111111111110001;
    LogicCell40 \pid_side.pid_prereg_esr_RNIDHBS3_30_LC_14_9_4  (
            .in0(N__61890),
            .in1(N__69989),
            .in2(N__58131),
            .in3(N__61959),
            .lcout(\pid_side.N_102 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_esr_RNIIATS_12_LC_14_9_6 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_esr_RNIIATS_12_LC_14_9_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_esr_RNIIATS_12_LC_14_9_6 .LUT_INIT=16'b0010001010101010;
    LogicCell40 \pid_side.pid_prereg_esr_RNIIATS_12_LC_14_9_6  (
            .in0(N__61891),
            .in1(N__71712),
            .in2(_gnd_net_),
            .in3(N__69501),
            .lcout(\pid_side.N_76 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.source_pid_1_esr_12_LC_14_10_0 .C_ON=1'b0;
    defparam \pid_side.source_pid_1_esr_12_LC_14_10_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.source_pid_1_esr_12_LC_14_10_0 .LUT_INIT=16'b1111001000000000;
    LogicCell40 \pid_side.source_pid_1_esr_12_LC_14_10_0  (
            .in0(N__61892),
            .in1(N__71710),
            .in2(N__70010),
            .in3(N__69498),
            .lcout(side_order_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87022),
            .ce(N__58291),
            .sr(N__58247));
    defparam \pid_side.source_pid_1_esr_13_LC_14_10_1 .C_ON=1'b0;
    defparam \pid_side.source_pid_1_esr_13_LC_14_10_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.source_pid_1_esr_13_LC_14_10_1 .LUT_INIT=16'b1010101010111011;
    LogicCell40 \pid_side.source_pid_1_esr_13_LC_14_10_1  (
            .in0(N__71709),
            .in1(N__70001),
            .in2(_gnd_net_),
            .in3(N__61893),
            .lcout(side_order_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87022),
            .ce(N__58291),
            .sr(N__58247));
    defparam \pid_side.un11lto30_i_a2_3_c_RNO_LC_14_10_2 .C_ON=1'b0;
    defparam \pid_side.un11lto30_i_a2_3_c_RNO_LC_14_10_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.un11lto30_i_a2_3_c_RNO_LC_14_10_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_side.un11lto30_i_a2_3_c_RNO_LC_14_10_2  (
            .in0(N__72692),
            .in1(N__71708),
            .in2(N__72723),
            .in3(N__69497),
            .lcout(\pid_side.un11lto30_i_a2_2_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_esr_RNIB2E2_28_LC_14_10_3 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_esr_RNIB2E2_28_LC_14_10_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_esr_RNIB2E2_28_LC_14_10_3 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \pid_side.pid_prereg_esr_RNIB2E2_28_LC_14_10_3  (
            .in0(N__70041),
            .in1(N__70000),
            .in2(_gnd_net_),
            .in3(N__69534),
            .lcout(\pid_side.un11lto30_i_a2_6_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.state_RNINK4U_0_LC_14_10_4 .C_ON=1'b0;
    defparam \pid_side.state_RNINK4U_0_LC_14_10_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.state_RNINK4U_0_LC_14_10_4 .LUT_INIT=16'b1111111100000010;
    LogicCell40 \pid_side.state_RNINK4U_0_LC_14_10_4  (
            .in0(N__59953),
            .in1(N__72613),
            .in2(N__59863),
            .in3(N__79922),
            .lcout(\pid_side.state_RNINK4UZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.state_RNIQ7UK_0_LC_14_10_6 .C_ON=1'b0;
    defparam \pid_side.state_RNIQ7UK_0_LC_14_10_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.state_RNIQ7UK_0_LC_14_10_6 .LUT_INIT=16'b0000000000001010;
    LogicCell40 \pid_side.state_RNIQ7UK_0_LC_14_10_6  (
            .in0(N__59954),
            .in1(_gnd_net_),
            .in2(N__59864),
            .in3(N__72614),
            .lcout(\pid_side.state_ns_0 ),
            .ltout(\pid_side.state_ns_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.state_RNINK4U_0_0_LC_14_10_7 .C_ON=1'b0;
    defparam \pid_side.state_RNINK4U_0_0_LC_14_10_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.state_RNINK4U_0_0_LC_14_10_7 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \pid_side.state_RNINK4U_0_0_LC_14_10_7  (
            .in0(N__79923),
            .in1(_gnd_net_),
            .in2(N__58206),
            .in3(_gnd_net_),
            .lcout(\pid_side.state_ns_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_7_LC_14_11_0 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_7_LC_14_11_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_7_LC_14_11_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_7_LC_14_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__66507),
            .lcout(\pid_side.error_i_acumm_preregZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87031),
            .ce(N__69892),
            .sr(N__79619));
    defparam \pid_side.error_i_acumm_prereg_esr_RNIJ04N_0_10_LC_14_11_1 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIJ04N_0_10_LC_14_11_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIJ04N_0_10_LC_14_11_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_RNIJ04N_0_10_LC_14_11_1  (
            .in0(_gnd_net_),
            .in1(N__65758),
            .in2(_gnd_net_),
            .in3(N__62005),
            .lcout(\pid_side.error_i_acumm_prereg_esr_RNIJ04N_0Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_RNIGSJV_7_LC_14_11_2 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIGSJV_7_LC_14_11_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIGSJV_7_LC_14_11_2 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_RNIGSJV_7_LC_14_11_2  (
            .in0(N__65804),
            .in1(N__62263),
            .in2(_gnd_net_),
            .in3(N__62281),
            .lcout(),
            .ltout(\pid_side.error_i_acumm_prereg_esr_RNIGSJVZ0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_RNIBT1C4_12_LC_14_11_3 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIBT1C4_12_LC_14_11_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIBT1C4_12_LC_14_11_3 .LUT_INIT=16'b0000010011001100;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_RNIBT1C4_12_LC_14_11_3  (
            .in0(N__61989),
            .in1(N__68365),
            .in2(N__58359),
            .in3(N__58356),
            .lcout(\pid_side.error_i_acumm_prereg_esr_RNIBT1C4Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_10_LC_14_11_4 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_10_LC_14_11_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_10_LC_14_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_10_LC_14_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__72933),
            .lcout(\pid_side.error_i_acumm_preregZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87031),
            .ce(N__69892),
            .sr(N__79619));
    defparam \pid_side.error_i_acumm_prereg_esr_RNIJ04N_10_LC_14_11_5 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIJ04N_10_LC_14_11_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIJ04N_10_LC_14_11_5 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_RNIJ04N_10_LC_14_11_5  (
            .in0(_gnd_net_),
            .in1(N__65759),
            .in2(_gnd_net_),
            .in3(N__62006),
            .lcout(\pid_side.error_i_acumm_prereg_esr_RNIJ04NZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_11_LC_14_11_6 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_11_LC_14_11_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_11_LC_14_11_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_11_LC_14_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78875),
            .lcout(\pid_side.error_i_acumm_preregZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87031),
            .ce(N__69892),
            .sr(N__79619));
    defparam \pid_side.error_i_acumm_prereg_esr_8_LC_14_11_7 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_8_LC_14_11_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_8_LC_14_11_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_8_LC_14_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__66468),
            .lcout(\pid_side.error_i_acumm_preregZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87031),
            .ce(N__69892),
            .sr(N__79619));
    defparam \pid_side.error_p_reg_esr_RNINKTC1_0_7_LC_14_12_0 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNINKTC1_0_7_LC_14_12_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNINKTC1_0_7_LC_14_12_0 .LUT_INIT=16'b0101101010010110;
    LogicCell40 \pid_side.error_p_reg_esr_RNINKTC1_0_7_LC_14_12_0  (
            .in0(N__58394),
            .in1(N__58379),
            .in2(N__84416),
            .in3(N__81268),
            .lcout(\pid_side.error_p_reg_esr_RNINKTC1_0Z0Z_7 ),
            .ltout(\pid_side.error_p_reg_esr_RNINKTC1_0Z0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNIODMH3_0_6_LC_14_12_1 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIODMH3_0_6_LC_14_12_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIODMH3_0_6_LC_14_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_p_reg_esr_RNIODMH3_0_6_LC_14_12_1  (
            .in0(_gnd_net_),
            .in1(N__58344),
            .in2(N__58350),
            .in3(N__66505),
            .lcout(\pid_side.error_p_reg_esr_RNIODMH3_0Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNISPEI_6_LC_14_12_2 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNISPEI_6_LC_14_12_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNISPEI_6_LC_14_12_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNISPEI_6_LC_14_12_2  (
            .in0(_gnd_net_),
            .in1(N__58378),
            .in2(_gnd_net_),
            .in3(N__81267),
            .lcout(\pid_side.N_2362_i ),
            .ltout(\pid_side.N_2362_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNIIFTC1_6_LC_14_12_3 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIIFTC1_6_LC_14_12_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIIFTC1_6_LC_14_12_3 .LUT_INIT=16'b1010111100101011;
    LogicCell40 \pid_side.error_p_reg_esr_RNIIFTC1_6_LC_14_12_3  (
            .in0(N__78591),
            .in1(N__78609),
            .in2(N__58347),
            .in3(N__81380),
            .lcout(\pid_side.error_p_reg_esr_RNIIFTC1Z0Z_6 ),
            .ltout(\pid_side.error_p_reg_esr_RNIIFTC1Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNIODMH3_6_LC_14_12_4 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIODMH3_6_LC_14_12_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIODMH3_6_LC_14_12_4 .LUT_INIT=16'b1111101010100000;
    LogicCell40 \pid_side.error_p_reg_esr_RNIODMH3_6_LC_14_12_4  (
            .in0(N__66506),
            .in1(_gnd_net_),
            .in2(N__58404),
            .in3(N__58401),
            .lcout(\pid_side.error_p_reg_esr_RNIODMH3Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_6_LC_14_12_5 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_6_LC_14_12_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_6_LC_14_12_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_6_LC_14_12_5  (
            .in0(N__81270),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_d_reg_prevZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87041),
            .ce(N__83399),
            .sr(N__83229));
    defparam \pid_side.error_p_reg_esr_RNINKTC1_7_LC_14_12_6 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNINKTC1_7_LC_14_12_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNINKTC1_7_LC_14_12_6 .LUT_INIT=16'b1111010101110001;
    LogicCell40 \pid_side.error_p_reg_esr_RNINKTC1_7_LC_14_12_6  (
            .in0(N__58395),
            .in1(N__58380),
            .in2(N__84417),
            .in3(N__81269),
            .lcout(\pid_side.error_p_reg_esr_RNINKTC1Z0Z_7 ),
            .ltout(\pid_side.error_p_reg_esr_RNINKTC1Z0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNIKF8V6_7_LC_14_12_7 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIKF8V6_7_LC_14_12_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIKF8V6_7_LC_14_12_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_p_reg_esr_RNIKF8V6_7_LC_14_12_7  (
            .in0(N__69311),
            .in1(N__62225),
            .in2(N__58368),
            .in3(N__66466),
            .lcout(\pid_side.error_p_reg_esr_RNIKF8V6Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_0_19_LC_14_13_0 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_0_19_LC_14_13_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_0_19_LC_14_13_0 .LUT_INIT=16'b1010100000001000;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_0_19_LC_14_13_0  (
            .in0(N__76656),
            .in1(N__74923),
            .in2(N__76942),
            .in3(N__58473),
            .lcout(),
            .ltout(\pid_side.error_i_reg_9_rn_0_19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_19_LC_14_13_1 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_19_LC_14_13_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_esr_19_LC_14_13_1 .LUT_INIT=16'b0011000011111100;
    LogicCell40 \pid_side.error_i_reg_esr_19_LC_14_13_1  (
            .in0(_gnd_net_),
            .in1(N__71286),
            .in2(N__58365),
            .in3(N__58515),
            .lcout(\pid_side.error_i_regZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87050),
            .ce(N__75289),
            .sr(N__79635));
    defparam \pid_side.error_i_reg_esr_RNO_0_14_LC_14_13_2 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_0_14_LC_14_13_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_0_14_LC_14_13_2 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_0_14_LC_14_13_2  (
            .in0(N__76241),
            .in1(N__71557),
            .in2(_gnd_net_),
            .in3(N__62318),
            .lcout(),
            .ltout(\pid_side.m2_2_03_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_14_LC_14_13_3 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_14_LC_14_13_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_esr_14_LC_14_13_3 .LUT_INIT=16'b1000000011000100;
    LogicCell40 \pid_side.error_i_reg_esr_14_LC_14_13_3  (
            .in0(N__76863),
            .in1(N__76658),
            .in2(N__58362),
            .in3(N__58410),
            .lcout(\pid_side.error_i_regZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87050),
            .ce(N__75289),
            .sr(N__79635));
    defparam \pid_side.error_i_reg_esr_RNO_0_27_LC_14_13_4 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_0_27_LC_14_13_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_0_27_LC_14_13_4 .LUT_INIT=16'b0000100010101000;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_0_27_LC_14_13_4  (
            .in0(N__76655),
            .in1(N__74921),
            .in2(N__76941),
            .in3(N__58533),
            .lcout(\pid_side.error_i_reg_9_rn_0_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_1_21_LC_14_13_5 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_1_21_LC_14_13_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_1_21_LC_14_13_5 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_1_21_LC_14_13_5  (
            .in0(N__74922),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__76853),
            .lcout(),
            .ltout(\pid_side.g3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_21_LC_14_13_6 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_21_LC_14_13_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_esr_21_LC_14_13_6 .LUT_INIT=16'b1010000010001000;
    LogicCell40 \pid_side.error_i_reg_esr_21_LC_14_13_6  (
            .in0(N__76657),
            .in1(N__58458),
            .in2(N__58452),
            .in3(N__59229),
            .lcout(\pid_side.error_i_regZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87050),
            .ce(N__75289),
            .sr(N__79635));
    defparam \pid_side.error_i_reg_esr_1_LC_14_13_7 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_1_LC_14_13_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_esr_1_LC_14_13_7 .LUT_INIT=16'b1000000011010000;
    LogicCell40 \pid_side.error_i_reg_esr_1_LC_14_13_7  (
            .in0(N__71558),
            .in1(N__70584),
            .in2(N__70979),
            .in3(N__67029),
            .lcout(\pid_side.error_i_regZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87050),
            .ce(N__75289),
            .sr(N__79635));
    defparam \pid_side.error_cry_3_0_c_RNI2JS52_LC_14_14_0 .C_ON=1'b0;
    defparam \pid_side.error_cry_3_0_c_RNI2JS52_LC_14_14_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_3_0_c_RNI2JS52_LC_14_14_0 .LUT_INIT=16'b0010010100101111;
    LogicCell40 \pid_side.error_cry_3_0_c_RNI2JS52_LC_14_14_0  (
            .in0(N__77903),
            .in1(N__75830),
            .in2(N__78423),
            .in3(N__74767),
            .lcout(),
            .ltout(\pid_side.m37_1_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_4_c_RNI8D2P3_LC_14_14_1 .C_ON=1'b0;
    defparam \pid_side.error_cry_4_c_RNI8D2P3_LC_14_14_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_4_c_RNI8D2P3_LC_14_14_1 .LUT_INIT=16'b1010000111110001;
    LogicCell40 \pid_side.error_cry_4_c_RNI8D2P3_LC_14_14_1  (
            .in0(N__80982),
            .in1(N__74655),
            .in2(N__58449),
            .in3(N__74591),
            .lcout(\pid_side.N_38_1 ),
            .ltout(\pid_side.N_38_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_2_22_LC_14_14_2 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_2_22_LC_14_14_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_2_22_LC_14_14_2 .LUT_INIT=16'b0000000100100011;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_2_22_LC_14_14_2  (
            .in0(N__80535),
            .in1(N__75697),
            .in2(N__58446),
            .in3(N__62552),
            .lcout(\pid_side.error_i_reg_esr_RNO_2Z0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_3_22_LC_14_14_3 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_3_22_LC_14_14_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_3_22_LC_14_14_3 .LUT_INIT=16'b1111010011110111;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_3_22_LC_14_14_3  (
            .in0(N__62553),
            .in1(N__80537),
            .in2(N__75741),
            .in3(N__62532),
            .lcout(),
            .ltout(\pid_side.error_i_reg_esr_RNO_3Z0Z_22_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_1_22_LC_14_14_4 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_1_22_LC_14_14_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_1_22_LC_14_14_4 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_1_22_LC_14_14_4  (
            .in0(N__62510),
            .in1(_gnd_net_),
            .in2(N__58443),
            .in3(N__58440),
            .lcout(\pid_side.error_i_reg_esr_RNO_1Z0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_2_14_LC_14_14_5 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_2_14_LC_14_14_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_2_14_LC_14_14_5 .LUT_INIT=16'b0100001101110011;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_2_14_LC_14_14_5  (
            .in0(N__62554),
            .in1(N__80536),
            .in2(N__80396),
            .in3(N__62533),
            .lcout(),
            .ltout(\pid_side.m136_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_1_14_LC_14_14_6 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_1_14_LC_14_14_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_1_14_LC_14_14_6 .LUT_INIT=16'b0000111001011110;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_1_14_LC_14_14_6  (
            .in0(N__75701),
            .in1(N__58424),
            .in2(N__58413),
            .in3(N__74929),
            .lcout(\pid_side.m18_2_03_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_1_0_c_RNIEAJ82_LC_14_15_0 .C_ON=1'b0;
    defparam \pid_side.error_cry_1_0_c_RNIEAJ82_LC_14_15_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_1_0_c_RNIEAJ82_LC_14_15_0 .LUT_INIT=16'b1011101010111111;
    LogicCell40 \pid_side.error_cry_1_0_c_RNIEAJ82_LC_14_15_0  (
            .in0(N__80974),
            .in1(N__75900),
            .in2(N__78419),
            .in3(N__75828),
            .lcout(\pid_side.error_cry_1_0_c_RNIEAJZ0Z82 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_1_0_c_RNIEAJ82_0_LC_14_15_1 .C_ON=1'b0;
    defparam \pid_side.error_cry_1_0_c_RNIEAJ82_0_LC_14_15_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_1_0_c_RNIEAJ82_0_LC_14_15_1 .LUT_INIT=16'b0000000000011101;
    LogicCell40 \pid_side.error_cry_1_0_c_RNIEAJ82_0_LC_14_15_1  (
            .in0(N__75829),
            .in1(N__78411),
            .in2(N__75908),
            .in3(N__80975),
            .lcout(),
            .ltout(\pid_side.error_cry_1_0_c_RNIEAJ82Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_1_0_c_RNIEKSB6_LC_14_15_2 .C_ON=1'b0;
    defparam \pid_side.error_cry_1_0_c_RNIEKSB6_LC_14_15_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_1_0_c_RNIEKSB6_LC_14_15_2 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \pid_side.error_cry_1_0_c_RNIEKSB6_LC_14_15_2  (
            .in0(_gnd_net_),
            .in1(N__58485),
            .in2(N__58479),
            .in3(N__70296),
            .lcout(\pid_side.N_39_0 ),
            .ltout(\pid_side.N_39_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_0_c_RNIPC708_LC_14_15_3 .C_ON=1'b0;
    defparam \pid_side.error_cry_0_c_RNIPC708_LC_14_15_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_0_c_RNIPC708_LC_14_15_3 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \pid_side.error_cry_0_c_RNIPC708_LC_14_15_3  (
            .in0(_gnd_net_),
            .in1(N__80515),
            .in2(N__58476),
            .in3(N__62350),
            .lcout(\pid_side.N_53_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_1_19_LC_14_15_4 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_1_19_LC_14_15_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_1_19_LC_14_15_4 .LUT_INIT=16'b0001000000010011;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_1_19_LC_14_15_4  (
            .in0(N__62351),
            .in1(N__80390),
            .in2(N__80567),
            .in3(N__62429),
            .lcout(\pid_side.m7_2_03 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_2_15_LC_14_15_5 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_2_15_LC_14_15_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_2_15_LC_14_15_5 .LUT_INIT=16'b0100001101110011;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_2_15_LC_14_15_5  (
            .in0(N__62430),
            .in1(N__80519),
            .in2(N__80397),
            .in3(N__62454),
            .lcout(),
            .ltout(\pid_side.m134_0_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_1_15_LC_14_15_6 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_1_15_LC_14_15_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_1_15_LC_14_15_6 .LUT_INIT=16'b0001111100011010;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_1_15_LC_14_15_6  (
            .in0(N__75749),
            .in1(N__74926),
            .in2(N__58464),
            .in3(N__62400),
            .lcout(),
            .ltout(\pid_side.m19_2_03_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_15_LC_14_15_7 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_15_LC_14_15_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_esr_15_LC_14_15_7 .LUT_INIT=16'b1000110000000100;
    LogicCell40 \pid_side.error_i_reg_esr_15_LC_14_15_7  (
            .in0(N__76943),
            .in1(N__76618),
            .in2(N__58461),
            .in3(N__62358),
            .lcout(\pid_side.error_i_regZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87068),
            .ce(N__75301),
            .sr(N__79651));
    defparam \pid_side.error_cry_5_c_RNIN1DB2_LC_14_16_0 .C_ON=1'b0;
    defparam \pid_side.error_cry_5_c_RNIN1DB2_LC_14_16_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_5_c_RNIN1DB2_LC_14_16_0 .LUT_INIT=16'b1010101111111011;
    LogicCell40 \pid_side.error_cry_5_c_RNIN1DB2_LC_14_16_0  (
            .in0(N__80962),
            .in1(N__74177),
            .in2(N__78416),
            .in3(N__74583),
            .lcout(),
            .ltout(\pid_side.error_cry_5_c_RNIN1DBZ0Z2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_5_c_RNIL5AI6_LC_14_16_1 .C_ON=1'b0;
    defparam \pid_side.error_cry_5_c_RNIL5AI6_LC_14_16_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_5_c_RNIL5AI6_LC_14_16_1 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \pid_side.error_cry_5_c_RNIL5AI6_LC_14_16_1  (
            .in0(_gnd_net_),
            .in1(N__70773),
            .in2(N__58545),
            .in3(N__58542),
            .lcout(\pid_side.N_49_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_5_c_RNIN1DB2_0_LC_14_16_2 .C_ON=1'b0;
    defparam \pid_side.error_cry_5_c_RNIN1DB2_0_LC_14_16_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_5_c_RNIN1DB2_0_LC_14_16_2 .LUT_INIT=16'b0000000101010001;
    LogicCell40 \pid_side.error_cry_5_c_RNIN1DB2_0_LC_14_16_2  (
            .in0(N__80961),
            .in1(N__74176),
            .in2(N__78415),
            .in3(N__74582),
            .lcout(\pid_side.error_cry_5_c_RNIN1DB2Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_0_7_LC_14_16_3 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_0_7_LC_14_16_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_0_7_LC_14_16_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_0_7_LC_14_16_3  (
            .in0(N__62431),
            .in1(N__80538),
            .in2(_gnd_net_),
            .in3(N__62456),
            .lcout(),
            .ltout(\pid_side.N_103_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_7_LC_14_16_4 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_7_LC_14_16_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_esr_7_LC_14_16_4 .LUT_INIT=16'b1000110000000100;
    LogicCell40 \pid_side.error_i_reg_esr_7_LC_14_16_4  (
            .in0(N__75702),
            .in1(N__75477),
            .in2(N__58536),
            .in3(N__62466),
            .lcout(\pid_side.error_i_regZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87079),
            .ce(N__75368),
            .sr(N__79659));
    defparam \pid_side.error_cry_7_c_RNI06B4E_LC_14_16_5 .C_ON=1'b0;
    defparam \pid_side.error_cry_7_c_RNI06B4E_LC_14_16_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_7_c_RNI06B4E_LC_14_16_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \pid_side.error_cry_7_c_RNI06B4E_LC_14_16_5  (
            .in0(N__62399),
            .in1(N__71460),
            .in2(_gnd_net_),
            .in3(N__62455),
            .lcout(\pid_side.N_50_1 ),
            .ltout(\pid_side.N_50_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_11_LC_14_16_6 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_11_LC_14_16_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_esr_11_LC_14_16_6 .LUT_INIT=16'b0100010000001100;
    LogicCell40 \pid_side.error_i_reg_esr_11_LC_14_16_6  (
            .in0(N__58532),
            .in1(N__75476),
            .in2(N__58518),
            .in3(N__75703),
            .lcout(\pid_side.error_i_regZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87079),
            .ce(N__75368),
            .sr(N__79659));
    defparam \pid_side.error_i_reg_esr_27_LC_14_16_7 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_27_LC_14_16_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_esr_27_LC_14_16_7 .LUT_INIT=16'b0111011100100010;
    LogicCell40 \pid_side.error_i_reg_esr_27_LC_14_16_7  (
            .in0(N__68290),
            .in1(N__58511),
            .in2(_gnd_net_),
            .in3(N__58500),
            .lcout(\pid_side.error_i_regZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87079),
            .ce(N__75368),
            .sr(N__79659));
    defparam \pid_front.state_0_LC_14_17_0 .C_ON=1'b0;
    defparam \pid_front.state_0_LC_14_17_0 .SEQ_MODE=4'b1000;
    defparam \pid_front.state_0_LC_14_17_0 .LUT_INIT=16'b0000000000001100;
    LogicCell40 \pid_front.state_0_LC_14_17_0  (
            .in0(_gnd_net_),
            .in1(N__59949),
            .in2(N__60184),
            .in3(N__60060),
            .lcout(\pid_front.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87093),
            .ce(),
            .sr(N__79666));
    defparam \pid_front.state_1_LC_14_17_1 .C_ON=1'b0;
    defparam \pid_front.state_1_LC_14_17_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.state_1_LC_14_17_1 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \pid_front.state_1_LC_14_17_1  (
            .in0(_gnd_net_),
            .in1(N__60165),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87093),
            .ce(),
            .sr(N__79666));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNIG6P4_4_LC_14_17_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNIG6P4_4_LC_14_17_4 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNIG6P4_4_LC_14_17_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_RNIG6P4_4_LC_14_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58491),
            .lcout(drone_H_disp_side_i_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNIH7P4_5_LC_14_17_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNIH7P4_5_LC_14_17_5 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNIH7P4_5_LC_14_17_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_RNIH7P4_5_LC_14_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58575),
            .lcout(drone_H_disp_side_i_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNII8P4_6_LC_14_17_6 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNII8P4_6_LC_14_17_6 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNII8P4_6_LC_14_17_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_RNII8P4_6_LC_14_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58569),
            .lcout(drone_H_disp_side_i_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNIJ9P4_7_LC_14_17_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNIJ9P4_7_LC_14_17_7 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNIJ9P4_7_LC_14_17_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_RNIJ9P4_7_LC_14_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58563),
            .lcout(drone_H_disp_side_i_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_3_21_LC_14_18_0 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_3_21_LC_14_18_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_3_21_LC_14_18_0 .LUT_INIT=16'b1100000111110001;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_3_21_LC_14_18_0  (
            .in0(N__74067),
            .in1(N__71970),
            .in2(N__62655),
            .in3(N__74502),
            .lcout(\pid_side.N_88_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_xy_ki_esr_1_LC_14_18_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_ki_esr_1_LC_14_18_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_ki_esr_1_LC_14_18_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_xy_ki_esr_1_LC_14_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84210),
            .lcout(xy_ki_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87109),
            .ce(N__78703),
            .sr(N__79673));
    defparam \pid_side.error_i_reg_esr_RNO_4_17_LC_14_18_2 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_4_17_LC_14_18_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_4_17_LC_14_18_2 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_4_17_LC_14_18_2  (
            .in0(N__71966),
            .in1(N__80725),
            .in2(N__80595),
            .in3(N__74403),
            .lcout(\pid_side.error_i_reg_esr_RNO_4Z0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_5_17_LC_14_18_3 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_5_17_LC_14_18_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_5_17_LC_14_18_3 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_5_17_LC_14_18_3  (
            .in0(N__74402),
            .in1(N__80554),
            .in2(N__80766),
            .in3(N__71967),
            .lcout(\pid_side.error_i_reg_esr_RNO_5Z0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_xy_ki_esr_0_LC_14_18_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_ki_esr_0_LC_14_18_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_ki_esr_0_LC_14_18_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_xy_ki_esr_0_LC_14_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__83828),
            .lcout(xy_ki_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87109),
            .ce(N__78703),
            .sr(N__79673));
    defparam \Commands_frame_decoder.source_xy_ki_2_rep2_esr_LC_14_18_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_ki_2_rep2_esr_LC_14_18_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_ki_2_rep2_esr_LC_14_18_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_xy_ki_2_rep2_esr_LC_14_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__77574),
            .lcout(xy_ki_2_rep2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87109),
            .ce(N__78703),
            .sr(N__79673));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_1_LC_14_19_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_1_LC_14_19_0 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_1_LC_14_19_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_1_LC_14_19_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59196),
            .lcout(drone_H_disp_front_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87123),
            .ce(N__59246),
            .sr(N__79679));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_2_LC_14_19_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_2_LC_14_19_1 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_2_LC_14_19_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_2_LC_14_19_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59104),
            .lcout(drone_H_disp_front_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87123),
            .ce(N__59246),
            .sr(N__79679));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_3_LC_14_19_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_3_LC_14_19_2 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_3_LC_14_19_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_3_LC_14_19_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59023),
            .lcout(drone_H_disp_front_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87123),
            .ce(N__59246),
            .sr(N__79679));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_4_LC_14_19_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_4_LC_14_19_3 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_4_LC_14_19_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_4_LC_14_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58929),
            .lcout(\dron_frame_decoder_1.drone_H_disp_front_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87123),
            .ce(N__59246),
            .sr(N__79679));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_5_LC_14_19_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_5_LC_14_19_4 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_5_LC_14_19_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_5_LC_14_19_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58833),
            .lcout(\dron_frame_decoder_1.drone_H_disp_front_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87123),
            .ce(N__59246),
            .sr(N__79679));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_6_LC_14_19_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_6_LC_14_19_5 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_6_LC_14_19_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_6_LC_14_19_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58753),
            .lcout(\dron_frame_decoder_1.drone_H_disp_front_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87123),
            .ce(N__59246),
            .sr(N__79679));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_7_LC_14_19_6 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_7_LC_14_19_6 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_7_LC_14_19_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_7_LC_14_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58644),
            .lcout(\dron_frame_decoder_1.drone_H_disp_front_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87123),
            .ce(N__59246),
            .sr(N__79679));
    defparam \pid_front.m12_1_LC_14_20_1 .C_ON=1'b0;
    defparam \pid_front.m12_1_LC_14_20_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.m12_1_LC_14_20_1 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \pid_front.m12_1_LC_14_20_1  (
            .in0(N__78399),
            .in1(N__78091),
            .in2(_gnd_net_),
            .in3(N__77232),
            .lcout(\pid_front.m0_0_03 ),
            .ltout(\pid_front.m0_0_03_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_3_16_LC_14_20_2 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_3_16_LC_14_20_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_3_16_LC_14_20_2 .LUT_INIT=16'b0011000000010001;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_3_16_LC_14_20_2  (
            .in0(N__63150),
            .in1(N__80347),
            .in2(N__58578),
            .in3(N__77759),
            .lcout(\pid_front.m4_2_03 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_0_LC_14_20_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_0_LC_14_20_3 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_0_LC_14_20_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_0_LC_14_20_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59302),
            .lcout(drone_H_disp_front_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87138),
            .ce(N__59250),
            .sr(N__79681));
    defparam \dron_frame_decoder_1.source_H_disp_front_fast_esr_0_LC_14_20_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_fast_esr_0_LC_14_20_4 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_fast_esr_0_LC_14_20_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_fast_esr_0_LC_14_20_4  (
            .in0(N__59303),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(dron_frame_decoder_1_source_H_disp_front_fast_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87138),
            .ce(N__59250),
            .sr(N__79681));
    defparam \pid_front.m61_0_bm_LC_14_20_5 .C_ON=1'b0;
    defparam \pid_front.m61_0_bm_LC_14_20_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.m61_0_bm_LC_14_20_5 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \pid_front.m61_0_bm_LC_14_20_5  (
            .in0(N__72008),
            .in1(N__80764),
            .in2(N__77782),
            .in3(N__77233),
            .lcout(\pid_front.m61_0_bm_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_2_21_LC_14_20_7 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_2_21_LC_14_20_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_2_21_LC_14_20_7 .LUT_INIT=16'b0010001111100011;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_2_21_LC_14_20_7  (
            .in0(N__74676),
            .in1(N__76300),
            .in2(N__77030),
            .in3(N__62748),
            .lcout(\pid_side.un4_error_i_reg_31_ns_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_0_0_c_RNILPEB2_LC_14_21_0 .C_ON=1'b0;
    defparam \pid_front.error_cry_0_0_c_RNILPEB2_LC_14_21_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_0_0_c_RNILPEB2_LC_14_21_0 .LUT_INIT=16'b1010000110101011;
    LogicCell40 \pid_front.error_cry_0_0_c_RNILPEB2_LC_14_21_0  (
            .in0(N__59214),
            .in1(N__67838),
            .in2(N__77897),
            .in3(N__67784),
            .lcout(\pid_front.N_12_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_3_0_c_RNIJ5832_0_LC_14_21_1 .C_ON=1'b0;
    defparam \pid_front.error_cry_3_0_c_RNIJ5832_0_LC_14_21_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_3_0_c_RNIJ5832_0_LC_14_21_1 .LUT_INIT=16'b0000010000000111;
    LogicCell40 \pid_front.error_cry_3_0_c_RNIJ5832_0_LC_14_21_1  (
            .in0(N__67638),
            .in1(N__78218),
            .in2(N__78103),
            .in3(N__62969),
            .lcout(\pid_front.error_cry_3_0_c_RNIJ5832Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_1_c_RNI1AE71_LC_14_21_2 .C_ON=1'b0;
    defparam \pid_front.error_cry_1_c_RNI1AE71_LC_14_21_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_1_c_RNI1AE71_LC_14_21_2 .LUT_INIT=16'b0010010101110101;
    LogicCell40 \pid_front.error_cry_1_c_RNI1AE71_LC_14_21_2  (
            .in0(N__78217),
            .in1(N__77118),
            .in2(N__77896),
            .in3(N__77060),
            .lcout(\pid_front.m11_0_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_4_c_RNI7DKG1_LC_14_21_3 .C_ON=1'b0;
    defparam \pid_front.error_cry_4_c_RNI7DKG1_LC_14_21_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_4_c_RNI7DKG1_LC_14_21_3 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \pid_front.error_cry_4_c_RNI7DKG1_LC_14_21_3  (
            .in0(N__78220),
            .in1(N__62968),
            .in2(_gnd_net_),
            .in3(N__59436),
            .lcout(\pid_front.N_48_1 ),
            .ltout(\pid_front.N_48_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_1_0_c_RNIOOIF3_0_LC_14_21_4 .C_ON=1'b0;
    defparam \pid_front.error_cry_1_0_c_RNIOOIF3_0_LC_14_21_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_1_0_c_RNIOOIF3_0_LC_14_21_4 .LUT_INIT=16'b0010001000110000;
    LogicCell40 \pid_front.error_cry_1_0_c_RNIOOIF3_0_LC_14_21_4  (
            .in0(N__72263),
            .in1(N__77755),
            .in2(N__59208),
            .in3(N__78090),
            .lcout(),
            .ltout(\pid_front.error_cry_1_0_c_RNIOOIF3Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_0_0_c_RNI5BKA9_LC_14_21_5 .C_ON=1'b0;
    defparam \pid_front.error_cry_0_0_c_RNI5BKA9_LC_14_21_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_0_0_c_RNI5BKA9_LC_14_21_5 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \pid_front.error_cry_0_0_c_RNI5BKA9_LC_14_21_5  (
            .in0(_gnd_net_),
            .in1(N__70857),
            .in2(N__59391),
            .in3(N__59385),
            .lcout(\pid_front.N_116_0 ),
            .ltout(\pid_front.N_116_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_0_c_RNIKMQ0B_LC_14_21_6 .C_ON=1'b0;
    defparam \pid_front.error_cry_0_c_RNIKMQ0B_LC_14_21_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_0_c_RNIKMQ0B_LC_14_21_6 .LUT_INIT=16'b0010011100000101;
    LogicCell40 \pid_front.error_cry_0_c_RNIKMQ0B_LC_14_21_6  (
            .in0(N__76301),
            .in1(N__71501),
            .in2(N__59388),
            .in3(N__71022),
            .lcout(\pid_front.m9_2_03_3_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_1_0_c_RNIOOIF3_LC_14_21_7 .C_ON=1'b0;
    defparam \pid_front.error_cry_1_0_c_RNIOOIF3_LC_14_21_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_1_0_c_RNIOOIF3_LC_14_21_7 .LUT_INIT=16'b1111110111111000;
    LogicCell40 \pid_front.error_cry_1_0_c_RNIOOIF3_LC_14_21_7  (
            .in0(N__78089),
            .in1(N__72262),
            .in2(N__77781),
            .in3(N__72223),
            .lcout(\pid_front.error_cry_1_0_c_RNIOOIFZ0Z3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_4_c_RNI5OS71_LC_14_22_0 .C_ON=1'b0;
    defparam \pid_front.error_cry_4_c_RNI5OS71_LC_14_22_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_4_c_RNI5OS71_LC_14_22_0 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \pid_front.error_cry_4_c_RNI5OS71_LC_14_22_0  (
            .in0(N__78249),
            .in1(N__59435),
            .in2(_gnd_net_),
            .in3(N__67313),
            .lcout(\pid_front.N_21_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_6_c_RNI1ADU1_LC_14_22_1 .C_ON=1'b0;
    defparam \pid_front.error_cry_6_c_RNI1ADU1_LC_14_22_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_6_c_RNI1ADU1_LC_14_22_1 .LUT_INIT=16'b1111001011110111;
    LogicCell40 \pid_front.error_cry_6_c_RNI1ADU1_LC_14_22_1  (
            .in0(N__78250),
            .in1(N__67380),
            .in2(N__78092),
            .in3(N__67165),
            .lcout(\pid_front.error_cry_6_c_RNI1ADUZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_6_c_RNI1ADU1_0_LC_14_22_2 .C_ON=1'b0;
    defparam \pid_front.error_cry_6_c_RNI1ADU1_0_LC_14_22_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_6_c_RNI1ADU1_0_LC_14_22_2 .LUT_INIT=16'b0000001100010001;
    LogicCell40 \pid_front.error_cry_6_c_RNI1ADU1_0_LC_14_22_2  (
            .in0(N__67166),
            .in1(N__78061),
            .in2(N__67397),
            .in3(N__78251),
            .lcout(),
            .ltout(\pid_front.error_cry_6_c_RNI1ADU1Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_4_c_RNI7CN45_LC_14_22_3 .C_ON=1'b0;
    defparam \pid_front.error_cry_4_c_RNI7CN45_LC_14_22_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_4_c_RNI7CN45_LC_14_22_3 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \pid_front.error_cry_4_c_RNI7CN45_LC_14_22_3  (
            .in0(_gnd_net_),
            .in1(N__59379),
            .in2(N__59373),
            .in3(N__59370),
            .lcout(\pid_front.N_22_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_1_16_LC_14_22_4 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_1_16_LC_14_22_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_1_16_LC_14_22_4 .LUT_INIT=16'b1010001000000010;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_1_16_LC_14_22_4  (
            .in0(N__76611),
            .in1(N__59397),
            .in2(N__77029),
            .in3(N__59364),
            .lcout(),
            .ltout(\pid_front.error_i_reg_9_rn_0_16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_16_LC_14_22_5 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_16_LC_14_22_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_esr_16_LC_14_22_5 .LUT_INIT=16'b0101000011111010;
    LogicCell40 \pid_front.error_i_reg_esr_16_LC_14_22_5  (
            .in0(N__71271),
            .in1(_gnd_net_),
            .in2(N__59355),
            .in3(N__59340),
            .lcout(\pid_front.error_i_regZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87170),
            .ce(N__72353),
            .sr(N__79689));
    defparam \pid_front.error_i_reg_esr_RNO_0_16_LC_14_22_6 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_0_16_LC_14_22_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_0_16_LC_14_22_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_0_16_LC_14_22_6  (
            .in0(N__71556),
            .in1(N__62901),
            .in2(_gnd_net_),
            .in3(N__63101),
            .lcout(\pid_front.error_i_reg_esr_RNO_0Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_8_c_RNIQ06A1_LC_14_23_0 .C_ON=1'b0;
    defparam \pid_front.error_cry_8_c_RNIQ06A1_LC_14_23_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_8_c_RNIQ06A1_LC_14_23_0 .LUT_INIT=16'b0101000001011111;
    LogicCell40 \pid_front.error_cry_8_c_RNIQ06A1_LC_14_23_0  (
            .in0(N__67215),
            .in1(_gnd_net_),
            .in2(N__78417),
            .in3(N__72093),
            .lcout(\pid_front.N_36_0 ),
            .ltout(\pid_front.N_36_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_6_c_RNITTOU2_LC_14_23_1 .C_ON=1'b0;
    defparam \pid_front.error_cry_6_c_RNITTOU2_LC_14_23_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_6_c_RNITTOU2_LC_14_23_1 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \pid_front.error_cry_6_c_RNITTOU2_LC_14_23_1  (
            .in0(N__72038),
            .in1(_gnd_net_),
            .in2(N__59409),
            .in3(N__59403),
            .lcout(\pid_front.N_37_1 ),
            .ltout(\pid_front.N_37_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_0_14_LC_14_23_2 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_0_14_LC_14_23_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_0_14_LC_14_23_2 .LUT_INIT=16'b1111000001010101;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_0_14_LC_14_23_2  (
            .in0(N__71123),
            .in1(_gnd_net_),
            .in2(N__59406),
            .in3(N__71544),
            .lcout(\pid_front.N_136 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_6_c_RNIU0FF1_LC_14_23_3 .C_ON=1'b0;
    defparam \pid_front.error_cry_6_c_RNIU0FF1_LC_14_23_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_6_c_RNIU0FF1_LC_14_23_3 .LUT_INIT=16'b0100010001110111;
    LogicCell40 \pid_front.error_cry_6_c_RNIU0FF1_LC_14_23_3  (
            .in0(N__67390),
            .in1(N__78246),
            .in2(_gnd_net_),
            .in3(N__67164),
            .lcout(\pid_front.N_18_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_1_22_LC_14_23_4 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_1_22_LC_14_23_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_1_22_LC_14_23_4 .LUT_INIT=16'b1100010101010101;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_1_22_LC_14_23_4  (
            .in0(N__71124),
            .in1(N__59618),
            .in2(N__76319),
            .in3(N__71545),
            .lcout(\pid_front.m26_2_03_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_2_16_LC_14_23_5 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_2_16_LC_14_23_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_2_16_LC_14_23_5 .LUT_INIT=16'b1000000011011111;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_2_16_LC_14_23_5  (
            .in0(N__72039),
            .in1(N__62859),
            .in2(N__77794),
            .in3(N__71122),
            .lcout(\pid_front.error_i_reg_esr_RNO_2_0_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_4_c_RNI81RM1_0_LC_14_23_6 .C_ON=1'b0;
    defparam \pid_front.error_cry_4_c_RNI81RM1_0_LC_14_23_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_4_c_RNI81RM1_0_LC_14_23_6 .LUT_INIT=16'b0000001000000111;
    LogicCell40 \pid_front.error_cry_4_c_RNI81RM1_0_LC_14_23_6  (
            .in0(N__78245),
            .in1(N__59437),
            .in2(N__78099),
            .in3(N__67305),
            .lcout(\pid_front.error_cry_4_c_RNI81RM1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_8_c_RNIO00A1_LC_14_23_7 .C_ON=1'b0;
    defparam \pid_front.error_cry_8_c_RNIO00A1_LC_14_23_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_8_c_RNIO00A1_LC_14_23_7 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \pid_front.error_cry_8_c_RNIO00A1_LC_14_23_7  (
            .in0(N__80778),
            .in1(N__67214),
            .in2(_gnd_net_),
            .in3(N__67163),
            .lcout(\pid_front.N_45_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_4_21_LC_14_24_0 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_4_21_LC_14_24_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_4_21_LC_14_24_0 .LUT_INIT=16'b0010010101110101;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_4_21_LC_14_24_0  (
            .in0(N__78252),
            .in1(N__67307),
            .in2(N__77904),
            .in3(N__67391),
            .lcout(),
            .ltout(\pid_front.error_i_reg_esr_RNO_4Z0Z_21_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_1_21_LC_14_24_1 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_1_21_LC_14_24_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_1_21_LC_14_24_1 .LUT_INIT=16'b1011000010110101;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_1_21_LC_14_24_1  (
            .in0(N__77902),
            .in1(N__67233),
            .in2(N__59535),
            .in3(N__67179),
            .lcout(\pid_front.N_88_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_3_21_LC_14_24_2 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_3_21_LC_14_24_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_3_21_LC_14_24_2 .LUT_INIT=16'b0100010001110111;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_3_21_LC_14_24_2  (
            .in0(N__77405),
            .in1(N__80377),
            .in2(_gnd_net_),
            .in3(N__71169),
            .lcout(\pid_front.g0_5_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_2_21_LC_14_24_3 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_2_21_LC_14_24_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_2_21_LC_14_24_3 .LUT_INIT=16'b0001010111010101;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_2_21_LC_14_24_3  (
            .in0(N__71170),
            .in1(N__77901),
            .in2(N__78407),
            .in3(N__72120),
            .lcout(),
            .ltout(\pid_front.N_126_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_0_21_LC_14_24_4 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_0_21_LC_14_24_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_0_21_LC_14_24_4 .LUT_INIT=16'b1110011011000100;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_0_21_LC_14_24_4  (
            .in0(N__80382),
            .in1(N__59532),
            .in2(N__59526),
            .in3(N__59523),
            .lcout(),
            .ltout(\pid_front.m25_2_03_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_21_LC_14_24_5 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_21_LC_14_24_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_esr_21_LC_14_24_5 .LUT_INIT=16'b1000101000000010;
    LogicCell40 \pid_front.error_i_reg_esr_21_LC_14_24_5  (
            .in0(N__76640),
            .in1(N__76954),
            .in2(N__59517),
            .in3(N__59514),
            .lcout(\pid_front.error_i_regZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87199),
            .ce(N__72412),
            .sr(N__79695));
    defparam \pid_front.error_i_reg_esr_12_LC_14_24_6 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_12_LC_14_24_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_esr_12_LC_14_24_6 .LUT_INIT=16'b1000110100000000;
    LogicCell40 \pid_front.error_i_reg_esr_12_LC_14_24_6  (
            .in0(N__76953),
            .in1(N__63057),
            .in2(N__63009),
            .in3(N__76641),
            .lcout(\pid_front.error_i_regZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87199),
            .ce(N__72412),
            .sr(N__79695));
    defparam \pid_front.error_cry_3_0_c_RNIGS9K1_LC_14_25_0 .C_ON=1'b0;
    defparam \pid_front.error_cry_3_0_c_RNIGS9K1_LC_14_25_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_3_0_c_RNIGS9K1_LC_14_25_0 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \pid_front.error_cry_3_0_c_RNIGS9K1_LC_14_25_0  (
            .in0(N__78247),
            .in1(N__67663),
            .in2(_gnd_net_),
            .in3(N__62986),
            .lcout(\pid_front.N_25_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_18_LC_14_25_1 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_18_LC_14_25_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_esr_18_LC_14_25_1 .LUT_INIT=16'b0111011100100010;
    LogicCell40 \pid_front.error_i_reg_esr_18_LC_14_25_1  (
            .in0(N__71281),
            .in1(N__63023),
            .in2(_gnd_net_),
            .in3(N__62841),
            .lcout(\pid_front.error_i_regZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87218),
            .ce(N__72407),
            .sr(N__79702));
    defparam \pid_front.error_cry_4_c_RNI81RM1_LC_14_25_4 .C_ON=1'b0;
    defparam \pid_front.error_cry_4_c_RNI81RM1_LC_14_25_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_4_c_RNI81RM1_LC_14_25_4 .LUT_INIT=16'b1111001011110111;
    LogicCell40 \pid_front.error_cry_4_c_RNI81RM1_LC_14_25_4  (
            .in0(N__78248),
            .in1(N__59455),
            .in2(N__78105),
            .in3(N__67306),
            .lcout(),
            .ltout(\pid_front.error_cry_4_c_RNI81RMZ0Z1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_4_c_RNI0VV15_LC_14_25_5 .C_ON=1'b0;
    defparam \pid_front.error_cry_4_c_RNI0VV15_LC_14_25_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_4_c_RNI0VV15_LC_14_25_5 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \pid_front.error_cry_4_c_RNI0VV15_LC_14_25_5  (
            .in0(_gnd_net_),
            .in1(N__59640),
            .in2(N__59634),
            .in3(N__59631),
            .lcout(\pid_front.N_38_1 ),
            .ltout(\pid_front.N_38_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_4_c_RNI2J198_LC_14_25_6 .C_ON=1'b0;
    defparam \pid_front.error_cry_4_c_RNI2J198_LC_14_25_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_4_c_RNI2J198_LC_14_25_6 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \pid_front.error_cry_4_c_RNI2J198_LC_14_25_6  (
            .in0(_gnd_net_),
            .in1(N__80568),
            .in2(N__59622),
            .in3(N__59619),
            .lcout(\pid_front.N_39_1 ),
            .ltout(\pid_front.N_39_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_10_LC_14_25_7 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_10_LC_14_25_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_esr_10_LC_14_25_7 .LUT_INIT=16'b1000101000000010;
    LogicCell40 \pid_front.error_i_reg_esr_10_LC_14_25_7  (
            .in0(N__75532),
            .in1(N__75753),
            .in2(N__59604),
            .in3(N__62766),
            .lcout(\pid_front.error_i_regZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87218),
            .ce(N__72407),
            .sr(N__79702));
    defparam \pid_front.error_i_reg_esr_RNO_2_14_LC_14_26_0 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_2_14_LC_14_26_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_2_14_LC_14_26_0 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_2_14_LC_14_26_0  (
            .in0(N__77767),
            .in1(N__67587),
            .in2(_gnd_net_),
            .in3(N__62827),
            .lcout(\pid_front.m2_2_03 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_4_c_RNIMVJS7_LC_14_26_1 .C_ON=1'b0;
    defparam \pid_front.error_cry_4_c_RNIMVJS7_LC_14_26_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_4_c_RNIMVJS7_LC_14_26_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \pid_front.error_cry_4_c_RNIMVJS7_LC_14_26_1  (
            .in0(N__77783),
            .in1(N__62790),
            .in2(_gnd_net_),
            .in3(N__59592),
            .lcout(\pid_front.N_110 ),
            .ltout(\pid_front.N_110_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_1_14_LC_14_26_2 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_1_14_LC_14_26_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_1_14_LC_14_26_2 .LUT_INIT=16'b1000110000000100;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_1_14_LC_14_26_2  (
            .in0(N__77012),
            .in1(N__76637),
            .in2(N__59586),
            .in3(N__59583),
            .lcout(),
            .ltout(\pid_front.error_i_reg_9_rn_1_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_14_LC_14_26_3 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_14_LC_14_26_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_esr_14_LC_14_26_3 .LUT_INIT=16'b0011000011111100;
    LogicCell40 \pid_front.error_i_reg_esr_14_LC_14_26_3  (
            .in0(_gnd_net_),
            .in1(N__70978),
            .in2(N__59577),
            .in3(N__59574),
            .lcout(\pid_front.error_i_regZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87231),
            .ce(N__72408),
            .sr(N__79706));
    defparam \pid_front.error_i_reg_esr_RNO_0_22_LC_14_26_5 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_0_22_LC_14_26_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_0_22_LC_14_26_5 .LUT_INIT=16'b0010000000101111;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_0_22_LC_14_26_5  (
            .in0(N__62828),
            .in1(N__77411),
            .in2(N__76326),
            .in3(N__67928),
            .lcout(),
            .ltout(\pid_front.m10_2_03_3_i_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_22_LC_14_26_6 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_22_LC_14_26_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_esr_22_LC_14_26_6 .LUT_INIT=16'b1000000011000100;
    LogicCell40 \pid_front.error_i_reg_esr_22_LC_14_26_6  (
            .in0(N__77013),
            .in1(N__76638),
            .in2(N__59556),
            .in3(N__59553),
            .lcout(\pid_front.error_i_regZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87231),
            .ce(N__72408),
            .sr(N__79706));
    defparam \pid_front.state_RNIQUOP1_0_LC_14_28_0 .C_ON=1'b0;
    defparam \pid_front.state_RNIQUOP1_0_LC_14_28_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.state_RNIQUOP1_0_LC_14_28_0 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \pid_front.state_RNIQUOP1_0_LC_14_28_0  (
            .in0(N__59952),
            .in1(N__70602),
            .in2(N__59973),
            .in3(N__60203),
            .lcout(),
            .ltout(\pid_front.N_196_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.state_RNIGSDC2_0_LC_14_28_1 .C_ON=1'b0;
    defparam \pid_front.state_RNIGSDC2_0_LC_14_28_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.state_RNIGSDC2_0_LC_14_28_1 .LUT_INIT=16'b1111111101110100;
    LogicCell40 \pid_front.state_RNIGSDC2_0_LC_14_28_1  (
            .in0(N__60204),
            .in1(N__60114),
            .in2(N__60009),
            .in3(N__79933),
            .lcout(\pid_front.error_i_acumm_1_sqmuxa_1_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.m153_e_5_LC_14_28_3 .C_ON=1'b0;
    defparam \pid_side.m153_e_5_LC_14_28_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.m153_e_5_LC_14_28_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \pid_side.m153_e_5_LC_14_28_3  (
            .in0(N__67586),
            .in1(N__80981),
            .in2(N__77002),
            .in3(N__80793),
            .lcout(pid_side_m153_e_5),
            .ltout(pid_side_m153_e_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.state_RNIMFDR1_0_LC_14_28_4 .C_ON=1'b0;
    defparam \pid_side.state_RNIMFDR1_0_LC_14_28_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.state_RNIMFDR1_0_LC_14_28_4 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \pid_side.state_RNIMFDR1_0_LC_14_28_4  (
            .in0(N__59951),
            .in1(N__70601),
            .in2(N__59874),
            .in3(N__59871),
            .lcout(\pid_side.N_196_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_15_c_RNO_LC_15_2_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_15_c_RNO_LC_15_2_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_15_c_RNO_LC_15_2_0 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_15_c_RNO_LC_15_2_0  (
            .in0(N__59679),
            .in1(N__64916),
            .in2(N__60423),
            .in3(N__64946),
            .lcout(\ppm_encoder_1.counter24_0_I_15_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_4_LC_15_2_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_4_LC_15_2_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_4_LC_15_2_1 .LUT_INIT=16'b1111110011111110;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_4_LC_15_2_1  (
            .in0(N__63422),
            .in1(N__61852),
            .in2(N__59775),
            .in3(N__59757),
            .lcout(),
            .ltout(\ppm_encoder_1.pulses2count_9_i_2_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_4_LC_15_2_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_4_LC_15_2_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_4_LC_15_2_2 .LUT_INIT=16'b0000010100000001;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_4_LC_15_2_2  (
            .in0(N__59736),
            .in1(N__64391),
            .in2(N__59721),
            .in3(N__59717),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__86975),
            .ce(N__68758),
            .sr(N__79572));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_5_LC_15_2_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_5_LC_15_2_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_5_LC_15_2_3 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_5_LC_15_2_3  (
            .in0(N__64390),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59673),
            .lcout(),
            .ltout(\ppm_encoder_1.pulses2count_esr_RNO_2Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_5_LC_15_2_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_5_LC_15_2_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_5_LC_15_2_4 .LUT_INIT=16'b1111101011111110;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_5_LC_15_2_4  (
            .in0(N__60474),
            .in1(N__63423),
            .in2(N__60462),
            .in3(N__60459),
            .lcout(),
            .ltout(\ppm_encoder_1.pulses2count_9_i_2_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_5_LC_15_2_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_5_LC_15_2_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_5_LC_15_2_5 .LUT_INIT=16'b0000000000000011;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_5_LC_15_2_5  (
            .in0(_gnd_net_),
            .in1(N__60438),
            .in2(N__60426),
            .in3(N__61854),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__86975),
            .ce(N__68758),
            .sr(N__79572));
    defparam \ppm_encoder_1.pulses2count_esr_0_LC_15_2_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_0_LC_15_2_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_0_LC_15_2_6 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_0_LC_15_2_6  (
            .in0(N__61853),
            .in1(N__60414),
            .in2(_gnd_net_),
            .in3(N__63510),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__86975),
            .ce(N__68758),
            .sr(N__79572));
    defparam \ppm_encoder_1.counter24_0_I_39_c_RNO_LC_15_3_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_39_c_RNO_LC_15_3_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_39_c_RNO_LC_15_3_0 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_39_c_RNO_LC_15_3_0  (
            .in0(N__60327),
            .in1(N__65553),
            .in2(N__60399),
            .in3(N__65577),
            .lcout(\ppm_encoder_1.counter24_0_I_39_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_12_LC_15_3_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_12_LC_15_3_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_12_LC_15_3_1 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_12_LC_15_3_1  (
            .in0(N__60375),
            .in1(N__68902),
            .in2(N__68820),
            .in3(N__60345),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__86981),
            .ce(N__68766),
            .sr(N__79579));
    defparam \ppm_encoder_1.pulses2count_esr_11_LC_15_3_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_11_LC_15_3_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_11_LC_15_3_2 .LUT_INIT=16'b1111111111101100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_11_LC_15_3_2  (
            .in0(N__68901),
            .in1(N__60321),
            .in2(N__60306),
            .in3(N__68819),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__86981),
            .ce(N__68766),
            .sr(N__79579));
    defparam \ppm_encoder_1.counter24_0_I_9_c_RNO_LC_15_3_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_9_c_RNO_LC_15_3_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_9_c_RNO_LC_15_3_4 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_9_c_RNO_LC_15_3_4  (
            .in0(N__68455),
            .in1(N__68778),
            .in2(N__68139),
            .in3(N__68410),
            .lcout(\ppm_encoder_1.counter24_0_I_9_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_27_c_RNO_LC_15_4_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_27_c_RNO_LC_15_4_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_27_c_RNO_LC_15_4_0 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_27_c_RNO_LC_15_4_0  (
            .in0(N__60210),
            .in1(N__64801),
            .in2(N__60618),
            .in3(N__64822),
            .lcout(\ppm_encoder_1.counter24_0_I_27_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_8_LC_15_4_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_8_LC_15_4_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_8_LC_15_4_1 .LUT_INIT=16'b0000001100000001;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_8_LC_15_4_1  (
            .in0(N__64436),
            .in1(N__60648),
            .in2(N__60261),
            .in3(N__60243),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__86987),
            .ce(N__68762),
            .sr(N__79586));
    defparam \ppm_encoder_1.pulses2count_esr_9_LC_15_4_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_9_LC_15_4_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_9_LC_15_4_2 .LUT_INIT=16'b0000010100000001;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_9_LC_15_4_2  (
            .in0(N__61779),
            .in1(N__64437),
            .in2(N__60636),
            .in3(N__63498),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__86987),
            .ce(N__68762),
            .sr(N__79586));
    defparam \ppm_encoder_1.pulses2count_esr_18_LC_15_4_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_18_LC_15_4_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_18_LC_15_4_3 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_18_LC_15_4_3  (
            .in0(N__64435),
            .in1(N__60609),
            .in2(_gnd_net_),
            .in3(N__64584),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__86987),
            .ce(N__68762),
            .sr(N__79586));
    defparam \ppm_encoder_1.pulses2count_esr_10_LC_15_4_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_10_LC_15_4_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_10_LC_15_4_5 .LUT_INIT=16'b0000000000100011;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_10_LC_15_4_5  (
            .in0(N__60576),
            .in1(N__60543),
            .in2(N__64448),
            .in3(N__60768),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__86987),
            .ce(N__68762),
            .sr(N__79586));
    defparam \ppm_encoder_1.counter24_0_I_33_c_RNO_LC_15_4_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_33_c_RNO_LC_15_4_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_33_c_RNO_LC_15_4_6 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_33_c_RNO_LC_15_4_6  (
            .in0(N__60537),
            .in1(N__64753),
            .in2(N__64782),
            .in3(N__60531),
            .lcout(\ppm_encoder_1.counter24_0_I_33_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.ppm_output_reg_RNO_0_LC_15_5_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.ppm_output_reg_RNO_0_LC_15_5_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.ppm_output_reg_RNO_0_LC_15_5_1 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \ppm_encoder_1.ppm_output_reg_RNO_0_LC_15_5_1  (
            .in0(N__60480),
            .in1(N__65508),
            .in2(N__61242),
            .in3(N__61163),
            .lcout(\ppm_encoder_1.ppm_output_reg_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter_RNIQM6H_12_LC_15_5_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter_RNIQM6H_12_LC_15_5_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter_RNIQM6H_12_LC_15_5_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \ppm_encoder_1.counter_RNIQM6H_12_LC_15_5_2  (
            .in0(N__68555),
            .in1(N__65551),
            .in2(N__68517),
            .in3(N__65575),
            .lcout(\ppm_encoder_1.un1_PPM_STATE_0_sqmuxa_0_i_a2_18_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter_RNIS9KG_8_LC_15_5_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter_RNIS9KG_8_LC_15_5_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter_RNIS9KG_8_LC_15_5_3 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \ppm_encoder_1.counter_RNIS9KG_8_LC_15_5_3  (
            .in0(N__64780),
            .in1(N__64802),
            .in2(N__64758),
            .in3(N__64823),
            .lcout(),
            .ltout(\ppm_encoder_1.un1_PPM_STATE_0_sqmuxa_0_i_a2_18_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter_RNIG7H22_2_LC_15_5_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter_RNIG7H22_2_LC_15_5_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter_RNIG7H22_2_LC_15_5_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \ppm_encoder_1.counter_RNIG7H22_2_LC_15_5_4  (
            .in0(N__60501),
            .in1(N__68394),
            .in2(N__60489),
            .in3(N__60486),
            .lcout(\ppm_encoder_1.N_486_18 ),
            .ltout(\ppm_encoder_1.N_486_18_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter_RNI09RH2_18_LC_15_5_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter_RNI09RH2_18_LC_15_5_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter_RNI09RH2_18_LC_15_5_5 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \ppm_encoder_1.counter_RNI09RH2_18_LC_15_5_5  (
            .in0(N__61238),
            .in1(N__65509),
            .in2(N__61221),
            .in3(N__61217),
            .lcout(\ppm_encoder_1.counter_RNI09RH2Z0Z_18 ),
            .ltout(\ppm_encoder_1.counter_RNI09RH2Z0Z_18_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNIGCO83_LC_15_5_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNIGCO83_LC_15_5_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNIGCO83_LC_15_5_6 .LUT_INIT=16'b1111111111110010;
    LogicCell40 \ppm_encoder_1.counter24_0_I_57_c_RNIGCO83_LC_15_5_6  (
            .in0(N__61164),
            .in1(N__61110),
            .in2(N__61083),
            .in3(N__66037),
            .lcout(\ppm_encoder_1.counter24_0_I_57_c_RNIGCOZ0Z83 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIJAMT_17_LC_15_6_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIJAMT_17_LC_15_6_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIJAMT_17_LC_15_6_1 .LUT_INIT=16'b1111000001111000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIJAMT_17_LC_15_6_1  (
            .in0(N__63438),
            .in1(N__64576),
            .in2(N__64635),
            .in3(N__64290),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_3_rep2_RNIA6041_LC_15_6_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_3_rep2_RNIA6041_LC_15_6_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_3_rep2_RNIA6041_LC_15_6_2 .LUT_INIT=16'b1110111010101010;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_3_rep2_RNIA6041_LC_15_6_2  (
            .in0(N__61014),
            .in1(N__60925),
            .in2(_gnd_net_),
            .in3(N__63860),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_3_rep2_RNIAZ0Z6041 ),
            .ltout(\ppm_encoder_1.CHOOSE_CHANNEL_3_rep2_RNIAZ0Z6041_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_10_LC_15_6_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_10_LC_15_6_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_10_LC_15_6_3 .LUT_INIT=16'b1111110011111110;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_10_LC_15_6_3  (
            .in0(N__63441),
            .in1(N__60723),
            .in2(N__60801),
            .in3(N__60794),
            .lcout(\ppm_encoder_1.pulses2count_9_i_0_2_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_10_LC_15_6_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_10_LC_15_6_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_10_LC_15_6_4 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_10_LC_15_6_4  (
            .in0(N__60758),
            .in1(N__61420),
            .in2(_gnd_net_),
            .in3(N__61639),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_2Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_8_LC_15_6_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_8_LC_15_6_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_8_LC_15_6_5 .LUT_INIT=16'b0000000000001010;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_8_LC_15_6_5  (
            .in0(N__61640),
            .in1(_gnd_net_),
            .in2(N__61448),
            .in3(N__60717),
            .lcout(),
            .ltout(\ppm_encoder_1.pulses2count_esr_RNO_2Z0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_8_LC_15_6_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_8_LC_15_6_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_8_LC_15_6_6 .LUT_INIT=16'b1111111111110100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_8_LC_15_6_6  (
            .in0(N__60684),
            .in1(N__63439),
            .in2(N__60651),
            .in3(N__61836),
            .lcout(\ppm_encoder_1.pulses2count_9_i_2_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_9_LC_15_6_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_9_LC_15_6_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_9_LC_15_6_7 .LUT_INIT=16'b1111110011111110;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_9_LC_15_6_7  (
            .in0(N__63440),
            .in1(N__61869),
            .in2(N__61851),
            .in3(N__61809),
            .lcout(\ppm_encoder_1.pulses2count_9_i_2_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_6_LC_15_7_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_6_LC_15_7_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_6_LC_15_7_1 .LUT_INIT=16'b0101100000001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_6_LC_15_7_1  (
            .in0(N__61626),
            .in1(N__61766),
            .in2(N__61450),
            .in3(N__61731),
            .lcout(\ppm_encoder_1.pulses2count_9_0_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_6_LC_15_7_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_6_LC_15_7_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_6_LC_15_7_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_6_LC_15_7_4  (
            .in0(_gnd_net_),
            .in1(N__64431),
            .in2(_gnd_net_),
            .in3(N__61695),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_2Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_13_LC_15_7_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_13_LC_15_7_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_13_LC_15_7_5 .LUT_INIT=16'b0101100000001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_13_LC_15_7_5  (
            .in0(N__61625),
            .in1(N__61488),
            .in2(N__61449),
            .in3(N__61308),
            .lcout(\ppm_encoder_1.pulses2count_9_0_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un11lto30_i_a2_0_c_LC_15_8_0 .C_ON=1'b1;
    defparam \pid_side.un11lto30_i_a2_0_c_LC_15_8_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.un11lto30_i_a2_0_c_LC_15_8_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_side.un11lto30_i_a2_0_c_LC_15_8_0  (
            .in0(_gnd_net_),
            .in1(N__61275),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_8_0_),
            .carryout(\pid_side.un11lto30_i_a2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un11lto30_i_a2_1_c_LC_15_8_1 .C_ON=1'b1;
    defparam \pid_side.un11lto30_i_a2_1_c_LC_15_8_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.un11lto30_i_a2_1_c_LC_15_8_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_side.un11lto30_i_a2_1_c_LC_15_8_1  (
            .in0(_gnd_net_),
            .in1(N__61269),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pid_side.un11lto30_i_a2 ),
            .carryout(\pid_side.un11lto30_i_a2_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un11lto30_i_a2_2_c_LC_15_8_2 .C_ON=1'b1;
    defparam \pid_side.un11lto30_i_a2_2_c_LC_15_8_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.un11lto30_i_a2_2_c_LC_15_8_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_side.un11lto30_i_a2_2_c_LC_15_8_2  (
            .in0(_gnd_net_),
            .in1(N__61263),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pid_side.un11lto30_i_a2_0 ),
            .carryout(\pid_side.un11lto30_i_a2_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un11lto30_i_a2_3_c_LC_15_8_3 .C_ON=1'b1;
    defparam \pid_side.un11lto30_i_a2_3_c_LC_15_8_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.un11lto30_i_a2_3_c_LC_15_8_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_side.un11lto30_i_a2_3_c_LC_15_8_3  (
            .in0(_gnd_net_),
            .in1(N__61251),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pid_side.un11lto30_i_a2_1 ),
            .carryout(\pid_side.un11lto30_i_a2_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un11lto30_i_a2_4_c_LC_15_8_4 .C_ON=1'b1;
    defparam \pid_side.un11lto30_i_a2_4_c_LC_15_8_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.un11lto30_i_a2_4_c_LC_15_8_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_side.un11lto30_i_a2_4_c_LC_15_8_4  (
            .in0(_gnd_net_),
            .in1(N__72735),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pid_side.un11lto30_i_a2_2 ),
            .carryout(\pid_side.un11lto30_i_a2_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un11lto30_i_a2_5_c_LC_15_8_5 .C_ON=1'b1;
    defparam \pid_side.un11lto30_i_a2_5_c_LC_15_8_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.un11lto30_i_a2_5_c_LC_15_8_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_side.un11lto30_i_a2_5_c_LC_15_8_5  (
            .in0(_gnd_net_),
            .in1(N__61916),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pid_side.un11lto30_i_a2_3 ),
            .carryout(\pid_side.un11lto30_i_a2_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un11lto30_i_a2_6_c_LC_15_8_6 .C_ON=1'b1;
    defparam \pid_side.un11lto30_i_a2_6_c_LC_15_8_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.un11lto30_i_a2_6_c_LC_15_8_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_side.un11lto30_i_a2_6_c_LC_15_8_6  (
            .in0(_gnd_net_),
            .in1(N__61941),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pid_side.un11lto30_i_a2_4 ),
            .carryout(\pid_side.un11lto30_i_a2_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un11lto30_i_a2_7_c_LC_15_8_7 .C_ON=1'b1;
    defparam \pid_side.un11lto30_i_a2_7_c_LC_15_8_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.un11lto30_i_a2_7_c_LC_15_8_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_side.un11lto30_i_a2_7_c_LC_15_8_7  (
            .in0(_gnd_net_),
            .in1(N__61935),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pid_side.un11lto30_i_a2_5 ),
            .carryout(\pid_side.un11lto30_i_a2_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un11lto30_i_a2_7_c_RNILAF8_LC_15_9_0 .C_ON=1'b0;
    defparam \pid_side.un11lto30_i_a2_7_c_RNILAF8_LC_15_9_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.un11lto30_i_a2_7_c_RNILAF8_LC_15_9_0 .LUT_INIT=16'b0000100000001111;
    LogicCell40 \pid_side.un11lto30_i_a2_7_c_RNILAF8_LC_15_9_0  (
            .in0(N__71711),
            .in1(N__69500),
            .in2(N__70011),
            .in3(N__61962),
            .lcout(\pid_side.source_pid_1_sqmuxa_1_0_o2_sx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_esr_RNIEHAB5_0_LC_15_9_2 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_esr_RNIEHAB5_0_LC_15_9_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_esr_RNIEHAB5_0_LC_15_9_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \pid_side.pid_prereg_esr_RNIEHAB5_0_LC_15_9_2  (
            .in0(N__61947),
            .in1(N__71591),
            .in2(N__68382),
            .in3(N__61889),
            .lcout(\pid_side.N_389 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_esr_RNIQVTS_0_LC_15_9_3 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_esr_RNIQVTS_0_LC_15_9_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_esr_RNIQVTS_0_LC_15_9_3 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \pid_side.pid_prereg_esr_RNIQVTS_0_LC_15_9_3  (
            .in0(N__69499),
            .in1(N__69412),
            .in2(_gnd_net_),
            .in3(N__69194),
            .lcout(\pid_side.source_pid_1_sqmuxa_1_0_a4_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_esr_RNI2L63_24_LC_15_9_6 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_esr_RNI2L63_24_LC_15_9_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_esr_RNI2L63_24_LC_15_9_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_side.pid_prereg_esr_RNI2L63_24_LC_15_9_6  (
            .in0(N__69606),
            .in1(N__69639),
            .in2(N__69576),
            .in3(N__69678),
            .lcout(\pid_side.un11lto30_i_a2_5_and ),
            .ltout(\pid_side.un11lto30_i_a2_5_and_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_esr_RNI9ACR_15_LC_15_9_7 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_esr_RNI9ACR_15_LC_15_9_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_esr_RNI9ACR_15_LC_15_9_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \pid_side.pid_prereg_esr_RNI9ACR_15_LC_15_9_7  (
            .in0(N__61934),
            .in1(N__72669),
            .in2(N__61920),
            .in3(N__61917),
            .lcout(\pid_side.N_98 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_10_LC_15_10_6 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_10_LC_15_10_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_10_LC_15_10_6 .LUT_INIT=16'b1100110010100000;
    LogicCell40 \pid_side.error_i_acumm_10_LC_15_10_6  (
            .in0(N__65928),
            .in1(N__62007),
            .in2(N__72641),
            .in3(N__65894),
            .lcout(\pid_side.error_i_acummZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87032),
            .ce(N__66107),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_3_LC_15_11_0 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_3_LC_15_11_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_3_LC_15_11_0 .LUT_INIT=16'b1111001000000010;
    LogicCell40 \pid_side.error_i_acumm_3_LC_15_11_0  (
            .in0(N__72620),
            .in1(N__66043),
            .in2(N__65895),
            .in3(N__65829),
            .lcout(\pid_side.error_i_acummZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87042),
            .ce(N__66100),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_1_LC_15_11_1 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_1_LC_15_11_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_1_LC_15_11_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \pid_side.error_i_acumm_1_LC_15_11_1  (
            .in0(_gnd_net_),
            .in1(N__65664),
            .in2(_gnd_net_),
            .in3(N__65884),
            .lcout(\pid_side.error_i_acummZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87042),
            .ce(N__66100),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_RNI6B4A1_0_LC_15_11_2 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_RNI6B4A1_0_LC_15_11_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_acumm_prereg_esr_RNI6B4A1_0_LC_15_11_2 .LUT_INIT=16'b1111111000000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_RNI6B4A1_0_LC_15_11_2  (
            .in0(N__65663),
            .in1(N__62246),
            .in2(N__65655),
            .in3(N__65828),
            .lcout(\pid_side.un10lt9_1 ),
            .ltout(\pid_side.un10lt9_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_RNIDUN92_0_4_LC_15_11_3 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIDUN92_0_4_LC_15_11_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIDUN92_0_4_LC_15_11_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_RNIDUN92_0_4_LC_15_11_3  (
            .in0(N__66125),
            .in1(N__68989),
            .in2(N__61992),
            .in3(N__65743),
            .lcout(\pid_side.error_i_acumm16lt9_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_2_LC_15_11_4 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_2_LC_15_11_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_2_LC_15_11_4 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \pid_side.error_i_acumm_2_LC_15_11_4  (
            .in0(N__65885),
            .in1(N__65654),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_i_acummZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87042),
            .ce(N__66100),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_RNIDUN92_4_LC_15_11_5 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIDUN92_4_LC_15_11_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIDUN92_4_LC_15_11_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_RNIDUN92_4_LC_15_11_5  (
            .in0(N__68990),
            .in1(N__65744),
            .in2(N__66129),
            .in3(N__61983),
            .lcout(),
            .ltout(\pid_side.un10lt9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_RNITQB93_7_LC_15_11_6 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_RNITQB93_7_LC_15_11_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_acumm_prereg_esr_RNITQB93_7_LC_15_11_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_RNITQB93_7_LC_15_11_6  (
            .in0(N__62264),
            .in1(N__65794),
            .in2(N__61977),
            .in3(N__62282),
            .lcout(),
            .ltout(\pid_side.un10lt11_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_RNIGIQP9_12_LC_15_11_7 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIGIQP9_12_LC_15_11_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIGIQP9_12_LC_15_11_7 .LUT_INIT=16'b0101010011111111;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_RNIGIQP9_12_LC_15_11_7  (
            .in0(N__68366),
            .in1(N__61974),
            .in2(N__61965),
            .in3(N__65637),
            .lcout(\pid_side.error_i_acumm_prereg_esr_RNIGIQP9Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_12_LC_15_12_0 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_12_LC_15_12_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_12_LC_15_12_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \pid_side.error_i_acumm_12_LC_15_12_0  (
            .in0(N__72519),
            .in1(N__68367),
            .in2(_gnd_net_),
            .in3(N__65890),
            .lcout(\pid_side.error_i_acummZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87051),
            .ce(N__66093),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_7_LC_15_12_1 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_7_LC_15_12_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_7_LC_15_12_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \pid_side.error_i_acumm_7_LC_15_12_1  (
            .in0(N__65891),
            .in1(N__72521),
            .in2(_gnd_net_),
            .in3(N__62283),
            .lcout(\pid_side.error_i_acummZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87051),
            .ce(N__66093),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_8_LC_15_12_2 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_8_LC_15_12_2 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_8_LC_15_12_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \pid_side.error_i_acumm_8_LC_15_12_2  (
            .in0(N__72520),
            .in1(N__62265),
            .in2(_gnd_net_),
            .in3(N__65892),
            .lcout(\pid_side.error_i_acummZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87051),
            .ce(N__66093),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_9_LC_15_12_3 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_9_LC_15_12_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_9_LC_15_12_3 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \pid_side.error_i_acumm_9_LC_15_12_3  (
            .in0(N__65893),
            .in1(_gnd_net_),
            .in2(N__65805),
            .in3(N__72522),
            .lcout(\pid_side.error_i_acummZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87051),
            .ce(N__66093),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_0_LC_15_12_4 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_0_LC_15_12_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_0_LC_15_12_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \pid_side.error_i_acumm_0_LC_15_12_4  (
            .in0(_gnd_net_),
            .in1(N__62247),
            .in2(_gnd_net_),
            .in3(N__65889),
            .lcout(\pid_side.error_i_acummZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87051),
            .ce(N__66093),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNIS1ID3_7_LC_15_12_5 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIS1ID3_7_LC_15_12_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIS1ID3_7_LC_15_12_5 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_side.error_p_reg_esr_RNIS1ID3_7_LC_15_12_5  (
            .in0(N__62229),
            .in1(N__62214),
            .in2(_gnd_net_),
            .in3(N__66467),
            .lcout(\pid_side.error_p_reg_esr_RNIS1ID3Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.data_Aux_RNO_0_0_LC_15_12_7 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_RNO_0_0_LC_15_12_7 .SEQ_MODE=4'b0000;
    defparam \uart_drone.data_Aux_RNO_0_0_LC_15_12_7 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \uart_drone.data_Aux_RNO_0_0_LC_15_12_7  (
            .in0(N__62208),
            .in1(N__62145),
            .in2(_gnd_net_),
            .in3(N__62085),
            .lcout(\uart_drone.data_Auxce_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_0_0_c_RNI3DS82_LC_15_13_0 .C_ON=1'b0;
    defparam \pid_side.error_cry_0_0_c_RNI3DS82_LC_15_13_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_0_0_c_RNI3DS82_LC_15_13_0 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \pid_side.error_cry_0_0_c_RNI3DS82_LC_15_13_0  (
            .in0(N__76009),
            .in1(N__75074),
            .in2(_gnd_net_),
            .in3(N__75904),
            .lcout(\pid_side.N_27_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_0_c_RNIRRMQ1_LC_15_13_1 .C_ON=1'b0;
    defparam \pid_side.error_cry_0_c_RNIRRMQ1_LC_15_13_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_0_c_RNIRRMQ1_LC_15_13_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \pid_side.error_cry_0_c_RNIRRMQ1_LC_15_13_1  (
            .in0(N__80944),
            .in1(N__62496),
            .in2(_gnd_net_),
            .in3(N__62334),
            .lcout(\pid_side.N_15_0 ),
            .ltout(\pid_side.N_15_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_0_16_LC_15_13_2 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_0_16_LC_15_13_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_0_16_LC_15_13_2 .LUT_INIT=16'b0100010000000101;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_0_16_LC_15_13_2  (
            .in0(N__76242),
            .in1(N__80222),
            .in2(N__62010),
            .in3(N__71559),
            .lcout(),
            .ltout(\pid_side.m4_2_03_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_16_LC_15_13_3 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_16_LC_15_13_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_esr_16_LC_15_13_3 .LUT_INIT=16'b1000000011000100;
    LogicCell40 \pid_side.error_i_reg_esr_16_LC_15_13_3  (
            .in0(N__76864),
            .in1(N__76659),
            .in2(N__62337),
            .in3(N__66891),
            .lcout(\pid_side.error_i_regZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87060),
            .ce(N__75290),
            .sr(N__79644));
    defparam \pid_side.error_i_reg_esr_0_LC_15_13_4 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_0_LC_15_13_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_esr_0_LC_15_13_4 .LUT_INIT=16'b1000100000001010;
    LogicCell40 \pid_side.error_i_reg_esr_0_LC_15_13_4  (
            .in0(N__70968),
            .in1(N__80223),
            .in2(N__67107),
            .in3(N__71561),
            .lcout(\pid_side.error_i_regZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87060),
            .ce(N__75290),
            .sr(N__79644));
    defparam \pid_side.error_cry_2_c_RNIB5P21_LC_15_13_5 .C_ON=1'b0;
    defparam \pid_side.error_cry_2_c_RNIB5P21_LC_15_13_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_2_c_RNIB5P21_LC_15_13_5 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \pid_side.error_cry_2_c_RNIB5P21_LC_15_13_5  (
            .in0(N__76010),
            .in1(N__75193),
            .in2(_gnd_net_),
            .in3(N__75023),
            .lcout(\pid_side.N_30_1 ),
            .ltout(\pid_side.N_30_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_2_c_RNIIVPE3_LC_15_13_6 .C_ON=1'b0;
    defparam \pid_side.error_cry_2_c_RNIIVPE3_LC_15_13_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_2_c_RNIIVPE3_LC_15_13_6 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \pid_side.error_cry_2_c_RNIIVPE3_LC_15_13_6  (
            .in0(_gnd_net_),
            .in1(N__80943),
            .in2(N__62328),
            .in3(N__62603),
            .lcout(\pid_side.N_63 ),
            .ltout(\pid_side.N_63_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_2_LC_15_13_7 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_2_LC_15_13_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_esr_2_LC_15_13_7 .LUT_INIT=16'b1000110000000100;
    LogicCell40 \pid_side.error_i_reg_esr_2_LC_15_13_7  (
            .in0(N__71560),
            .in1(N__70969),
            .in2(N__62325),
            .in3(N__62322),
            .lcout(\pid_side.error_i_regZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87060),
            .ce(N__75290),
            .sr(N__79644));
    defparam \pid_side.error_d_reg_prev_esr_RNI1FKL1_0_22_LC_15_14_0 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI1FKL1_0_22_LC_15_14_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI1FKL1_0_22_LC_15_14_0 .LUT_INIT=16'b0001100011100111;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI1FKL1_0_22_LC_15_14_0  (
            .in0(N__84593),
            .in1(N__83569),
            .in2(N__73212),
            .in3(N__66841),
            .lcout(\pid_side.un1_pid_prereg_0_23 ),
            .ltout(\pid_side.un1_pid_prereg_0_23_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI0R7B3_22_LC_15_14_1 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI0R7B3_22_LC_15_14_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI0R7B3_22_LC_15_14_1 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI0R7B3_22_LC_15_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__62289),
            .in3(N__62378),
            .lcout(\pid_side.error_d_reg_prev_esr_RNI0R7B3Z0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIVBJL1_22_LC_15_14_2 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIVBJL1_22_LC_15_14_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIVBJL1_22_LC_15_14_2 .LUT_INIT=16'b1110111100001000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIVBJL1_22_LC_15_14_2  (
            .in0(N__84592),
            .in1(N__83568),
            .in2(N__73211),
            .in3(N__72828),
            .lcout(\pid_side.un1_pid_prereg_0_22 ),
            .ltout(\pid_side.un1_pid_prereg_0_22_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNISFDM6_22_LC_15_14_3 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNISFDM6_22_LC_15_14_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNISFDM6_22_LC_15_14_3 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNISFDM6_22_LC_15_14_3  (
            .in0(N__73239),
            .in1(N__62387),
            .in2(N__62286),
            .in3(N__72795),
            .lcout(\pid_side.error_d_reg_prev_esr_RNISFDM6Z0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI2HLL1_0_22_LC_15_14_4 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI2HLL1_0_22_LC_15_14_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI2HLL1_0_22_LC_15_14_4 .LUT_INIT=16'b0001100011100111;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI2HLL1_0_22_LC_15_14_4  (
            .in0(N__84591),
            .in1(N__83567),
            .in2(N__73210),
            .in3(N__66723),
            .lcout(\pid_side.un1_pid_prereg_0_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI1FKL1_22_LC_15_14_5 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI1FKL1_22_LC_15_14_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI1FKL1_22_LC_15_14_5 .LUT_INIT=16'b1011101010100010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI1FKL1_22_LC_15_14_5  (
            .in0(N__66842),
            .in1(N__73204),
            .in2(N__83574),
            .in3(N__84594),
            .lcout(\pid_side.un1_pid_prereg_0_24 ),
            .ltout(\pid_side.un1_pid_prereg_0_24_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI3RHM6_22_LC_15_14_6 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI3RHM6_22_LC_15_14_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI3RHM6_22_LC_15_14_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI3RHM6_22_LC_15_14_6  (
            .in0(N__62388),
            .in1(N__62379),
            .in2(N__62367),
            .in3(N__66286),
            .lcout(\pid_side.error_d_reg_prev_esr_RNI3RHM6Z0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI30AB3_22_LC_15_14_7 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI30AB3_22_LC_15_14_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI30AB3_22_LC_15_14_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI30AB3_22_LC_15_14_7  (
            .in0(N__66287),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__66323),
            .lcout(\pid_side.error_d_reg_prev_esr_RNI30AB3Z0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_1_c_RNIGFRK_LC_15_15_0 .C_ON=1'b0;
    defparam \pid_side.error_cry_1_c_RNIGFRK_LC_15_15_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_1_c_RNIGFRK_LC_15_15_0 .LUT_INIT=16'b0100010001110111;
    LogicCell40 \pid_side.error_cry_1_c_RNIGFRK_LC_15_15_0  (
            .in0(N__75129),
            .in1(N__75997),
            .in2(_gnd_net_),
            .in3(N__75192),
            .lcout(\pid_side.N_11_0 ),
            .ltout(\pid_side.N_11_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_0_c_RNI622C1_LC_15_15_1 .C_ON=1'b0;
    defparam \pid_side.error_cry_0_c_RNI622C1_LC_15_15_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_0_c_RNI622C1_LC_15_15_1 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \pid_side.error_cry_0_c_RNI622C1_LC_15_15_1  (
            .in0(N__80939),
            .in1(_gnd_net_),
            .in2(N__62364),
            .in3(N__62477),
            .lcout(\pid_side.N_15_1 ),
            .ltout(\pid_side.N_15_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_0_15_LC_15_15_2 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_0_15_LC_15_15_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_0_15_LC_15_15_2 .LUT_INIT=16'b0000000000000011;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_0_15_LC_15_15_2  (
            .in0(_gnd_net_),
            .in1(N__75743),
            .in2(N__62361),
            .in3(N__71518),
            .lcout(\pid_side.m3_2_03 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_3_LC_15_15_3 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_3_LC_15_15_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_esr_3_LC_15_15_3 .LUT_INIT=16'b0010000001110000;
    LogicCell40 \pid_side.error_i_reg_esr_3_LC_15_15_3  (
            .in0(N__71519),
            .in1(N__62352),
            .in2(N__70980),
            .in3(N__62433),
            .lcout(\pid_side.error_i_regZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87080),
            .ce(N__75329),
            .sr(N__79660));
    defparam \pid_side.error_cry_0_c_RNII52K_LC_15_15_4 .C_ON=1'b0;
    defparam \pid_side.error_cry_0_c_RNII52K_LC_15_15_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_0_c_RNII52K_LC_15_15_4 .LUT_INIT=16'b0001000111011101;
    LogicCell40 \pid_side.error_cry_0_c_RNII52K_LC_15_15_4  (
            .in0(N__73868),
            .in1(N__75996),
            .in2(_gnd_net_),
            .in3(N__81047),
            .lcout(\pid_side.N_14_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_0_6_LC_15_15_5 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_0_6_LC_15_15_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_0_6_LC_15_15_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_0_6_LC_15_15_5  (
            .in0(N__80615),
            .in1(N__62566),
            .in2(_gnd_net_),
            .in3(N__62535),
            .lcout(),
            .ltout(\pid_side.N_110_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_6_LC_15_15_6 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_6_LC_15_15_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_esr_6_LC_15_15_6 .LUT_INIT=16'b1000100000001100;
    LogicCell40 \pid_side.error_i_reg_esr_6_LC_15_15_6  (
            .in0(N__62514),
            .in1(N__75475),
            .in2(N__62499),
            .in3(N__75744),
            .lcout(\pid_side.error_i_regZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87080),
            .ce(N__75329),
            .sr(N__79660));
    defparam \pid_side.error_cry_0_c_RNIC9PK_LC_15_15_7 .C_ON=1'b0;
    defparam \pid_side.error_cry_0_c_RNIC9PK_LC_15_15_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_0_c_RNIC9PK_LC_15_15_7 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \pid_side.error_cry_0_c_RNIC9PK_LC_15_15_7  (
            .in0(N__75995),
            .in1(N__73867),
            .in2(_gnd_net_),
            .in3(N__75128),
            .lcout(\pid_side.N_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_0_c_RNIC7AM1_LC_15_16_0 .C_ON=1'b0;
    defparam \pid_side.error_cry_0_c_RNIC7AM1_LC_15_16_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_0_c_RNIC7AM1_LC_15_16_0 .LUT_INIT=16'b0000001000000111;
    LogicCell40 \pid_side.error_cry_0_c_RNIC7AM1_LC_15_16_0  (
            .in0(N__71988),
            .in1(N__62478),
            .in2(N__80616),
            .in3(N__67043),
            .lcout(\pid_side.N_104 ),
            .ltout(\pid_side.N_104_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_2_23_LC_15_16_1 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_2_23_LC_15_16_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_2_23_LC_15_16_1 .LUT_INIT=16'b0001101100011011;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_2_23_LC_15_16_1  (
            .in0(N__75718),
            .in1(N__80607),
            .in2(N__62460),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\pid_side.un4_error_i_reg_33_bm_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_1_23_LC_15_16_2 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_1_23_LC_15_16_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_1_23_LC_15_16_2 .LUT_INIT=16'b0001101000011111;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_1_23_LC_15_16_2  (
            .in0(N__75748),
            .in1(N__62457),
            .in2(N__62436),
            .in3(N__62432),
            .lcout(),
            .ltout(\pid_side.error_i_reg_esr_RNO_1Z0Z_23_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_23_LC_15_16_3 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_23_LC_15_16_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_esr_23_LC_15_16_3 .LUT_INIT=16'b1100010010000000;
    LogicCell40 \pid_side.error_i_reg_esr_23_LC_15_16_3  (
            .in0(N__76945),
            .in1(N__76615),
            .in2(N__62406),
            .in3(N__62619),
            .lcout(\pid_side.error_i_regZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87094),
            .ce(N__75331),
            .sr(N__79667));
    defparam \pid_side.error_cry_9_c_RNIL6R82_0_LC_15_16_4 .C_ON=1'b0;
    defparam \pid_side.error_cry_9_c_RNIL6R82_0_LC_15_16_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_9_c_RNIL6R82_0_LC_15_16_4 .LUT_INIT=16'b0000001100010001;
    LogicCell40 \pid_side.error_cry_9_c_RNIL6R82_0_LC_15_16_4  (
            .in0(N__74884),
            .in1(N__71987),
            .in2(N__74419),
            .in3(N__80755),
            .lcout(),
            .ltout(\pid_side.error_cry_9_c_RNIL6R82Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_7_c_RNI53TC7_LC_15_16_5 .C_ON=1'b0;
    defparam \pid_side.error_cry_7_c_RNI53TC7_LC_15_16_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_7_c_RNI53TC7_LC_15_16_5 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \pid_side.error_cry_7_c_RNI53TC7_LC_15_16_5  (
            .in0(_gnd_net_),
            .in1(N__62664),
            .in2(N__62403),
            .in3(N__62613),
            .lcout(\pid_side.N_46_1 ),
            .ltout(\pid_side.N_46_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_0_23_LC_15_16_6 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_0_23_LC_15_16_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_0_23_LC_15_16_6 .LUT_INIT=16'b0010111010101010;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_0_23_LC_15_16_6  (
            .in0(N__74885),
            .in1(N__75717),
            .in2(N__62622),
            .in3(N__71530),
            .lcout(\pid_side.error_i_reg_esr_RNO_0Z0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_9_c_RNIL6R82_LC_15_16_7 .C_ON=1'b0;
    defparam \pid_side.error_cry_9_c_RNIL6R82_LC_15_16_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_9_c_RNIL6R82_LC_15_16_7 .LUT_INIT=16'b1111001011110111;
    LogicCell40 \pid_side.error_cry_9_c_RNIL6R82_LC_15_16_7  (
            .in0(N__80754),
            .in1(N__74409),
            .in2(N__72032),
            .in3(N__74883),
            .lcout(\pid_side.error_cry_9_c_RNIL6RZ0Z82 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_3_0_c_RNIJIPS1_0_LC_15_17_0 .C_ON=1'b0;
    defparam \pid_side.error_cry_3_0_c_RNIJIPS1_0_LC_15_17_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_3_0_c_RNIJIPS1_0_LC_15_17_0 .LUT_INIT=16'b0000000100001101;
    LogicCell40 \pid_side.error_cry_3_0_c_RNIJIPS1_0_LC_15_17_0  (
            .in0(N__74756),
            .in1(N__76005),
            .in2(N__80971),
            .in3(N__75811),
            .lcout(\pid_side.error_cry_3_0_c_RNIJIPS1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_3_0_c_RNIJIPS1_LC_15_17_1 .C_ON=1'b0;
    defparam \pid_side.error_cry_3_0_c_RNIJIPS1_LC_15_17_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_3_0_c_RNIJIPS1_LC_15_17_1 .LUT_INIT=16'b1101110011011111;
    LogicCell40 \pid_side.error_cry_3_0_c_RNIJIPS1_LC_15_17_1  (
            .in0(N__75812),
            .in1(N__80938),
            .in2(N__76011),
            .in3(N__74757),
            .lcout(),
            .ltout(\pid_side.error_cry_3_0_c_RNIJIPSZ0Z1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_3_0_c_RNI9IF26_LC_15_17_2 .C_ON=1'b0;
    defparam \pid_side.error_cry_3_0_c_RNI9IF26_LC_15_17_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_3_0_c_RNI9IF26_LC_15_17_2 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \pid_side.error_cry_3_0_c_RNI9IF26_LC_15_17_2  (
            .in0(_gnd_net_),
            .in1(N__62607),
            .in2(N__62592),
            .in3(N__62589),
            .lcout(\pid_side.N_28_1 ),
            .ltout(\pid_side.N_28_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_0_c_RNI94F58_LC_15_17_3 .C_ON=1'b0;
    defparam \pid_side.error_cry_0_c_RNI94F58_LC_15_17_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_0_c_RNI94F58_LC_15_17_3 .LUT_INIT=16'b0000010110101111;
    LogicCell40 \pid_side.error_cry_0_c_RNI94F58_LC_15_17_3  (
            .in0(N__80475),
            .in1(_gnd_net_),
            .in2(N__62583),
            .in3(N__67108),
            .lcout(\pid_side.error_cry_0_c_RNI94FZ0Z58 ),
            .ltout(\pid_side.error_cry_0_c_RNI94FZ0Z58_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_0_20_LC_15_17_4 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_0_20_LC_15_17_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_0_20_LC_15_17_4 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_0_20_LC_15_17_4  (
            .in0(_gnd_net_),
            .in1(N__76271),
            .in2(N__62580),
            .in3(N__67434),
            .lcout(),
            .ltout(\pid_side.m8_2_03_3_i_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_20_LC_15_17_5 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_20_LC_15_17_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_esr_20_LC_15_17_5 .LUT_INIT=16'b1000000011000100;
    LogicCell40 \pid_side.error_i_reg_esr_20_LC_15_17_5  (
            .in0(N__76944),
            .in1(N__76581),
            .in2(N__62577),
            .in3(N__62574),
            .lcout(\pid_side.error_i_regZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87110),
            .ce(N__75330),
            .sr(N__79674));
    defparam \pid_side.error_i_reg_esr_RNO_1_20_LC_15_17_6 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_1_20_LC_15_17_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_1_20_LC_15_17_6 .LUT_INIT=16'b1111111100100000;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_1_20_LC_15_17_6  (
            .in0(N__71974),
            .in1(N__74322),
            .in2(N__80383),
            .in3(N__62676),
            .lcout(\pid_side.m24_2_03_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_7_20_LC_15_18_0 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_7_20_LC_15_18_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_7_20_LC_15_18_0 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_7_20_LC_15_18_0  (
            .in0(N__67569),
            .in1(N__77890),
            .in2(_gnd_net_),
            .in3(N__77406),
            .lcout(),
            .ltout(\pid_side.G_5_0_a5_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_5_20_LC_15_18_1 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_5_20_LC_15_18_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_5_20_LC_15_18_1 .LUT_INIT=16'b0101000000110000;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_5_20_LC_15_18_1  (
            .in0(N__74166),
            .in1(N__74056),
            .in2(N__62682),
            .in3(N__78418),
            .lcout(),
            .ltout(\pid_side.N_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_2_20_LC_15_18_2 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_2_20_LC_15_18_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_2_20_LC_15_18_2 .LUT_INIT=16'b1111000011111101;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_2_20_LC_15_18_2  (
            .in0(N__67570),
            .in1(N__62670),
            .in2(N__62679),
            .in3(N__74905),
            .lcout(\pid_side.G_5_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_4_20_LC_15_18_3 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_4_20_LC_15_18_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_4_20_LC_15_18_3 .LUT_INIT=16'b0000010100000101;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_4_20_LC_15_18_3  (
            .in0(N__77891),
            .in1(_gnd_net_),
            .in2(N__77412),
            .in3(_gnd_net_),
            .lcout(\pid_side.G_5_0_a5_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_7_12_LC_15_18_4 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_7_12_LC_15_18_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_7_12_LC_15_18_4 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_7_12_LC_15_18_4  (
            .in0(N__80704),
            .in1(N__74049),
            .in2(_gnd_net_),
            .in3(N__74164),
            .lcout(\pid_side.N_6_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_7_c_RNIRL6R2_LC_15_18_6 .C_ON=1'b0;
    defparam \pid_side.error_cry_7_c_RNIRL6R2_LC_15_18_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_7_c_RNIRL6R2_LC_15_18_6 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \pid_side.error_cry_7_c_RNIRL6R2_LC_15_18_6  (
            .in0(N__80702),
            .in1(N__74048),
            .in2(_gnd_net_),
            .in3(N__74489),
            .lcout(\pid_side.N_45_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_7_21_LC_15_18_7 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_7_21_LC_15_18_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_7_21_LC_15_18_7 .LUT_INIT=16'b0001001111010011;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_7_21_LC_15_18_7  (
            .in0(N__74165),
            .in1(N__80703),
            .in2(N__78104),
            .in3(N__74574),
            .lcout(\pid_side.m87_0_ns_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam GB_BUFFER_reset_system_g_THRU_LUT4_0_LC_15_19_0.C_ON=1'b0;
    defparam GB_BUFFER_reset_system_g_THRU_LUT4_0_LC_15_19_0.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_reset_system_g_THRU_LUT4_0_LC_15_19_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 GB_BUFFER_reset_system_g_THRU_LUT4_0_LC_15_19_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__79915),
            .lcout(GB_BUFFER_reset_system_g_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_3_12_LC_15_19_1 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_3_12_LC_15_19_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_3_12_LC_15_19_1 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_3_12_LC_15_19_1  (
            .in0(N__77761),
            .in1(N__62628),
            .in2(_gnd_net_),
            .in3(N__74904),
            .lcout(\pid_side.N_9_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_11_21_LC_15_19_3 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_11_21_LC_15_19_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_11_21_LC_15_19_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_11_21_LC_15_19_3  (
            .in0(N__80721),
            .in1(N__81057),
            .in2(_gnd_net_),
            .in3(N__73872),
            .lcout(),
            .ltout(\pid_side.g2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_6_21_LC_15_19_4 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_6_21_LC_15_19_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_6_21_LC_15_19_4 .LUT_INIT=16'b0000000000110000;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_6_21_LC_15_19_4  (
            .in0(_gnd_net_),
            .in1(N__77760),
            .in2(N__62751),
            .in3(N__71969),
            .lcout(\pid_side.N_117_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_3_17_LC_15_19_5 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_3_17_LC_15_19_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_3_17_LC_15_19_5 .LUT_INIT=16'b0000100000001011;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_3_17_LC_15_19_5  (
            .in0(N__70572),
            .in1(N__71517),
            .in2(N__76268),
            .in3(N__67019),
            .lcout(\pid_side.m5_2_03 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_2_25_LC_15_19_6 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_2_25_LC_15_19_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_2_25_LC_15_19_6 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_2_25_LC_15_19_6  (
            .in0(N__71516),
            .in1(N__71968),
            .in2(N__80774),
            .in3(N__76208),
            .lcout(\pid_front.error_i_reg_esr_RNO_2Z0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_2_LC_15_20_0 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_2_LC_15_20_0 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_esr_2_LC_15_20_0 .LUT_INIT=16'b1000000011010000;
    LogicCell40 \pid_front.error_i_reg_esr_2_LC_15_20_0  (
            .in0(N__71526),
            .in1(N__62829),
            .in2(N__70973),
            .in3(N__62786),
            .lcout(\pid_front.error_i_regZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87156),
            .ce(N__72413),
            .sr(N__79687));
    defparam \pid_front.error_i_reg_esr_3_LC_15_20_1 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_3_LC_15_20_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_esr_3_LC_15_20_1 .LUT_INIT=16'b0001101100000000;
    LogicCell40 \pid_front.error_i_reg_esr_3_LC_15_20_1  (
            .in0(N__71502),
            .in1(N__76095),
            .in2(N__76383),
            .in3(N__70957),
            .lcout(\pid_front.error_i_regZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87156),
            .ce(N__72413),
            .sr(N__79687));
    defparam \pid_side.error_cry_0_c_RNIODGI_LC_15_20_2 .C_ON=1'b0;
    defparam \pid_side.error_cry_0_c_RNIODGI_LC_15_20_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_0_c_RNIODGI_LC_15_20_2 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \pid_side.error_cry_0_c_RNIODGI_LC_15_20_2  (
            .in0(N__80738),
            .in1(N__81059),
            .in2(N__80973),
            .in3(N__73877),
            .lcout(\pid_side.m1_0_03 ),
            .ltout(\pid_side.m1_0_03_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_1_5_LC_15_20_3 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_1_5_LC_15_20_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_1_5_LC_15_20_3 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_1_5_LC_15_20_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__62712),
            .in3(N__71525),
            .lcout(\pid_side.N_117 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_2_17_LC_15_20_5 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_2_17_LC_15_20_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_2_17_LC_15_20_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_2_17_LC_15_20_5  (
            .in0(N__62709),
            .in1(N__62700),
            .in2(_gnd_net_),
            .in3(N__74906),
            .lcout(),
            .ltout(\pid_side.N_131_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_0_17_LC_15_20_6 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_0_17_LC_15_20_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_0_17_LC_15_20_6 .LUT_INIT=16'b1000110000000100;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_0_17_LC_15_20_6  (
            .in0(N__77024),
            .in1(N__76513),
            .in2(N__62691),
            .in3(N__62688),
            .lcout(\pid_side.error_i_reg_9_rn_1_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_0_0_c_RNIIEHM2_LC_15_21_0 .C_ON=1'b0;
    defparam \pid_front.error_cry_0_0_c_RNIIEHM2_LC_15_21_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_0_0_c_RNIIEHM2_LC_15_21_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \pid_front.error_cry_0_0_c_RNIIEHM2_LC_15_21_0  (
            .in0(N__78057),
            .in1(N__63161),
            .in2(_gnd_net_),
            .in3(N__62924),
            .lcout(\pid_front.N_63 ),
            .ltout(\pid_front.N_63_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_1_18_LC_15_21_1 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_1_18_LC_15_21_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_1_18_LC_15_21_1 .LUT_INIT=16'b0100010100000001;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_1_18_LC_15_21_1  (
            .in0(N__80363),
            .in1(N__77762),
            .in2(N__62847),
            .in3(N__62823),
            .lcout(),
            .ltout(\pid_front.m6_2_03_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_0_18_LC_15_21_2 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_0_18_LC_15_21_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_0_18_LC_15_21_2 .LUT_INIT=16'b1010001010000000;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_0_18_LC_15_21_2  (
            .in0(N__76558),
            .in1(N__77022),
            .in2(N__62844),
            .in3(N__71183),
            .lcout(\pid_front.error_i_reg_9_rn_0_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_0_0_c_RNIL4UN4_LC_15_21_3 .C_ON=1'b0;
    defparam \pid_front.error_cry_0_0_c_RNIL4UN4_LC_15_21_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_0_0_c_RNIL4UN4_LC_15_21_3 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \pid_front.error_cry_0_0_c_RNIL4UN4_LC_15_21_3  (
            .in0(N__77404),
            .in1(N__62822),
            .in2(_gnd_net_),
            .in3(N__62782),
            .lcout(\pid_front.N_41_0 ),
            .ltout(\pid_front.N_41_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_0_26_LC_15_21_4 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_0_26_LC_15_21_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_0_26_LC_15_21_4 .LUT_INIT=16'b1010001010000000;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_0_26_LC_15_21_4  (
            .in0(N__76559),
            .in1(N__77023),
            .in2(N__62754),
            .in3(N__71184),
            .lcout(\pid_front.error_i_reg_9_rn_0_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_0_0_c_RNI44H31_LC_15_21_5 .C_ON=1'b0;
    defparam \pid_front.error_cry_0_0_c_RNI44H31_LC_15_21_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_0_0_c_RNI44H31_LC_15_21_5 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \pid_front.error_cry_0_0_c_RNI44H31_LC_15_21_5  (
            .in0(N__78221),
            .in1(N__67726),
            .in2(_gnd_net_),
            .in3(N__67789),
            .lcout(\pid_front.N_27_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_2_c_RNIB1241_LC_15_21_6 .C_ON=1'b0;
    defparam \pid_front.error_cry_2_c_RNIB1241_LC_15_21_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_2_c_RNIB1241_LC_15_21_6 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \pid_front.error_cry_2_c_RNIB1241_LC_15_21_6  (
            .in0(N__78219),
            .in1(N__77067),
            .in2(_gnd_net_),
            .in3(N__67846),
            .lcout(\pid_front.N_30_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_0_0_c_RNISQ6J3_LC_15_21_7 .C_ON=1'b0;
    defparam \pid_front.error_cry_0_0_c_RNISQ6J3_LC_15_21_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_0_0_c_RNISQ6J3_LC_15_21_7 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \pid_front.error_cry_0_0_c_RNISQ6J3_LC_15_21_7  (
            .in0(N__70858),
            .in1(N__77763),
            .in2(_gnd_net_),
            .in3(N__71021),
            .lcout(\pid_front.N_93_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_2_12_LC_15_22_0 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_2_12_LC_15_22_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_2_12_LC_15_22_0 .LUT_INIT=16'b0000110001110111;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_2_12_LC_15_22_0  (
            .in0(N__62900),
            .in1(N__80364),
            .in2(N__63149),
            .in3(N__77737),
            .lcout(),
            .ltout(\pid_front.m129_0_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_1_12_LC_15_22_1 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_1_12_LC_15_22_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_1_12_LC_15_22_1 .LUT_INIT=16'b0000111110101100;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_1_12_LC_15_22_1  (
            .in0(N__63120),
            .in1(N__63097),
            .in2(N__63012),
            .in3(N__76280),
            .lcout(\pid_front.m16_2_03_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_3_0_c_RNIJ5832_LC_15_22_2 .C_ON=1'b0;
    defparam \pid_front.error_cry_3_0_c_RNIJ5832_LC_15_22_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_3_0_c_RNIJ5832_LC_15_22_2 .LUT_INIT=16'b1111001011110111;
    LogicCell40 \pid_front.error_cry_3_0_c_RNIJ5832_LC_15_22_2  (
            .in0(N__78208),
            .in1(N__67662),
            .in2(N__78093),
            .in3(N__62976),
            .lcout(\pid_front.error_cry_3_0_c_RNIJZ0Z5832 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_4_c_RNI46QMA_LC_15_22_3 .C_ON=1'b0;
    defparam \pid_front.error_cry_4_c_RNI46QMA_LC_15_22_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_4_c_RNI46QMA_LC_15_22_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \pid_front.error_cry_4_c_RNI46QMA_LC_15_22_3  (
            .in0(N__77394),
            .in1(N__62899),
            .in2(_gnd_net_),
            .in3(N__63096),
            .lcout(\pid_front.N_29_1 ),
            .ltout(\pid_front.N_29_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_1_24_LC_15_22_4 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_1_24_LC_15_22_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_1_24_LC_15_22_4 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_1_24_LC_15_22_4  (
            .in0(_gnd_net_),
            .in1(N__80365),
            .in2(N__62931),
            .in3(N__68063),
            .lcout(\pid_front.N_89_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_3_0_c_RNI76F08_LC_15_22_5 .C_ON=1'b0;
    defparam \pid_front.error_cry_3_0_c_RNI76F08_LC_15_22_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_3_0_c_RNI76F08_LC_15_22_5 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \pid_front.error_cry_3_0_c_RNI76F08_LC_15_22_5  (
            .in0(N__77736),
            .in1(N__63141),
            .in2(_gnd_net_),
            .in3(N__62898),
            .lcout(\pid_front.error_cry_3_0_c_RNI76FZ0Z08 ),
            .ltout(\pid_front.error_cry_3_0_c_RNI76FZ0Z08_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_0_20_LC_15_22_6 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_0_20_LC_15_22_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_0_20_LC_15_22_6 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_0_20_LC_15_22_6  (
            .in0(N__76279),
            .in1(_gnd_net_),
            .in2(N__62928),
            .in3(N__68249),
            .lcout(\pid_front.m8_2_03_3_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_3_0_c_RNIAF1A5_LC_15_22_7 .C_ON=1'b0;
    defparam \pid_front.error_cry_3_0_c_RNIAF1A5_LC_15_22_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_3_0_c_RNIAF1A5_LC_15_22_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \pid_front.error_cry_3_0_c_RNIAF1A5_LC_15_22_7  (
            .in0(N__62925),
            .in1(N__62913),
            .in2(_gnd_net_),
            .in3(N__62907),
            .lcout(\pid_front.N_28_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_0_LC_15_23_0 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_0_LC_15_23_0 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_esr_0_LC_15_23_0 .LUT_INIT=16'b1000000011010000;
    LogicCell40 \pid_front.error_i_reg_esr_0_LC_15_23_0  (
            .in0(N__71547),
            .in1(N__63077),
            .in2(N__70977),
            .in3(N__63148),
            .lcout(\pid_front.error_i_regZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87200),
            .ce(N__72414),
            .sr(N__79696));
    defparam \pid_front.error_cry_10_c_RNIMQN12_LC_15_23_2 .C_ON=1'b0;
    defparam \pid_front.error_cry_10_c_RNIMQN12_LC_15_23_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_10_c_RNIMQN12_LC_15_23_2 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \pid_front.error_cry_10_c_RNIMQN12_LC_15_23_2  (
            .in0(N__72040),
            .in1(N__62858),
            .in2(_gnd_net_),
            .in3(N__71174),
            .lcout(\pid_front.N_57_0 ),
            .ltout(\pid_front.N_57_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_0_24_LC_15_23_3 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_0_24_LC_15_23_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_0_24_LC_15_23_3 .LUT_INIT=16'b1101000101010101;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_0_24_LC_15_23_3  (
            .in0(N__71175),
            .in1(N__76282),
            .in2(N__63204),
            .in3(N__80603),
            .lcout(),
            .ltout(\pid_front.N_59_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_24_LC_15_23_4 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_24_LC_15_23_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_esr_24_LC_15_23_4 .LUT_INIT=16'b1000110000000100;
    LogicCell40 \pid_front.error_i_reg_esr_24_LC_15_23_4  (
            .in0(N__76979),
            .in1(N__76628),
            .in2(N__63201),
            .in3(N__63198),
            .lcout(\pid_front.error_i_regZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87200),
            .ce(N__72414),
            .sr(N__79696));
    defparam \pid_front.error_cry_0_c_RNIP4BI2_LC_15_23_5 .C_ON=1'b0;
    defparam \pid_front.error_cry_0_c_RNIP4BI2_LC_15_23_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_0_c_RNIP4BI2_LC_15_23_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \pid_front.error_cry_0_c_RNIP4BI2_LC_15_23_5  (
            .in0(N__78082),
            .in1(N__63177),
            .in2(_gnd_net_),
            .in3(N__63165),
            .lcout(\pid_front.N_15_0 ),
            .ltout(\pid_front.N_15_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_0_c_RNI20AR3_LC_15_23_6 .C_ON=1'b0;
    defparam \pid_front.error_cry_0_c_RNI20AR3_LC_15_23_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_0_c_RNI20AR3_LC_15_23_6 .LUT_INIT=16'b1100110000001111;
    LogicCell40 \pid_front.error_cry_0_c_RNI20AR3_LC_15_23_6  (
            .in0(_gnd_net_),
            .in1(N__63076),
            .in2(N__63123),
            .in3(N__77403),
            .lcout(\pid_front.N_32_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_2_20_LC_15_24_0 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_2_20_LC_15_24_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_2_20_LC_15_24_0 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_2_20_LC_15_24_0  (
            .in0(N__80378),
            .in1(N__77787),
            .in2(_gnd_net_),
            .in3(N__71168),
            .lcout(),
            .ltout(\pid_front.m138_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_1_20_LC_15_24_1 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_1_20_LC_15_24_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_1_20_LC_15_24_1 .LUT_INIT=16'b1101101011010000;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_1_20_LC_15_24_1  (
            .in0(N__76320),
            .in1(N__63119),
            .in2(N__63105),
            .in3(N__63102),
            .lcout(\pid_front.m24_2_03_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_0_12_LC_15_24_5 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_0_12_LC_15_24_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_0_12_LC_15_24_5 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_0_12_LC_15_24_5  (
            .in0(N__76321),
            .in1(N__71546),
            .in2(_gnd_net_),
            .in3(N__63078),
            .lcout(\pid_front.m0_2_03 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_20_LC_15_25_2 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_20_LC_15_25_2 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_esr_20_LC_15_25_2 .LUT_INIT=16'b1100010100000000;
    LogicCell40 \pid_front.error_i_reg_esr_20_LC_15_25_2  (
            .in0(N__63051),
            .in1(N__63045),
            .in2(N__77014),
            .in3(N__76642),
            .lcout(\pid_front.error_i_regZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87232),
            .ce(N__72390),
            .sr(N__79707));
    defparam \pid_front.error_i_reg_esr_26_LC_15_25_6 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_26_LC_15_25_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_esr_26_LC_15_25_6 .LUT_INIT=16'b0111011100100010;
    LogicCell40 \pid_front.error_i_reg_esr_26_LC_15_25_6  (
            .in0(N__68280),
            .in1(N__63024),
            .in2(_gnd_net_),
            .in3(N__63966),
            .lcout(\pid_front.error_i_regZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87232),
            .ce(N__72390),
            .sr(N__79707));
    defparam \ppm_encoder_1.pulses2count_esr_16_LC_16_1_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_16_LC_16_1_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_16_LC_16_1_2 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_16_LC_16_1_2  (
            .in0(N__63942),
            .in1(N__64504),
            .in2(_gnd_net_),
            .in3(N__64397),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__86976),
            .ce(N__68768),
            .sr(N__79573));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_3_LC_16_2_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_3_LC_16_2_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_3_LC_16_2_1 .LUT_INIT=16'b0000000010001101;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_3_LC_16_2_1  (
            .in0(N__64289),
            .in1(N__64487),
            .in2(N__63912),
            .in3(N__79998),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__86982),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNISSER_LC_16_2_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNISSER_LC_16_2_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNISSER_LC_16_2_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNISSER_LC_16_2_2  (
            .in0(_gnd_net_),
            .in1(N__63859),
            .in2(_gnd_net_),
            .in3(N__63805),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNISSERZ0 ),
            .ltout(\ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNISSERZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_1_LC_16_2_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_1_LC_16_2_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_1_LC_16_2_3 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_1_LC_16_2_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__63693),
            .in3(N__63689),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_0_LC_16_2_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_0_LC_16_2_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_0_LC_16_2_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_0_LC_16_2_4  (
            .in0(N__63645),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__64388),
            .lcout(),
            .ltout(\ppm_encoder_1.pulses2count_esr_RNO_2Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_0_LC_16_2_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_0_LC_16_2_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_0_LC_16_2_5 .LUT_INIT=16'b1111101011111110;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_0_LC_16_2_5  (
            .in0(N__63406),
            .in1(N__63621),
            .in2(N__63597),
            .in3(N__63590),
            .lcout(\ppm_encoder_1.pulses2count_9_0_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNI4LP01_9_LC_16_2_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI4LP01_9_LC_16_2_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI4LP01_9_LC_16_2_6 .LUT_INIT=16'b1010101001101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI4LP01_9_LC_16_2_6  (
            .in0(N__63504),
            .in1(N__63405),
            .in2(N__64520),
            .in3(N__64288),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_2_LC_16_2_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_2_LC_16_2_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_2_LC_16_2_7 .LUT_INIT=16'b1111110011111110;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_2_LC_16_2_7  (
            .in0(N__64389),
            .in1(N__63270),
            .in2(N__63258),
            .in3(N__63235),
            .lcout(\ppm_encoder_1.pulses2count_9_i_3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_1_c_RNO_LC_16_3_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_1_c_RNO_LC_16_3_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_1_c_RNO_LC_16_3_0 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_1_c_RNO_LC_16_3_0  (
            .in0(N__63988),
            .in1(N__64737),
            .in2(N__64683),
            .in3(N__64015),
            .lcout(\ppm_encoder_1.counter24_0_I_1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_1_LC_16_3_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_1_LC_16_3_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_1_LC_16_3_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_1_LC_16_3_1  (
            .in0(N__68815),
            .in1(N__64719),
            .in2(N__64704),
            .in3(N__64689),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__86988),
            .ce(N__68767),
            .sr(N__79587));
    defparam \ppm_encoder_1.pulses2count_esr_15_LC_16_3_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_15_LC_16_3_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_15_LC_16_3_3 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_15_LC_16_3_3  (
            .in0(N__64674),
            .in1(N__64582),
            .in2(_gnd_net_),
            .in3(N__64395),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__86988),
            .ce(N__68767),
            .sr(N__79587));
    defparam \ppm_encoder_1.pulses2count_esr_17_LC_16_3_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_17_LC_16_3_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_17_LC_16_3_5 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_17_LC_16_3_5  (
            .in0(N__64634),
            .in1(N__64583),
            .in2(_gnd_net_),
            .in3(N__64396),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__86988),
            .ce(N__68767),
            .sr(N__79587));
    defparam \ppm_encoder_1.counter24_0_I_51_c_RNO_LC_16_3_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_51_c_RNO_LC_16_3_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_51_c_RNO_LC_16_3_6 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_51_c_RNO_LC_16_3_6  (
            .in0(N__64332),
            .in1(N__68435),
            .in2(N__64323),
            .in3(N__68480),
            .lcout(\ppm_encoder_1.counter24_0_I_51_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter_0_LC_16_4_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_0_LC_16_4_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_0_LC_16_4_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_0_LC_16_4_0  (
            .in0(_gnd_net_),
            .in1(N__64019),
            .in2(N__64255),
            .in3(N__64172),
            .lcout(\ppm_encoder_1.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_16_4_0_),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_0 ),
            .clk(N__86995),
            .ce(),
            .sr(N__65486));
    defparam \ppm_encoder_1.counter_1_LC_16_4_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_1_LC_16_4_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_1_LC_16_4_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_1_LC_16_4_1  (
            .in0(_gnd_net_),
            .in1(N__63992),
            .in2(_gnd_net_),
            .in3(N__63972),
            .lcout(\ppm_encoder_1.counterZ0Z_1 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_0 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_1 ),
            .clk(N__86995),
            .ce(),
            .sr(N__65486));
    defparam \ppm_encoder_1.counter_2_LC_16_4_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_2_LC_16_4_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_2_LC_16_4_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_2_LC_16_4_2  (
            .in0(_gnd_net_),
            .in1(N__68412),
            .in2(_gnd_net_),
            .in3(N__63969),
            .lcout(\ppm_encoder_1.counterZ0Z_2 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_1 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_2 ),
            .clk(N__86995),
            .ce(),
            .sr(N__65486));
    defparam \ppm_encoder_1.counter_3_LC_16_4_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_3_LC_16_4_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_3_LC_16_4_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_3_LC_16_4_3  (
            .in0(_gnd_net_),
            .in1(N__68457),
            .in2(_gnd_net_),
            .in3(N__64956),
            .lcout(\ppm_encoder_1.counterZ0Z_3 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_2 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_3 ),
            .clk(N__86995),
            .ce(),
            .sr(N__65486));
    defparam \ppm_encoder_1.counter_4_LC_16_4_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_4_LC_16_4_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_4_LC_16_4_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_4_LC_16_4_4  (
            .in0(_gnd_net_),
            .in1(N__64945),
            .in2(_gnd_net_),
            .in3(N__64926),
            .lcout(\ppm_encoder_1.counterZ0Z_4 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_3 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_4 ),
            .clk(N__86995),
            .ce(),
            .sr(N__65486));
    defparam \ppm_encoder_1.counter_5_LC_16_4_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_5_LC_16_4_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_5_LC_16_4_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_5_LC_16_4_5  (
            .in0(_gnd_net_),
            .in1(N__64915),
            .in2(_gnd_net_),
            .in3(N__64896),
            .lcout(\ppm_encoder_1.counterZ0Z_5 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_4 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_5 ),
            .clk(N__86995),
            .ce(),
            .sr(N__65486));
    defparam \ppm_encoder_1.counter_6_LC_16_4_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_6_LC_16_4_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_6_LC_16_4_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_6_LC_16_4_6  (
            .in0(_gnd_net_),
            .in1(N__64882),
            .in2(_gnd_net_),
            .in3(N__64863),
            .lcout(\ppm_encoder_1.counterZ0Z_6 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_5 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_6 ),
            .clk(N__86995),
            .ce(),
            .sr(N__65486));
    defparam \ppm_encoder_1.counter_7_LC_16_4_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_7_LC_16_4_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_7_LC_16_4_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_7_LC_16_4_7  (
            .in0(_gnd_net_),
            .in1(N__64843),
            .in2(_gnd_net_),
            .in3(N__64827),
            .lcout(\ppm_encoder_1.counterZ0Z_7 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_6 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_7 ),
            .clk(N__86995),
            .ce(),
            .sr(N__65486));
    defparam \ppm_encoder_1.counter_8_LC_16_5_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_8_LC_16_5_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_8_LC_16_5_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_8_LC_16_5_0  (
            .in0(_gnd_net_),
            .in1(N__64824),
            .in2(_gnd_net_),
            .in3(N__64806),
            .lcout(\ppm_encoder_1.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_16_5_0_),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_8 ),
            .clk(N__87001),
            .ce(),
            .sr(N__65479));
    defparam \ppm_encoder_1.counter_9_LC_16_5_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_9_LC_16_5_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_9_LC_16_5_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_9_LC_16_5_1  (
            .in0(_gnd_net_),
            .in1(N__64803),
            .in2(_gnd_net_),
            .in3(N__64785),
            .lcout(\ppm_encoder_1.counterZ0Z_9 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_8 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_9 ),
            .clk(N__87001),
            .ce(),
            .sr(N__65479));
    defparam \ppm_encoder_1.counter_10_LC_16_5_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_10_LC_16_5_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_10_LC_16_5_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_10_LC_16_5_2  (
            .in0(_gnd_net_),
            .in1(N__64781),
            .in2(_gnd_net_),
            .in3(N__64761),
            .lcout(\ppm_encoder_1.counterZ0Z_10 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_9 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_10 ),
            .clk(N__87001),
            .ce(),
            .sr(N__65479));
    defparam \ppm_encoder_1.counter_11_LC_16_5_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_11_LC_16_5_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_11_LC_16_5_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_11_LC_16_5_3  (
            .in0(_gnd_net_),
            .in1(N__64757),
            .in2(_gnd_net_),
            .in3(N__65580),
            .lcout(\ppm_encoder_1.counterZ0Z_11 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_10 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_11 ),
            .clk(N__87001),
            .ce(),
            .sr(N__65479));
    defparam \ppm_encoder_1.counter_12_LC_16_5_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_12_LC_16_5_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_12_LC_16_5_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_12_LC_16_5_4  (
            .in0(_gnd_net_),
            .in1(N__65576),
            .in2(_gnd_net_),
            .in3(N__65556),
            .lcout(\ppm_encoder_1.counterZ0Z_12 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_11 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_12 ),
            .clk(N__87001),
            .ce(),
            .sr(N__65479));
    defparam \ppm_encoder_1.counter_13_LC_16_5_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_13_LC_16_5_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_13_LC_16_5_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_13_LC_16_5_5  (
            .in0(_gnd_net_),
            .in1(N__65552),
            .in2(_gnd_net_),
            .in3(N__65532),
            .lcout(\ppm_encoder_1.counterZ0Z_13 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_12 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_13 ),
            .clk(N__87001),
            .ce(),
            .sr(N__65479));
    defparam \ppm_encoder_1.counter_14_LC_16_5_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_14_LC_16_5_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_14_LC_16_5_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_14_LC_16_5_6  (
            .in0(_gnd_net_),
            .in1(N__68556),
            .in2(_gnd_net_),
            .in3(N__65529),
            .lcout(\ppm_encoder_1.counterZ0Z_14 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_13 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_14 ),
            .clk(N__87001),
            .ce(),
            .sr(N__65479));
    defparam \ppm_encoder_1.counter_15_LC_16_5_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_15_LC_16_5_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_15_LC_16_5_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_15_LC_16_5_7  (
            .in0(_gnd_net_),
            .in1(N__68516),
            .in2(_gnd_net_),
            .in3(N__65526),
            .lcout(\ppm_encoder_1.counterZ0Z_15 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_14 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_15 ),
            .clk(N__87001),
            .ce(),
            .sr(N__65479));
    defparam \ppm_encoder_1.counter_16_LC_16_6_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_16_LC_16_6_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_16_LC_16_6_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_16_LC_16_6_0  (
            .in0(_gnd_net_),
            .in1(N__68479),
            .in2(_gnd_net_),
            .in3(N__65523),
            .lcout(\ppm_encoder_1.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_16_6_0_),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_16 ),
            .clk(N__87009),
            .ce(),
            .sr(N__65487));
    defparam \ppm_encoder_1.counter_17_LC_16_6_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_17_LC_16_6_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_17_LC_16_6_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_17_LC_16_6_1  (
            .in0(_gnd_net_),
            .in1(N__68434),
            .in2(_gnd_net_),
            .in3(N__65520),
            .lcout(\ppm_encoder_1.counterZ0Z_17 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_16 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_17 ),
            .clk(N__87009),
            .ce(),
            .sr(N__65487));
    defparam \ppm_encoder_1.counter_18_LC_16_6_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter_18_LC_16_6_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_18_LC_16_6_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ppm_encoder_1.counter_18_LC_16_6_2  (
            .in0(_gnd_net_),
            .in1(N__65510),
            .in2(_gnd_net_),
            .in3(N__65517),
            .lcout(\ppm_encoder_1.counterZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87009),
            .ce(),
            .sr(N__65487));
    defparam \pid_alt.source_data_valid_esr_LC_16_7_0 .C_ON=1'b0;
    defparam \pid_alt.source_data_valid_esr_LC_16_7_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_data_valid_esr_LC_16_7_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.source_data_valid_esr_LC_16_7_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__65436),
            .lcout(pid_altitude_dv),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87016),
            .ce(N__64971),
            .sr(N__79606));
    defparam \pid_side.error_i_acumm_prereg_esr_RNIQL8E1_14_LC_16_8_0 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIQL8E1_14_LC_16_8_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIQL8E1_14_LC_16_8_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_RNIQL8E1_14_LC_16_8_0  (
            .in0(N__65820),
            .in1(N__65714),
            .in2(N__69015),
            .in3(N__65702),
            .lcout(),
            .ltout(\pid_side.un10lto27_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_RNI5LOD5_0_14_LC_16_8_1 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_RNI5LOD5_0_14_LC_16_8_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_acumm_prereg_esr_RNI5LOD5_0_14_LC_16_8_1 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_RNI5LOD5_0_14_LC_16_8_1  (
            .in0(_gnd_net_),
            .in1(N__65625),
            .in2(N__65640),
            .in3(N__65682),
            .lcout(\pid_side.error_i_acumm_prereg_esr_RNI5LOD5_0Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_RNIOLAE1_18_LC_16_8_2 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIOLAE1_18_LC_16_8_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIOLAE1_18_LC_16_8_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_RNIOLAE1_18_LC_16_8_2  (
            .in0(N__65618),
            .in1(N__65606),
            .in2(N__68337),
            .in3(N__65591),
            .lcout(\pid_side.un10lto27_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_18_LC_16_8_3 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_18_LC_16_8_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_18_LC_16_8_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_18_LC_16_8_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70152),
            .lcout(\pid_side.error_i_acumm_preregZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87023),
            .ce(N__69891),
            .sr(N__79612));
    defparam \pid_side.error_i_acumm_prereg_esr_19_LC_16_8_4 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_19_LC_16_8_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_19_LC_16_8_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_19_LC_16_8_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73350),
            .lcout(\pid_side.error_i_acumm_preregZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87023),
            .ce(N__69891),
            .sr(N__79612));
    defparam \pid_side.error_i_acumm_prereg_esr_14_LC_16_8_5 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_14_LC_16_8_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_14_LC_16_8_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_14_LC_16_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82021),
            .lcout(\pid_side.error_i_acumm_preregZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87023),
            .ce(N__69891),
            .sr(N__79612));
    defparam \pid_side.error_i_acumm_prereg_esr_20_LC_16_8_6 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_20_LC_16_8_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_20_LC_16_8_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_20_LC_16_8_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73290),
            .lcout(\pid_side.error_i_acumm_preregZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87023),
            .ce(N__69891),
            .sr(N__79612));
    defparam \pid_side.error_i_acumm_prereg_esr_15_LC_16_8_7 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_15_LC_16_8_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_15_LC_16_8_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_15_LC_16_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78990),
            .lcout(\pid_side.error_i_acumm_preregZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87023),
            .ce(N__69891),
            .sr(N__79612));
    defparam \pid_side.error_i_acumm_prereg_esr_RNIOLAE1_0_18_LC_16_9_0 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIOLAE1_0_18_LC_16_9_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIOLAE1_0_18_LC_16_9_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_RNIOLAE1_0_18_LC_16_9_0  (
            .in0(N__65619),
            .in1(N__65607),
            .in2(N__65595),
            .in3(N__68336),
            .lcout(\pid_side.error_i_acumm16lto27_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_RNITJO21_26_LC_16_9_1 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_RNITJO21_26_LC_16_9_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_acumm_prereg_esr_RNITJO21_26_LC_16_9_1 .LUT_INIT=16'b0000000000000101;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_RNITJO21_26_LC_16_9_1  (
            .in0(N__68318),
            .in1(_gnd_net_),
            .in2(N__65676),
            .in3(N__65775),
            .lcout(\pid_side.error_i_acumm16lto27_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_RNIMLCE1_0_22_LC_16_9_2 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIMLCE1_0_22_LC_16_9_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIMLCE1_0_22_LC_16_9_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_RNIMLCE1_0_22_LC_16_9_2  (
            .in0(N__69036),
            .in1(N__66698),
            .in2(N__69027),
            .in3(N__69045),
            .lcout(),
            .ltout(\pid_side.error_i_acumm16lto27_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_RNI5LOD5_14_LC_16_9_3 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_RNI5LOD5_14_LC_16_9_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_acumm_prereg_esr_RNI5LOD5_14_LC_16_9_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_RNI5LOD5_14_LC_16_9_3  (
            .in0(N__65691),
            .in1(N__65730),
            .in2(N__65724),
            .in3(N__65721),
            .lcout(\pid_side.error_i_acumm16lto27_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_RNIQL8E1_0_14_LC_16_9_4 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIQL8E1_0_14_LC_16_9_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIQL8E1_0_14_LC_16_9_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_RNIQL8E1_0_14_LC_16_9_4  (
            .in0(N__65819),
            .in1(N__65715),
            .in2(N__69014),
            .in3(N__65703),
            .lcout(\pid_side.error_i_acumm16lto27_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_RNIMLCE1_22_LC_16_9_5 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIMLCE1_22_LC_16_9_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIMLCE1_22_LC_16_9_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_RNIMLCE1_22_LC_16_9_5  (
            .in0(N__69044),
            .in1(N__69023),
            .in2(N__66699),
            .in3(N__69035),
            .lcout(),
            .ltout(\pid_side.un10lto27_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_RNIJ95H2_26_LC_16_9_6 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIJ95H2_26_LC_16_9_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIJ95H2_26_LC_16_9_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_RNIJ95H2_26_LC_16_9_6  (
            .in0(N__65774),
            .in1(N__65672),
            .in2(N__65685),
            .in3(N__68317),
            .lcout(\pid_side.un10lto27_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_26_LC_16_9_7 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_26_LC_16_9_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_26_LC_16_9_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_26_LC_16_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__72826),
            .lcout(\pid_side.error_i_acumm_preregZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87033),
            .ce(N__69893),
            .sr(N__79620));
    defparam \pid_side.error_i_acumm_prereg_esr_1_LC_16_10_0 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_1_LC_16_10_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_1_LC_16_10_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_1_LC_16_10_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__72481),
            .lcout(\pid_side.error_i_acumm_preregZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87043),
            .ce(N__69894),
            .sr(N__79627));
    defparam \pid_side.error_i_acumm_prereg_esr_2_LC_16_10_1 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_2_LC_16_10_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_2_LC_16_10_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_2_LC_16_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82162),
            .lcout(\pid_side.error_i_acumm_preregZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87043),
            .ce(N__69894),
            .sr(N__79627));
    defparam \pid_side.error_i_acumm_prereg_esr_3_LC_16_10_2 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_3_LC_16_10_2 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_3_LC_16_10_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_3_LC_16_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81775),
            .lcout(\pid_side.error_i_acumm16lto3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87043),
            .ce(N__69894),
            .sr(N__79627));
    defparam \pid_side.error_i_acumm_prereg_esr_4_LC_16_10_3 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_4_LC_16_10_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_4_LC_16_10_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_4_LC_16_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81483),
            .lcout(\pid_side.error_i_acumm_preregZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87043),
            .ce(N__69894),
            .sr(N__79627));
    defparam \pid_side.error_i_acumm_prereg_esr_16_LC_16_10_4 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_16_LC_16_10_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_16_LC_16_10_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_16_LC_16_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__69792),
            .lcout(\pid_side.error_i_acumm_preregZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87043),
            .ce(N__69894),
            .sr(N__79627));
    defparam \pid_side.error_i_acumm_prereg_esr_6_LC_16_10_5 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_6_LC_16_10_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_6_LC_16_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_6_LC_16_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78538),
            .lcout(\pid_side.error_i_acumm_preregZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87043),
            .ce(N__69894),
            .sr(N__79627));
    defparam \pid_side.error_i_acumm_prereg_esr_9_LC_16_10_6 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_9_LC_16_10_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_9_LC_16_10_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_9_LC_16_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__66424),
            .lcout(\pid_side.error_i_acumm_preregZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87043),
            .ce(N__69894),
            .sr(N__79627));
    defparam \pid_side.error_i_acumm_prereg_esr_27_LC_16_10_7 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_27_LC_16_10_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_27_LC_16_10_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_27_LC_16_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__66843),
            .lcout(\pid_side.error_i_acumm_preregZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87043),
            .ce(N__69894),
            .sr(N__79627));
    defparam \pid_side.error_i_acumm_13_LC_16_11_1 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_13_LC_16_11_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_13_LC_16_11_1 .LUT_INIT=16'b1110101001000000;
    LogicCell40 \pid_side.error_i_acumm_13_LC_16_11_1  (
            .in0(N__65880),
            .in1(N__65924),
            .in2(N__72655),
            .in3(N__68322),
            .lcout(\pid_side.error_i_acummZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87052),
            .ce(N__66108),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_11_LC_16_11_2 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_11_LC_16_11_2 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_11_LC_16_11_2 .LUT_INIT=16'b1111000010001000;
    LogicCell40 \pid_side.error_i_acumm_11_LC_16_11_2  (
            .in0(N__65923),
            .in1(N__72643),
            .in2(N__65766),
            .in3(N__65879),
            .lcout(\pid_side.error_i_acummZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87052),
            .ce(N__66108),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_4_LC_16_11_3 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_4_LC_16_11_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_4_LC_16_11_3 .LUT_INIT=16'b1110101001000000;
    LogicCell40 \pid_side.error_i_acumm_4_LC_16_11_3  (
            .in0(N__65881),
            .in1(N__65925),
            .in2(N__72656),
            .in3(N__65745),
            .lcout(\pid_side.error_i_acummZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87052),
            .ce(N__66108),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_5_LC_16_11_4 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_5_LC_16_11_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_5_LC_16_11_4 .LUT_INIT=16'b1111000010001000;
    LogicCell40 \pid_side.error_i_acumm_5_LC_16_11_4  (
            .in0(N__65926),
            .in1(N__72644),
            .in2(N__68994),
            .in3(N__65882),
            .lcout(\pid_side.error_i_acummZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87052),
            .ce(N__66108),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_6_LC_16_11_5 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_6_LC_16_11_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_6_LC_16_11_5 .LUT_INIT=16'b1110101001000000;
    LogicCell40 \pid_side.error_i_acumm_6_LC_16_11_5  (
            .in0(N__65883),
            .in1(N__65927),
            .in2(N__72657),
            .in3(N__66124),
            .lcout(\pid_side.error_i_acummZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87052),
            .ce(N__66108),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_RNIF9KEA_28_LC_16_11_6 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIF9KEA_28_LC_16_11_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIF9KEA_28_LC_16_11_6 .LUT_INIT=16'b0000000011110010;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_RNIF9KEA_28_LC_16_11_6  (
            .in0(N__66063),
            .in1(N__66054),
            .in2(N__72548),
            .in3(N__65994),
            .lcout(\pid_side.error_i_acumm_2_sqmuxa_1 ),
            .ltout(\pid_side.error_i_acumm_2_sqmuxa_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_RNIQVDQK_28_LC_16_11_7 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIQVDQK_28_LC_16_11_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIQVDQK_28_LC_16_11_7 .LUT_INIT=16'b0010000010100000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_RNIQVDQK_28_LC_16_11_7  (
            .in0(N__72642),
            .in1(N__72544),
            .in2(N__65904),
            .in3(N__65901),
            .lcout(\pid_side.error_i_acumm_2_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI2HLL1_22_LC_16_12_0 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI2HLL1_22_LC_16_12_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI2HLL1_22_LC_16_12_0 .LUT_INIT=16'b1110111100001000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI2HLL1_22_LC_16_12_0  (
            .in0(N__83566),
            .in1(N__84623),
            .in2(N__73207),
            .in3(N__66722),
            .lcout(\pid_side.un1_pid_prereg_0_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI1QLO_22_LC_16_12_1 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI1QLO_22_LC_16_12_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI1QLO_22_LC_16_12_1 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI1QLO_22_LC_16_12_1  (
            .in0(N__84621),
            .in1(N__73182),
            .in2(_gnd_net_),
            .in3(N__83562),
            .lcout(\pid_side.un1_pid_prereg_370_1 ),
            .ltout(\pid_side.un1_pid_prereg_370_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIMN4E2_21_LC_16_12_2 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIMN4E2_21_LC_16_12_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIMN4E2_21_LC_16_12_2 .LUT_INIT=16'b1111110011000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIMN4E2_21_LC_16_12_2  (
            .in0(_gnd_net_),
            .in1(N__73104),
            .in2(N__65838),
            .in3(N__69836),
            .lcout(\pid_side.un1_pid_prereg_0_14 ),
            .ltout(\pid_side.un1_pid_prereg_0_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIK1TV8_22_LC_16_12_3 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIK1TV8_22_LC_16_12_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIK1TV8_22_LC_16_12_3 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIK1TV8_22_LC_16_12_3  (
            .in0(N__73419),
            .in1(N__73440),
            .in2(N__65835),
            .in3(N__68939),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIK1TV8Z0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIP2GL1_0_22_LC_16_12_4 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIP2GL1_0_22_LC_16_12_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIP2GL1_0_22_LC_16_12_4 .LUT_INIT=16'b0110010101011001;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIP2GL1_0_22_LC_16_12_4  (
            .in0(N__69236),
            .in1(N__73186),
            .in2(N__83573),
            .in3(N__84622),
            .lcout(\pid_side.un1_pid_prereg_0_15 ),
            .ltout(\pid_side.un1_pid_prereg_0_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIFQK34_22_LC_16_12_5 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIFQK34_22_LC_16_12_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIFQK34_22_LC_16_12_5 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIFQK34_22_LC_16_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__65832),
            .in3(N__68960),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIFQK34Z0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_esr_RNO_0_30_LC_16_12_6 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_esr_RNO_0_30_LC_16_12_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_esr_RNO_0_30_LC_16_12_6 .LUT_INIT=16'b1000011101111000;
    LogicCell40 \pid_side.pid_prereg_esr_RNO_0_30_LC_16_12_6  (
            .in0(N__66307),
            .in1(N__66290),
            .in2(N__66312),
            .in3(N__66291),
            .lcout(\pid_side.un1_pid_prereg_0_axb_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI72LM6_22_LC_16_12_7 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI72LM6_22_LC_16_12_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI72LM6_22_LC_16_12_7 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI72LM6_22_LC_16_12_7  (
            .in0(N__66327),
            .in1(N__66289),
            .in2(N__66311),
            .in3(N__66288),
            .lcout(\pid_side.error_d_reg_prev_esr_RNI72LM6Z0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNIARAI_0_LC_16_13_0 .C_ON=1'b1;
    defparam \pid_side.error_i_reg_esr_RNIARAI_0_LC_16_13_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNIARAI_0_LC_16_13_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \pid_side.error_i_reg_esr_RNIARAI_0_LC_16_13_0  (
            .in0(_gnd_net_),
            .in1(N__66254),
            .in2(N__66239),
            .in3(_gnd_net_),
            .lcout(\pid_side.un1_pid_prereg_0 ),
            .ltout(),
            .carryin(bfn_16_13_0_),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_0_c_RNITGKN_LC_16_13_1 .C_ON=1'b1;
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_0_c_RNITGKN_LC_16_13_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_0_c_RNITGKN_LC_16_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_0_c_RNITGKN_LC_16_13_1  (
            .in0(_gnd_net_),
            .in1(N__66222),
            .in2(N__66213),
            .in3(N__66201),
            .lcout(\pid_side.un1_error_i_acumm_prereg_cry_0_c_RNITGKN ),
            .ltout(),
            .carryin(\pid_side.un1_error_i_acumm_prereg_cry_0 ),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_1_c_RNI0LLN_LC_16_13_2 .C_ON=1'b1;
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_1_c_RNI0LLN_LC_16_13_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_1_c_RNI0LLN_LC_16_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_1_c_RNI0LLN_LC_16_13_2  (
            .in0(_gnd_net_),
            .in1(N__66198),
            .in2(N__66189),
            .in3(N__66180),
            .lcout(\pid_side.un1_error_i_acumm_prereg_cry_1_c_RNI0LLN ),
            .ltout(),
            .carryin(\pid_side.un1_error_i_acumm_prereg_cry_1 ),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_2_c_RNI3PMN_LC_16_13_3 .C_ON=1'b1;
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_2_c_RNI3PMN_LC_16_13_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_2_c_RNI3PMN_LC_16_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_2_c_RNI3PMN_LC_16_13_3  (
            .in0(_gnd_net_),
            .in1(N__66177),
            .in2(N__66168),
            .in3(N__66156),
            .lcout(\pid_side.un1_error_i_acumm_prereg_cry_2_c_RNI3PMN ),
            .ltout(),
            .carryin(\pid_side.un1_error_i_acumm_prereg_cry_2 ),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_3_c_RNI6TNN_LC_16_13_4 .C_ON=1'b1;
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_3_c_RNI6TNN_LC_16_13_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_3_c_RNI6TNN_LC_16_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_3_c_RNI6TNN_LC_16_13_4  (
            .in0(_gnd_net_),
            .in1(N__66153),
            .in2(N__66960),
            .in3(N__66144),
            .lcout(\pid_side.un1_error_i_acumm_prereg_cry_3_c_RNI6TNN ),
            .ltout(),
            .carryin(\pid_side.un1_error_i_acumm_prereg_cry_3 ),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_4_c_RNI91PN_LC_16_13_5 .C_ON=1'b1;
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_4_c_RNI91PN_LC_16_13_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_4_c_RNI91PN_LC_16_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_4_c_RNI91PN_LC_16_13_5  (
            .in0(_gnd_net_),
            .in1(N__66141),
            .in2(N__75390),
            .in3(N__66132),
            .lcout(\pid_side.un1_error_i_acumm_prereg_cry_4_c_RNI91PN ),
            .ltout(),
            .carryin(\pid_side.un1_error_i_acumm_prereg_cry_4 ),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_5_c_RNIC5QN_LC_16_13_6 .C_ON=1'b1;
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_5_c_RNIC5QN_LC_16_13_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_5_c_RNIC5QN_LC_16_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_5_c_RNIC5QN_LC_16_13_6  (
            .in0(_gnd_net_),
            .in1(N__66552),
            .in2(N__66543),
            .in3(N__66531),
            .lcout(\pid_side.un1_error_i_acumm_prereg_cry_5_c_RNIC5QN ),
            .ltout(),
            .carryin(\pid_side.un1_error_i_acumm_prereg_cry_5 ),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_6_c_RNIF9RN_LC_16_13_7 .C_ON=1'b1;
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_6_c_RNIF9RN_LC_16_13_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_6_c_RNIF9RN_LC_16_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_6_c_RNIF9RN_LC_16_13_7  (
            .in0(_gnd_net_),
            .in1(N__66528),
            .in2(N__66522),
            .in3(N__66480),
            .lcout(\pid_side.un1_error_i_acumm_prereg_cry_6_c_RNIF9RN ),
            .ltout(),
            .carryin(\pid_side.un1_error_i_acumm_prereg_cry_6 ),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_7_c_RNI9JMJ_LC_16_14_0 .C_ON=1'b1;
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_7_c_RNI9JMJ_LC_16_14_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_7_c_RNI9JMJ_LC_16_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_7_c_RNI9JMJ_LC_16_14_0  (
            .in0(_gnd_net_),
            .in1(N__66477),
            .in2(N__66930),
            .in3(N__66438),
            .lcout(\pid_side.un1_error_i_acumm_prereg_cry_7_c_RNI9JMJ ),
            .ltout(),
            .carryin(bfn_16_14_0_),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_8_c_RNILHTN_LC_16_14_1 .C_ON=1'b1;
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_8_c_RNILHTN_LC_16_14_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_8_c_RNILHTN_LC_16_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_8_c_RNILHTN_LC_16_14_1  (
            .in0(_gnd_net_),
            .in1(N__66435),
            .in2(N__66987),
            .in3(N__66402),
            .lcout(\pid_side.un1_error_i_acumm_prereg_cry_8_c_RNILHTN ),
            .ltout(),
            .carryin(\pid_side.un1_error_i_acumm_prereg_cry_8 ),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNI6OOI_10_LC_16_14_2 .C_ON=1'b1;
    defparam \pid_side.error_i_reg_esr_RNI6OOI_10_LC_16_14_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNI6OOI_10_LC_16_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_i_reg_esr_RNI6OOI_10_LC_16_14_2  (
            .in0(_gnd_net_),
            .in1(N__66399),
            .in2(N__66387),
            .in3(N__66375),
            .lcout(\pid_side.error_i_reg_esr_RNI6OOIZ0Z_10 ),
            .ltout(),
            .carryin(\pid_side.un1_error_i_acumm_prereg_cry_9 ),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNIGRJR_11_LC_16_14_3 .C_ON=1'b1;
    defparam \pid_side.error_i_reg_esr_RNIGRJR_11_LC_16_14_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNIGRJR_11_LC_16_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_i_reg_esr_RNIGRJR_11_LC_16_14_3  (
            .in0(_gnd_net_),
            .in1(N__66372),
            .in2(N__66363),
            .in3(N__66348),
            .lcout(\pid_side.error_i_reg_esr_RNIGRJRZ0Z_11 ),
            .ltout(),
            .carryin(\pid_side.un1_error_i_acumm_prereg_cry_10 ),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNIJVKR_12_LC_16_14_4 .C_ON=1'b1;
    defparam \pid_side.error_i_reg_esr_RNIJVKR_12_LC_16_14_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNIJVKR_12_LC_16_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_i_reg_esr_RNIJVKR_12_LC_16_14_4  (
            .in0(_gnd_net_),
            .in1(N__66345),
            .in2(N__67872),
            .in3(N__66333),
            .lcout(\pid_side.error_i_reg_esr_RNIJVKRZ0Z_12 ),
            .ltout(),
            .carryin(\pid_side.un1_error_i_acumm_prereg_cry_11 ),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNIM3MR_13_LC_16_14_5 .C_ON=1'b1;
    defparam \pid_side.error_i_reg_esr_RNIM3MR_13_LC_16_14_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNIM3MR_13_LC_16_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_i_reg_esr_RNIM3MR_13_LC_16_14_5  (
            .in0(_gnd_net_),
            .in1(N__66771),
            .in2(N__70725),
            .in3(N__66330),
            .lcout(\pid_side.error_i_reg_esr_RNIM3MRZ0Z_13 ),
            .ltout(),
            .carryin(\pid_side.un1_error_i_acumm_prereg_cry_12 ),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNIO6NR_14_LC_16_14_6 .C_ON=1'b1;
    defparam \pid_side.error_i_reg_esr_RNIO6NR_14_LC_16_14_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNIO6NR_14_LC_16_14_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_i_reg_esr_RNIO6NR_14_LC_16_14_6  (
            .in0(_gnd_net_),
            .in1(N__66681),
            .in2(N__66801),
            .in3(N__66669),
            .lcout(\pid_side.error_i_reg_esr_RNIO6NRZ0Z_14 ),
            .ltout(),
            .carryin(\pid_side.un1_error_i_acumm_prereg_cry_13 ),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNIQ9OR_15_LC_16_14_7 .C_ON=1'b1;
    defparam \pid_side.error_i_reg_esr_RNIQ9OR_15_LC_16_14_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNIQ9OR_15_LC_16_14_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_i_reg_esr_RNIQ9OR_15_LC_16_14_7  (
            .in0(_gnd_net_),
            .in1(N__66775),
            .in2(N__66666),
            .in3(N__66651),
            .lcout(\pid_side.error_i_reg_esr_RNIQ9ORZ0Z_15 ),
            .ltout(),
            .carryin(\pid_side.un1_error_i_acumm_prereg_cry_14 ),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNISCPR_16_LC_16_15_0 .C_ON=1'b1;
    defparam \pid_side.error_i_reg_esr_RNISCPR_16_LC_16_15_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNISCPR_16_LC_16_15_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_i_reg_esr_RNISCPR_16_LC_16_15_0  (
            .in0(_gnd_net_),
            .in1(N__66776),
            .in2(N__66648),
            .in3(N__66636),
            .lcout(\pid_side.error_i_reg_esr_RNISCPRZ0Z_16 ),
            .ltout(),
            .carryin(bfn_16_15_0_),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNIUFQR_17_LC_16_15_1 .C_ON=1'b1;
    defparam \pid_side.error_i_reg_esr_RNIUFQR_17_LC_16_15_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNIUFQR_17_LC_16_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_i_reg_esr_RNIUFQR_17_LC_16_15_1  (
            .in0(_gnd_net_),
            .in1(N__67461),
            .in2(N__66802),
            .in3(N__66633),
            .lcout(\pid_side.error_i_reg_esr_RNIUFQRZ0Z_17 ),
            .ltout(),
            .carryin(\pid_side.un1_error_i_acumm_prereg_cry_16 ),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNI0JRR_18_LC_16_15_2 .C_ON=1'b1;
    defparam \pid_side.error_i_reg_esr_RNI0JRR_18_LC_16_15_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNI0JRR_18_LC_16_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_i_reg_esr_RNI0JRR_18_LC_16_15_2  (
            .in0(_gnd_net_),
            .in1(N__66780),
            .in2(N__66630),
            .in3(N__66618),
            .lcout(\pid_side.error_i_reg_esr_RNI0JRRZ0Z_18 ),
            .ltout(),
            .carryin(\pid_side.un1_error_i_acumm_prereg_cry_17 ),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNI2MSR_19_LC_16_15_3 .C_ON=1'b1;
    defparam \pid_side.error_i_reg_esr_RNI2MSR_19_LC_16_15_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNI2MSR_19_LC_16_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_i_reg_esr_RNI2MSR_19_LC_16_15_3  (
            .in0(_gnd_net_),
            .in1(N__66615),
            .in2(N__66803),
            .in3(N__66603),
            .lcout(\pid_side.error_i_reg_esr_RNI2MSRZ0Z_19 ),
            .ltout(),
            .carryin(\pid_side.un1_error_i_acumm_prereg_cry_18 ),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNIRGUR_20_LC_16_15_4 .C_ON=1'b1;
    defparam \pid_side.error_i_reg_esr_RNIRGUR_20_LC_16_15_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNIRGUR_20_LC_16_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_i_reg_esr_RNIRGUR_20_LC_16_15_4  (
            .in0(_gnd_net_),
            .in1(N__66784),
            .in2(N__66600),
            .in3(N__66585),
            .lcout(\pid_side.error_i_reg_esr_RNIRGURZ0Z_20 ),
            .ltout(),
            .carryin(\pid_side.un1_error_i_acumm_prereg_cry_19 ),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNIK2OS_21_LC_16_15_5 .C_ON=1'b1;
    defparam \pid_side.error_i_reg_esr_RNIK2OS_21_LC_16_15_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNIK2OS_21_LC_16_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_i_reg_esr_RNIK2OS_21_LC_16_15_5  (
            .in0(_gnd_net_),
            .in1(N__66582),
            .in2(N__66804),
            .in3(N__66570),
            .lcout(\pid_side.error_i_reg_esr_RNIK2OSZ0Z_21 ),
            .ltout(),
            .carryin(\pid_side.un1_error_i_acumm_prereg_cry_20 ),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNIM5PS_22_LC_16_15_6 .C_ON=1'b1;
    defparam \pid_side.error_i_reg_esr_RNIM5PS_22_LC_16_15_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNIM5PS_22_LC_16_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_i_reg_esr_RNIM5PS_22_LC_16_15_6  (
            .in0(_gnd_net_),
            .in1(N__66788),
            .in2(N__66567),
            .in3(N__66879),
            .lcout(\pid_side.error_i_reg_esr_RNIM5PSZ0Z_22 ),
            .ltout(),
            .carryin(\pid_side.un1_error_i_acumm_prereg_cry_21 ),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNIO8QS_23_LC_16_15_7 .C_ON=1'b1;
    defparam \pid_side.error_i_reg_esr_RNIO8QS_23_LC_16_15_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNIO8QS_23_LC_16_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_i_reg_esr_RNIO8QS_23_LC_16_15_7  (
            .in0(_gnd_net_),
            .in1(N__66876),
            .in2(N__66805),
            .in3(N__66870),
            .lcout(\pid_side.error_i_reg_esr_RNIO8QSZ0Z_23 ),
            .ltout(),
            .carryin(\pid_side.un1_error_i_acumm_prereg_cry_22 ),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNIQBRS_24_LC_16_16_0 .C_ON=1'b1;
    defparam \pid_side.error_i_reg_esr_RNIQBRS_24_LC_16_16_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNIQBRS_24_LC_16_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_i_reg_esr_RNIQBRS_24_LC_16_16_0  (
            .in0(_gnd_net_),
            .in1(N__66792),
            .in2(N__70215),
            .in3(N__66867),
            .lcout(\pid_side.error_i_reg_esr_RNIQBRSZ0Z_24 ),
            .ltout(),
            .carryin(bfn_16_16_0_),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNISESS_25_LC_16_16_1 .C_ON=1'b1;
    defparam \pid_side.error_i_reg_esr_RNISESS_25_LC_16_16_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNISESS_25_LC_16_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_i_reg_esr_RNISESS_25_LC_16_16_1  (
            .in0(_gnd_net_),
            .in1(N__67446),
            .in2(N__66806),
            .in3(N__66864),
            .lcout(\pid_side.error_i_reg_esr_RNISESSZ0Z_25 ),
            .ltout(),
            .carryin(\pid_side.un1_error_i_acumm_prereg_cry_24 ),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNIUHTS_26_LC_16_16_2 .C_ON=1'b1;
    defparam \pid_side.error_i_reg_esr_RNIUHTS_26_LC_16_16_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNIUHTS_26_LC_16_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_i_reg_esr_RNIUHTS_26_LC_16_16_2  (
            .in0(_gnd_net_),
            .in1(N__66796),
            .in2(N__66861),
            .in3(N__66846),
            .lcout(\pid_side.error_i_reg_esr_RNIUHTSZ0Z_26 ),
            .ltout(),
            .carryin(\pid_side.un1_error_i_acumm_prereg_cry_25 ),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_26_c_RNI0LUS_LC_16_16_3 .C_ON=1'b1;
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_26_c_RNI0LUS_LC_16_16_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_26_c_RNI0LUS_LC_16_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_26_c_RNI0LUS_LC_16_16_3  (
            .in0(_gnd_net_),
            .in1(N__66818),
            .in2(N__66807),
            .in3(N__66822),
            .lcout(\pid_side.un1_error_i_acumm_prereg_cry_26_c_RNI0LUS ),
            .ltout(),
            .carryin(\pid_side.un1_error_i_acumm_prereg_cry_26 ),
            .carryout(\pid_side.un1_error_i_acumm_prereg_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_27_c_RNI1NVS_LC_16_16_4 .C_ON=1'b0;
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_27_c_RNI1NVS_LC_16_16_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_27_c_RNI1NVS_LC_16_16_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_side.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_27_c_RNI1NVS_LC_16_16_4  (
            .in0(N__66819),
            .in1(N__66800),
            .in2(_gnd_net_),
            .in3(N__66726),
            .lcout(\pid_side.un1_error_i_acumm_prereg_cry_27_c_RNI1NVS ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_28_LC_16_16_5 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_28_LC_16_16_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_28_LC_16_16_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_28_LC_16_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__66721),
            .lcout(\pid_side.error_i_acumm_preregZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87111),
            .ce(N__69900),
            .sr(N__79675));
    defparam \pid_side.error_i_acumm_prereg_esr_25_LC_16_16_7 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_25_LC_16_16_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_25_LC_16_16_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_25_LC_16_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__72892),
            .lcout(\pid_side.error_i_acumm_preregZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87111),
            .ce(N__69900),
            .sr(N__79675));
    defparam \pid_side.error_cry_0_c_RNIOJ1L2_LC_16_17_0 .C_ON=1'b0;
    defparam \pid_side.error_cry_0_c_RNIOJ1L2_LC_16_17_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_0_c_RNIOJ1L2_LC_16_17_0 .LUT_INIT=16'b0111001101000011;
    LogicCell40 \pid_side.error_cry_0_c_RNIOJ1L2_LC_16_17_0  (
            .in0(N__80213),
            .in1(N__77799),
            .in2(N__80395),
            .in3(N__67115),
            .lcout(),
            .ltout(\pid_side.m32_0_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_7_c_RNIKG31E_LC_16_17_1 .C_ON=1'b0;
    defparam \pid_side.error_cry_7_c_RNIKG31E_LC_16_17_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_7_c_RNIKG31E_LC_16_17_1 .LUT_INIT=16'b0000110100111101;
    LogicCell40 \pid_side.error_cry_7_c_RNIKG31E_LC_16_17_1  (
            .in0(N__67067),
            .in1(N__76270),
            .in2(N__66948),
            .in3(N__66909),
            .lcout(\pid_side.N_89_i ),
            .ltout(\pid_side.N_89_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_8_LC_16_17_2 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_8_LC_16_17_2 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_8_LC_16_17_2 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \pid_side.error_i_reg_8_LC_16_17_2  (
            .in0(N__66926),
            .in1(N__75474),
            .in2(N__66945),
            .in3(N__66942),
            .lcout(\pid_side.error_i_regZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87124),
            .ce(),
            .sr(N__79680));
    defparam \pid_side.error_cry_7_c_RNIDB5S4_LC_16_17_3 .C_ON=1'b0;
    defparam \pid_side.error_cry_7_c_RNIDB5S4_LC_16_17_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_7_c_RNIDB5S4_LC_16_17_3 .LUT_INIT=16'b1111010100000011;
    LogicCell40 \pid_side.error_cry_7_c_RNIDB5S4_LC_16_17_3  (
            .in0(N__74063),
            .in1(N__74181),
            .in2(N__80972),
            .in3(N__70260),
            .lcout(\pid_side.N_22_0 ),
            .ltout(\pid_side.N_22_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_3_16_LC_16_17_4 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_3_16_LC_16_17_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_3_16_LC_16_17_4 .LUT_INIT=16'b1100100001000000;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_3_16_LC_16_17_4  (
            .in0(N__80533),
            .in1(N__75690),
            .in2(N__66912),
            .in3(N__67065),
            .lcout(\pid_side.error_i_reg_esr_RNO_3Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_4_16_LC_16_17_5 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_4_16_LC_16_17_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_4_16_LC_16_17_5 .LUT_INIT=16'b1011111110001111;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_4_16_LC_16_17_5  (
            .in0(N__67066),
            .in1(N__80534),
            .in2(N__75739),
            .in3(N__66908),
            .lcout(),
            .ltout(\pid_side.error_i_reg_esr_RNO_4Z0Z_16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_1_16_LC_16_17_6 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_1_16_LC_16_17_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_1_16_LC_16_17_6 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_1_16_LC_16_17_6  (
            .in0(_gnd_net_),
            .in1(N__70239),
            .in2(N__66900),
            .in3(N__66897),
            .lcout(\pid_side.m20_2_03_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_3_17_LC_16_18_0 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_3_17_LC_16_18_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_3_17_LC_16_18_0 .LUT_INIT=16'b0010000000100011;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_3_17_LC_16_18_0  (
            .in0(N__71016),
            .in1(N__76269),
            .in2(N__71551),
            .in3(N__70869),
            .lcout(\pid_front.m5_2_03 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNI08RD_13_LC_16_18_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNI08RD_13_LC_16_18_1 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNI08RD_13_LC_16_18_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_RNI08RD_13_LC_16_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73973),
            .lcout(drone_H_disp_side_i_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_3_c_RNI6SLI2_LC_16_18_2 .C_ON=1'b0;
    defparam \pid_side.error_cry_3_c_RNI6SLI2_LC_16_18_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_3_c_RNI6SLI2_LC_16_18_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \pid_side.error_cry_3_c_RNI6SLI2_LC_16_18_2  (
            .in0(N__80959),
            .in1(N__67047),
            .in2(_gnd_net_),
            .in3(N__70289),
            .lcout(\pid_side.N_12_1 ),
            .ltout(\pid_side.N_12_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_0_c_RNI30FD3_LC_16_18_3 .C_ON=1'b0;
    defparam \pid_side.error_cry_0_c_RNI30FD3_LC_16_18_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_0_c_RNI30FD3_LC_16_18_3 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \pid_side.error_cry_0_c_RNI30FD3_LC_16_18_3  (
            .in0(N__80594),
            .in1(_gnd_net_),
            .in2(N__67008),
            .in3(N__70580),
            .lcout(\pid_side.N_93_0 ),
            .ltout(\pid_side.N_93_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_0_25_LC_16_18_4 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_0_25_LC_16_18_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_0_25_LC_16_18_4 .LUT_INIT=16'b1100010010000000;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_0_25_LC_16_18_4  (
            .in0(N__76840),
            .in1(N__76514),
            .in2(N__67005),
            .in3(N__66999),
            .lcout(\pid_side.error_i_reg_9_rn_1_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_3_25_LC_16_18_6 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_3_25_LC_16_18_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_3_25_LC_16_18_6 .LUT_INIT=16'b0101111111111111;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_3_25_LC_16_18_6  (
            .in0(N__80960),
            .in1(_gnd_net_),
            .in2(N__71550),
            .in3(N__80767),
            .lcout(),
            .ltout(\pid_side.un4_error_i_reg_35_am_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_2_25_LC_16_18_7 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_2_25_LC_16_18_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_2_25_LC_16_18_7 .LUT_INIT=16'b1111110100001000;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_2_25_LC_16_18_7  (
            .in0(N__75742),
            .in1(N__74404),
            .in2(N__67002),
            .in3(N__74868),
            .lcout(\pid_side.error_i_reg_esr_RNO_2_0_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_9_LC_16_19_0 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_9_LC_16_19_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_esr_9_LC_16_19_0 .LUT_INIT=16'b1000000011010000;
    LogicCell40 \pid_side.error_i_reg_esr_9_LC_16_19_0  (
            .in0(N__75738),
            .in1(N__66993),
            .in2(N__75481),
            .in3(N__70272),
            .lcout(\pid_side.error_i_regZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87157),
            .ce(N__75332),
            .sr(N__79688));
    defparam \pid_side.m101_e_LC_16_19_1 .C_ON=1'b0;
    defparam \pid_side.m101_e_LC_16_19_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.m101_e_LC_16_19_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_side.m101_e_LC_16_19_1  (
            .in0(N__70634),
            .in1(N__70710),
            .in2(N__70680),
            .in3(N__76913),
            .lcout(pid_side_N_166),
            .ltout(pid_side_N_166_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_4_LC_16_19_2 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_4_LC_16_19_2 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_esr_4_LC_16_19_2 .LUT_INIT=16'b1101000010000000;
    LogicCell40 \pid_side.error_i_reg_esr_4_LC_16_19_2  (
            .in0(N__76272),
            .in1(N__67430),
            .in2(N__66972),
            .in3(N__66969),
            .lcout(\pid_side.error_i_regZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87157),
            .ce(N__75332),
            .sr(N__79688));
    defparam \pid_front.m64_e_LC_16_19_3 .C_ON=1'b0;
    defparam \pid_front.m64_e_LC_16_19_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.m64_e_LC_16_19_3 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \pid_front.m64_e_LC_16_19_3  (
            .in0(N__70633),
            .in1(N__70709),
            .in2(_gnd_net_),
            .in3(N__70676),
            .lcout(pid_front_N_331),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_17_LC_16_19_4 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_17_LC_16_19_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_esr_17_LC_16_19_4 .LUT_INIT=16'b0111011100100010;
    LogicCell40 \pid_side.error_i_reg_esr_17_LC_16_19_4  (
            .in0(N__68202),
            .in1(N__70270),
            .in2(_gnd_net_),
            .in3(N__67467),
            .lcout(\pid_side.error_i_regZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87157),
            .ce(N__75332),
            .sr(N__79688));
    defparam \pid_side.error_i_reg_esr_25_LC_16_19_5 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_25_LC_16_19_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_esr_25_LC_16_19_5 .LUT_INIT=16'b0111011101000100;
    LogicCell40 \pid_side.error_i_reg_esr_25_LC_16_19_5  (
            .in0(N__70271),
            .in1(N__68190),
            .in2(_gnd_net_),
            .in3(N__67452),
            .lcout(\pid_side.error_i_regZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87157),
            .ce(N__75332),
            .sr(N__79688));
    defparam \pid_side.m61_0_bm_LC_16_19_6 .C_ON=1'b0;
    defparam \pid_side.m61_0_bm_LC_16_19_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.m61_0_bm_LC_16_19_6 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \pid_side.m61_0_bm_LC_16_19_6  (
            .in0(N__81058),
            .in1(N__80609),
            .in2(N__72057),
            .in3(N__80792),
            .lcout(\pid_side.m61_0_bmZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_5_c_RNIJV481_LC_16_20_0 .C_ON=1'b0;
    defparam \pid_front.error_cry_5_c_RNIJV481_LC_16_20_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_5_c_RNIJV481_LC_16_20_0 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \pid_front.error_cry_5_c_RNIJV481_LC_16_20_0  (
            .in0(N__78244),
            .in1(N__67320),
            .in2(_gnd_net_),
            .in3(N__67404),
            .lcout(\pid_front.N_47_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_5_13_LC_16_20_1 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_5_13_LC_16_20_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_5_13_LC_16_20_1 .LUT_INIT=16'b0000110001110111;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_5_13_LC_16_20_1  (
            .in0(N__67405),
            .in1(N__72036),
            .in2(N__67330),
            .in3(N__78380),
            .lcout(),
            .ltout(\pid_front.g0_15_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_2_13_LC_16_20_2 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_2_13_LC_16_20_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_2_13_LC_16_20_2 .LUT_INIT=16'b1011000010110101;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_2_13_LC_16_20_2  (
            .in0(N__72037),
            .in1(N__67237),
            .in2(N__67194),
            .in3(N__67183),
            .lcout(\pid_front.N_88_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_0_12_LC_16_20_3 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_0_12_LC_16_20_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_0_12_LC_16_20_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_0_12_LC_16_20_3  (
            .in0(N__72044),
            .in1(N__70251),
            .in2(_gnd_net_),
            .in3(N__67122),
            .lcout(\pid_side.N_129 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_4_12_LC_16_20_4 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_4_12_LC_16_20_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_4_12_LC_16_20_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_4_12_LC_16_20_4  (
            .in0(N__80613),
            .in1(N__67116),
            .in2(_gnd_net_),
            .in3(N__67071),
            .lcout(),
            .ltout(\pid_side.N_60_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_1_12_LC_16_20_5 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_1_12_LC_16_20_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_1_12_LC_16_20_5 .LUT_INIT=16'b1000101100000000;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_1_12_LC_16_20_5  (
            .in0(N__80190),
            .in1(N__77005),
            .in2(N__67050),
            .in3(N__76535),
            .lcout(),
            .ltout(\pid_side.error_i_reg_9_rn_1_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_12_LC_16_20_6 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_12_LC_16_20_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_esr_12_LC_16_20_6 .LUT_INIT=16'b0101000011111010;
    LogicCell40 \pid_side.error_i_reg_esr_12_LC_16_20_6  (
            .in0(N__70903),
            .in1(_gnd_net_),
            .in2(N__67881),
            .in3(N__67878),
            .lcout(\pid_side.error_i_regZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87171),
            .ce(N__75344),
            .sr(N__79690));
    defparam \pid_front.error_cry_1_0_c_RNIDPRQ1_LC_16_21_0 .C_ON=1'b0;
    defparam \pid_front.error_cry_1_0_c_RNIDPRQ1_LC_16_21_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_1_0_c_RNIDPRQ1_LC_16_21_0 .LUT_INIT=16'b1010111010111111;
    LogicCell40 \pid_front.error_cry_1_0_c_RNIDPRQ1_LC_16_21_0  (
            .in0(N__78045),
            .in1(N__78215),
            .in2(N__67746),
            .in3(N__67667),
            .lcout(\pid_front.error_cry_1_0_c_RNIDPRQZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_0_0_c_RNIJE041_LC_16_21_1 .C_ON=1'b0;
    defparam \pid_front.error_cry_0_0_c_RNIJE041_LC_16_21_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_0_0_c_RNIJE041_LC_16_21_1 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \pid_front.error_cry_0_0_c_RNIJE041_LC_16_21_1  (
            .in0(N__78214),
            .in1(N__67845),
            .in2(_gnd_net_),
            .in3(N__67788),
            .lcout(\pid_front.N_9_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_1_0_c_RNIDPRQ1_0_LC_16_21_2 .C_ON=1'b0;
    defparam \pid_front.error_cry_1_0_c_RNIDPRQ1_0_LC_16_21_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_1_0_c_RNIDPRQ1_0_LC_16_21_2 .LUT_INIT=16'b0000010000010101;
    LogicCell40 \pid_front.error_cry_1_0_c_RNIDPRQ1_0_LC_16_21_2  (
            .in0(N__78046),
            .in1(N__78216),
            .in2(N__67747),
            .in3(N__67668),
            .lcout(),
            .ltout(\pid_front.error_cry_1_0_c_RNIDPRQ1Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_0_0_c_RNID1OP4_LC_16_21_3 .C_ON=1'b0;
    defparam \pid_front.error_cry_0_0_c_RNID1OP4_LC_16_21_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_0_0_c_RNID1OP4_LC_16_21_3 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \pid_front.error_cry_0_0_c_RNID1OP4_LC_16_21_3  (
            .in0(_gnd_net_),
            .in1(N__67602),
            .in2(N__67596),
            .in3(N__67593),
            .lcout(\pid_front.N_39_0 ),
            .ltout(\pid_front.N_39_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_1_c_RNIKLQF7_LC_16_21_4 .C_ON=1'b0;
    defparam \pid_front.error_cry_1_c_RNIKLQF7_LC_16_21_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_1_c_RNIKLQF7_LC_16_21_4 .LUT_INIT=16'b0001010110011101;
    LogicCell40 \pid_front.error_cry_1_c_RNIKLQF7_LC_16_21_4  (
            .in0(N__77393),
            .in1(N__67579),
            .in2(N__67539),
            .in3(N__76372),
            .lcout(),
            .ltout(\pid_front.m53_0_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_1_c_RNI78AMF_LC_16_21_5 .C_ON=1'b0;
    defparam \pid_front.error_cry_1_c_RNI78AMF_LC_16_21_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_1_c_RNI78AMF_LC_16_21_5 .LUT_INIT=16'b0101111000001110;
    LogicCell40 \pid_front.error_cry_1_c_RNI78AMF_LC_16_21_5  (
            .in0(N__76281),
            .in1(N__76054),
            .in2(N__67536),
            .in3(N__71306),
            .lcout(\pid_front.N_54_0 ),
            .ltout(\pid_front.N_54_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_11_LC_16_21_6 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_11_LC_16_21_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_11_LC_16_21_6 .LUT_INIT=16'b0011101100001000;
    LogicCell40 \pid_front.error_i_reg_11_LC_16_21_6  (
            .in0(N__75488),
            .in1(N__67532),
            .in2(N__67497),
            .in3(N__67487),
            .lcout(\pid_front.error_i_regZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87186),
            .ce(),
            .sr(N__79693));
    defparam \pid_front.error_i_reg_esr_27_LC_16_22_0 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_27_LC_16_22_0 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_esr_27_LC_16_22_0 .LUT_INIT=16'b0000100011001000;
    LogicCell40 \pid_front.error_i_reg_esr_27_LC_16_22_0  (
            .in0(N__71133),
            .in1(N__76546),
            .in2(N__76984),
            .in3(N__67473),
            .lcout(\pid_front.error_i_regZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87201),
            .ce(N__72416),
            .sr(N__79697));
    defparam \pid_front.error_i_reg_esr_RNO_3_19_LC_16_22_1 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_3_19_LC_16_22_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_3_19_LC_16_22_1 .LUT_INIT=16'b0000000100001011;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_3_19_LC_16_22_1  (
            .in0(N__77739),
            .in1(N__76093),
            .in2(N__80340),
            .in3(N__76382),
            .lcout(),
            .ltout(\pid_front.m7_2_03_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_0_19_LC_16_22_2 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_0_19_LC_16_22_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_0_19_LC_16_22_2 .LUT_INIT=16'b1110001000000000;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_0_19_LC_16_22_2  (
            .in0(N__71132),
            .in1(N__76885),
            .in2(N__67974),
            .in3(N__76545),
            .lcout(),
            .ltout(\pid_front.error_i_reg_9_rn_0_19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_19_LC_16_22_3 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_19_LC_16_22_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_esr_19_LC_16_22_3 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \pid_front.error_i_reg_esr_19_LC_16_22_3  (
            .in0(_gnd_net_),
            .in1(N__71235),
            .in2(N__67971),
            .in3(N__67953),
            .lcout(\pid_front.error_i_regZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87201),
            .ce(N__72416),
            .sr(N__79697));
    defparam \pid_front.error_i_reg_9_sn_19_LC_16_22_4 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_9_sn_19_LC_16_22_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_9_sn_19_LC_16_22_4 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \pid_front.error_i_reg_9_sn_19_LC_16_22_4  (
            .in0(N__80287),
            .in1(N__76884),
            .in2(_gnd_net_),
            .in3(N__76544),
            .lcout(pid_front_error_i_reg_9_sn_19),
            .ltout(pid_front_error_i_reg_9_sn_19_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_2_19_LC_16_22_5 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_2_19_LC_16_22_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_2_19_LC_16_22_5 .LUT_INIT=16'b0100111101111111;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_2_19_LC_16_22_5  (
            .in0(N__76067),
            .in1(N__80599),
            .in2(N__67956),
            .in3(N__71307),
            .lcout(\pid_front.error_i_reg_esr_RNO_2Z0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_0_7_LC_16_22_7 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_0_7_LC_16_22_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_0_7_LC_16_22_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_0_7_LC_16_22_7  (
            .in0(N__76066),
            .in1(N__77738),
            .in2(_gnd_net_),
            .in3(N__76094),
            .lcout(\pid_front.N_103_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_6_LC_16_23_0 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_6_LC_16_23_0 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_esr_6_LC_16_23_0 .LUT_INIT=16'b1000000011010000;
    LogicCell40 \pid_front.error_i_reg_esr_6_LC_16_23_0  (
            .in0(N__75732),
            .in1(N__67947),
            .in2(N__75534),
            .in3(N__67935),
            .lcout(\pid_front.error_i_regZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87219),
            .ce(N__72415),
            .sr(N__79703));
    defparam \pid_front.error_i_reg_esr_7_LC_16_23_1 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_7_LC_16_23_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_esr_7_LC_16_23_1 .LUT_INIT=16'b1100010000000100;
    LogicCell40 \pid_front.error_i_reg_esr_7_LC_16_23_1  (
            .in0(N__67902),
            .in1(N__75518),
            .in2(N__75752),
            .in3(N__76344),
            .lcout(\pid_front.error_i_regZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87219),
            .ce(N__72415),
            .sr(N__79703));
    defparam \pid_front.error_i_reg_esr_9_LC_16_23_3 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_9_LC_16_23_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_esr_9_LC_16_23_3 .LUT_INIT=16'b1101000000010000;
    LogicCell40 \pid_front.error_i_reg_esr_9_LC_16_23_3  (
            .in0(N__72168),
            .in1(N__75733),
            .in2(N__75536),
            .in3(N__68097),
            .lcout(\pid_front.error_i_regZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87219),
            .ce(N__72415),
            .sr(N__79703));
    defparam \pid_front.error_i_reg_esr_RNO_1_25_LC_16_23_4 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_1_25_LC_16_23_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_1_25_LC_16_23_4 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_1_25_LC_16_23_4  (
            .in0(N__68112),
            .in1(N__72133),
            .in2(_gnd_net_),
            .in3(N__71179),
            .lcout(),
            .ltout(\pid_front.error_i_reg_esr_RNO_1Z0Z_25_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_0_25_LC_16_23_5 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_0_25_LC_16_23_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_0_25_LC_16_23_5 .LUT_INIT=16'b1000110000000100;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_0_25_LC_16_23_5  (
            .in0(N__76980),
            .in1(N__76552),
            .in2(N__68100),
            .in3(N__68096),
            .lcout(),
            .ltout(\pid_front.error_i_reg_9_rn_1_25_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_25_LC_16_23_6 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_25_LC_16_23_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_esr_25_LC_16_23_6 .LUT_INIT=16'b0101000011111010;
    LogicCell40 \pid_front.error_i_reg_esr_25_LC_16_23_6  (
            .in0(N__68294),
            .in1(_gnd_net_),
            .in2(N__68085),
            .in3(N__72167),
            .lcout(\pid_front.error_i_regZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87219),
            .ce(N__72415),
            .sr(N__79703));
    defparam \pid_front.error_i_reg_esr_8_LC_16_23_7 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_8_LC_16_23_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_esr_8_LC_16_23_7 .LUT_INIT=16'b1011000000010000;
    LogicCell40 \pid_front.error_i_reg_esr_8_LC_16_23_7  (
            .in0(N__75734),
            .in1(N__68070),
            .in2(N__75535),
            .in3(N__68064),
            .lcout(\pid_front.error_i_regZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87219),
            .ce(N__72415),
            .sr(N__79703));
    defparam \pid_front.error_i_reg_esr_RNO_0_13_LC_16_24_0 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_0_13_LC_16_24_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_0_13_LC_16_24_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_0_13_LC_16_24_0  (
            .in0(N__80614),
            .in1(N__68028),
            .in2(_gnd_net_),
            .in3(N__68037),
            .lcout(\pid_front.N_127 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_3_13_LC_16_24_1 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_3_13_LC_16_24_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_3_13_LC_16_24_1 .LUT_INIT=16'b0100000001111111;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_3_13_LC_16_24_1  (
            .in0(N__72132),
            .in1(N__80795),
            .in2(N__72063),
            .in3(N__71167),
            .lcout(\pid_front.N_126_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_1_13_LC_16_24_2 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_1_13_LC_16_24_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_1_13_LC_16_24_2 .LUT_INIT=16'b1000000010001010;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_1_13_LC_16_24_2  (
            .in0(N__76624),
            .in1(N__68301),
            .in2(N__77031),
            .in3(N__68022),
            .lcout(),
            .ltout(\pid_front.error_i_reg_9_rn_1_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_13_LC_16_24_3 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_13_LC_16_24_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_esr_13_LC_16_24_3 .LUT_INIT=16'b0011000011111100;
    LogicCell40 \pid_front.error_i_reg_esr_13_LC_16_24_3  (
            .in0(_gnd_net_),
            .in1(N__70964),
            .in2(N__68010),
            .in3(N__68007),
            .lcout(\pid_front.error_i_regZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87233),
            .ce(N__72422),
            .sr(N__79708));
    defparam \pid_front.error_cry_0_c_RNI3FL31_LC_16_24_4 .C_ON=1'b0;
    defparam \pid_front.error_cry_0_c_RNI3FL31_LC_16_24_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_0_c_RNI3FL31_LC_16_24_4 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \pid_front.error_cry_0_c_RNI3FL31_LC_16_24_4  (
            .in0(N__80794),
            .in1(N__77263),
            .in2(N__78097),
            .in3(N__77185),
            .lcout(\pid_front.m1_0_03 ),
            .ltout(\pid_front.m1_0_03_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_4_13_LC_16_24_5 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_4_13_LC_16_24_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_4_13_LC_16_24_5 .LUT_INIT=16'b0000000000110000;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_4_13_LC_16_24_5  (
            .in0(_gnd_net_),
            .in1(N__80338),
            .in2(N__68304),
            .in3(N__77780),
            .lcout(\pid_front.m1_2_03 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_1_17_LC_16_25_2 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_1_17_LC_16_25_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_1_17_LC_16_25_2 .LUT_INIT=16'b0101000000000000;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_1_17_LC_16_25_2  (
            .in0(N__76961),
            .in1(_gnd_net_),
            .in2(N__76322),
            .in3(N__76551),
            .lcout(\pid_front.error_i_reg_9_sn_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_9_sn_27_LC_16_25_3 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_9_sn_27_LC_16_25_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_9_sn_27_LC_16_25_3 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \pid_side.error_i_reg_9_sn_27_LC_16_25_3  (
            .in0(N__76547),
            .in1(N__76955),
            .in2(_gnd_net_),
            .in3(N__76311),
            .lcout(pid_side_error_i_reg_9_sn_27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_4_LC_16_25_4 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_4_LC_16_25_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_esr_4_LC_16_25_4 .LUT_INIT=16'b1011000010000000;
    LogicCell40 \pid_front.error_i_reg_esr_4_LC_16_25_4  (
            .in0(N__68253),
            .in1(N__76318),
            .in2(N__75533),
            .in3(N__68226),
            .lcout(\pid_front.error_i_regZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87245),
            .ce(N__72406),
            .sr(N__79711));
    defparam \pid_side.error_i_reg_esr_RNO_1_17_LC_16_25_5 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_1_17_LC_16_25_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_1_17_LC_16_25_5 .LUT_INIT=16'b0010000000100000;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_1_17_LC_16_25_5  (
            .in0(N__76549),
            .in1(N__76959),
            .in2(N__75750),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_i_reg_9_sn_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_1_25_LC_16_25_6 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_1_25_LC_16_25_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_1_25_LC_16_25_6 .LUT_INIT=16'b0011000000000000;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_1_25_LC_16_25_6  (
            .in0(_gnd_net_),
            .in1(N__75725),
            .in2(N__77004),
            .in3(N__76548),
            .lcout(\pid_side.error_i_reg_9_sn_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_2_13_LC_16_25_7 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_2_13_LC_16_25_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_2_13_LC_16_25_7 .LUT_INIT=16'b0000001000000010;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_2_13_LC_16_25_7  (
            .in0(N__76550),
            .in1(N__76960),
            .in2(N__75751),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_i_reg_9_sn_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_3_LC_17_3_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_3_LC_17_3_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_3_LC_17_3_0 .LUT_INIT=16'b1111111011101110;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_3_LC_17_3_0  (
            .in0(N__68813),
            .in1(N__68562),
            .in2(N__68178),
            .in3(N__68904),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__86996),
            .ce(N__68769),
            .sr(N__79593));
    defparam \ppm_encoder_1.pulses2count_esr_2_LC_17_3_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_2_LC_17_3_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_2_LC_17_3_3 .LUT_INIT=16'b0000000000110001;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_2_LC_17_3_3  (
            .in0(N__68903),
            .in1(N__68859),
            .in2(N__68853),
            .in3(N__68814),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__86996),
            .ce(N__68769),
            .sr(N__79593));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_3_LC_17_4_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_3_LC_17_4_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_3_LC_17_4_3 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_3_LC_17_4_3  (
            .in0(N__68676),
            .in1(N__68607),
            .in2(_gnd_net_),
            .in3(N__68594),
            .lcout(\ppm_encoder_1.pulses2count_9_0_0_3_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_45_c_RNO_LC_17_4_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_45_c_RNO_LC_17_4_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_45_c_RNO_LC_17_4_5 .LUT_INIT=16'b0110111111110110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_45_c_RNO_LC_17_4_5  (
            .in0(N__68554),
            .in1(N__68538),
            .in2(N__68526),
            .in3(N__68506),
            .lcout(\ppm_encoder_1.counter24_0_I_45_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter_RNIS9KG_2_LC_17_4_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter_RNIS9KG_2_LC_17_4_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter_RNIS9KG_2_LC_17_4_6 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \ppm_encoder_1.counter_RNIS9KG_2_LC_17_4_6  (
            .in0(N__68481),
            .in1(N__68456),
            .in2(N__68439),
            .in3(N__68411),
            .lcout(\ppm_encoder_1.un1_PPM_STATE_0_sqmuxa_0_i_a2_18_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_esr_RNIF3BO1_1_LC_17_8_4 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_esr_RNIF3BO1_1_LC_17_8_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_esr_RNIF3BO1_1_LC_17_8_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_side.pid_prereg_esr_RNIF3BO1_1_LC_17_8_4  (
            .in0(N__69373),
            .in1(N__69115),
            .in2(N__69085),
            .in3(N__69145),
            .lcout(\pid_side.source_pid_1_sqmuxa_1_0_a4_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_12_LC_17_9_0 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_12_LC_17_9_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_12_LC_17_9_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_12_LC_17_9_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78783),
            .lcout(\pid_side.un10lto12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87044),
            .ce(N__69895),
            .sr(N__79628));
    defparam \pid_side.error_i_acumm_prereg_esr_21_LC_17_9_1 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_21_LC_17_9_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_21_LC_17_9_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_21_LC_17_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73044),
            .lcout(\pid_side.error_i_acumm_preregZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87044),
            .ce(N__69895),
            .sr(N__79628));
    defparam \pid_side.error_i_acumm_prereg_esr_13_LC_17_9_2 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_13_LC_17_9_2 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_13_LC_17_9_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_13_LC_17_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81983),
            .lcout(\pid_side.error_i_acumm_preregZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87044),
            .ce(N__69895),
            .sr(N__79628));
    defparam \pid_side.error_i_acumm_prereg_esr_22_LC_17_9_3 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_22_LC_17_9_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_22_LC_17_9_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_22_LC_17_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__69840),
            .lcout(\pid_side.error_i_acumm_preregZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87044),
            .ce(N__69895),
            .sr(N__79628));
    defparam \pid_side.error_i_acumm_prereg_esr_23_LC_17_9_4 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_23_LC_17_9_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_23_LC_17_9_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_23_LC_17_9_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__69237),
            .lcout(\pid_side.error_i_acumm_preregZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87044),
            .ce(N__69895),
            .sr(N__79628));
    defparam \pid_side.error_i_acumm_prereg_esr_24_LC_17_9_5 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_24_LC_17_9_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_24_LC_17_9_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_24_LC_17_9_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68928),
            .lcout(\pid_side.error_i_acumm_preregZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87044),
            .ce(N__69895),
            .sr(N__79628));
    defparam \pid_side.error_i_acumm_prereg_esr_17_LC_17_9_6 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_17_LC_17_9_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_17_LC_17_9_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_17_LC_17_9_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70098),
            .lcout(\pid_side.error_i_acumm_preregZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87044),
            .ce(N__69895),
            .sr(N__79628));
    defparam \pid_side.error_i_acumm_prereg_esr_5_LC_17_9_7 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_5_LC_17_9_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_acumm_prereg_esr_5_LC_17_9_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_5_LC_17_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78513),
            .lcout(\pid_side.error_i_acumm_preregZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87044),
            .ce(N__69895),
            .sr(N__79628));
    defparam \pid_side.error_d_reg_prev_esr_RNIR5HL1_0_22_LC_17_10_0 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIR5HL1_0_22_LC_17_10_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIR5HL1_0_22_LC_17_10_0 .LUT_INIT=16'b0001100011100111;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIR5HL1_0_22_LC_17_10_0  (
            .in0(N__84625),
            .in1(N__83533),
            .in2(N__73209),
            .in3(N__68924),
            .lcout(\pid_side.un1_pid_prereg_0_17 ),
            .ltout(\pid_side.un1_pid_prereg_0_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIK81B3_22_LC_17_10_1 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIK81B3_22_LC_17_10_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIK81B3_22_LC_17_10_1 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIK81B3_22_LC_17_10_1  (
            .in0(N__69209),
            .in1(_gnd_net_),
            .in2(N__68967),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIK81B3Z0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI33ME7_22_LC_17_10_2 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI33ME7_22_LC_17_10_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI33ME7_22_LC_17_10_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI33ME7_22_LC_17_10_2  (
            .in0(N__68964),
            .in1(N__69208),
            .in2(N__68949),
            .in3(N__69251),
            .lcout(\pid_side.error_d_reg_prev_esr_RNI33ME7Z0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIR5HL1_22_LC_17_10_3 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIR5HL1_22_LC_17_10_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIR5HL1_22_LC_17_10_3 .LUT_INIT=16'b1011101010100010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIR5HL1_22_LC_17_10_3  (
            .in0(N__68923),
            .in1(N__73194),
            .in2(N__83552),
            .in3(N__84629),
            .lcout(\pid_side.un1_pid_prereg_0_18 ),
            .ltout(\pid_side.un1_pid_prereg_0_18_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNICN4M6_22_LC_17_10_4 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNICN4M6_22_LC_17_10_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNICN4M6_22_LC_17_10_4 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNICN4M6_22_LC_17_10_4  (
            .in0(N__69252),
            .in1(N__72848),
            .in2(N__69240),
            .in3(N__69210),
            .lcout(\pid_side.error_d_reg_prev_esr_RNICN4M6Z0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIP2GL1_22_LC_17_10_5 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIP2GL1_22_LC_17_10_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIP2GL1_22_LC_17_10_5 .LUT_INIT=16'b1110111100001000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIP2GL1_22_LC_17_10_5  (
            .in0(N__83532),
            .in1(N__84624),
            .in2(N__73208),
            .in3(N__69235),
            .lcout(\pid_side.un1_pid_prereg_0_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIT8IL1_0_22_LC_17_10_6 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIT8IL1_0_22_LC_17_10_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIT8IL1_0_22_LC_17_10_6 .LUT_INIT=16'b0101011010010101;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIT8IL1_0_22_LC_17_10_6  (
            .in0(N__72899),
            .in1(N__83537),
            .in2(N__84633),
            .in3(N__73190),
            .lcout(\pid_side.un1_pid_prereg_0_19 ),
            .ltout(\pid_side.un1_pid_prereg_0_19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIOE3B3_22_LC_17_10_7 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIOE3B3_22_LC_17_10_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIOE3B3_22_LC_17_10_7 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIOE3B3_22_LC_17_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__69198),
            .in3(N__72866),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIOE3B3Z0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un1_pid_prereg_0_cry_0_c_THRU_CRY_0_LC_17_11_0 .C_ON=1'b1;
    defparam \pid_side.un1_pid_prereg_0_cry_0_c_THRU_CRY_0_LC_17_11_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.un1_pid_prereg_0_cry_0_c_THRU_CRY_0_LC_17_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_side.un1_pid_prereg_0_cry_0_c_THRU_CRY_0_LC_17_11_0  (
            .in0(_gnd_net_),
            .in1(N__84500),
            .in2(N__84504),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_17_11_0_),
            .carryout(\pid_side.un1_pid_prereg_0_cry_0_c_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_esr_0_LC_17_11_1 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_0_LC_17_11_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_0_LC_17_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_0_LC_17_11_1  (
            .in0(_gnd_net_),
            .in1(N__73691),
            .in2(N__73674),
            .in3(N__69156),
            .lcout(\pid_side.pid_preregZ0Z_0 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_0_cry_0_c_THRU_CO ),
            .carryout(\pid_side.un1_pid_prereg_0_cry_0 ),
            .clk(N__87061),
            .ce(N__69896),
            .sr(N__79645));
    defparam \pid_side.pid_prereg_esr_1_LC_17_11_2 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_1_LC_17_11_2 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_1_LC_17_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_1_LC_17_11_2  (
            .in0(_gnd_net_),
            .in1(N__72453),
            .in2(N__72485),
            .in3(N__69120),
            .lcout(\pid_side.pid_preregZ0Z_1 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_0_cry_0 ),
            .carryout(\pid_side.un1_pid_prereg_0_cry_1 ),
            .clk(N__87061),
            .ce(N__69896),
            .sr(N__79645));
    defparam \pid_side.pid_prereg_esr_2_LC_17_11_3 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_2_LC_17_11_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_2_LC_17_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_2_LC_17_11_3  (
            .in0(_gnd_net_),
            .in1(N__82131),
            .in2(N__82166),
            .in3(N__69093),
            .lcout(\pid_side.pid_preregZ0Z_2 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_0_cry_1 ),
            .carryout(\pid_side.un1_pid_prereg_0_cry_2 ),
            .clk(N__87061),
            .ce(N__69896),
            .sr(N__79645));
    defparam \pid_side.pid_prereg_esr_3_LC_17_11_4 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_3_LC_17_11_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_3_LC_17_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_3_LC_17_11_4  (
            .in0(_gnd_net_),
            .in1(N__82199),
            .in2(N__81750),
            .in3(N__69048),
            .lcout(\pid_side.pid_preregZ0Z_3 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_0_cry_2 ),
            .carryout(\pid_side.un1_pid_prereg_0_cry_3 ),
            .clk(N__87061),
            .ce(N__69896),
            .sr(N__79645));
    defparam \pid_side.pid_prereg_esr_4_LC_17_11_5 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_4_LC_17_11_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_4_LC_17_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_4_LC_17_11_5  (
            .in0(_gnd_net_),
            .in1(N__81462),
            .in2(N__81447),
            .in3(N__69378),
            .lcout(\pid_side.pid_preregZ0Z_4 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_0_cry_3 ),
            .carryout(\pid_side.un1_pid_prereg_0_cry_4 ),
            .clk(N__87061),
            .ce(N__69896),
            .sr(N__79645));
    defparam \pid_side.pid_prereg_esr_5_LC_17_11_6 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_5_LC_17_11_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_5_LC_17_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_5_LC_17_11_6  (
            .in0(_gnd_net_),
            .in1(N__81605),
            .in2(N__81585),
            .in3(N__69342),
            .lcout(\pid_side.pid_preregZ0Z_5 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_0_cry_4 ),
            .carryout(\pid_side.un1_pid_prereg_0_cry_5 ),
            .clk(N__87061),
            .ce(N__69896),
            .sr(N__79645));
    defparam \pid_side.pid_prereg_esr_6_LC_17_11_7 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_6_LC_17_11_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_6_LC_17_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_6_LC_17_11_7  (
            .in0(_gnd_net_),
            .in1(N__78456),
            .in2(N__78633),
            .in3(N__69339),
            .lcout(\pid_side.pid_preregZ0Z_6 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_0_cry_5 ),
            .carryout(\pid_side.un1_pid_prereg_0_cry_6 ),
            .clk(N__87061),
            .ce(N__69896),
            .sr(N__79645));
    defparam \pid_side.pid_prereg_esr_7_LC_17_12_0 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_7_LC_17_12_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_7_LC_17_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_7_LC_17_12_0  (
            .in0(_gnd_net_),
            .in1(N__69336),
            .in2(N__72498),
            .in3(N__69327),
            .lcout(\pid_side.pid_preregZ0Z_7 ),
            .ltout(),
            .carryin(bfn_17_12_0_),
            .carryout(\pid_side.un1_pid_prereg_0_cry_7 ),
            .clk(N__87069),
            .ce(N__69897),
            .sr(N__79652));
    defparam \pid_side.pid_prereg_esr_8_LC_17_12_1 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_8_LC_17_12_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_8_LC_17_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_8_LC_17_12_1  (
            .in0(_gnd_net_),
            .in1(N__69324),
            .in2(N__69315),
            .in3(N__69297),
            .lcout(\pid_side.pid_preregZ0Z_8 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_0_cry_7 ),
            .carryout(\pid_side.un1_pid_prereg_0_cry_8 ),
            .clk(N__87069),
            .ce(N__69897),
            .sr(N__79652));
    defparam \pid_side.pid_prereg_esr_9_LC_17_12_2 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_9_LC_17_12_2 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_9_LC_17_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_9_LC_17_12_2  (
            .in0(_gnd_net_),
            .in1(N__69294),
            .in2(N__69284),
            .in3(N__69261),
            .lcout(\pid_side.pid_preregZ0Z_9 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_0_cry_8 ),
            .carryout(\pid_side.un1_pid_prereg_0_cry_9 ),
            .clk(N__87069),
            .ce(N__69897),
            .sr(N__79652));
    defparam \pid_side.pid_prereg_esr_10_LC_17_12_3 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_10_LC_17_12_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_10_LC_17_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_10_LC_17_12_3  (
            .in0(_gnd_net_),
            .in1(N__72978),
            .in2(N__73001),
            .in3(N__69258),
            .lcout(\pid_side.pid_preregZ0Z_10 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_0_cry_9 ),
            .carryout(\pid_side.un1_pid_prereg_0_cry_10 ),
            .clk(N__87069),
            .ce(N__69897),
            .sr(N__79652));
    defparam \pid_side.pid_prereg_esr_11_LC_17_12_4 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_11_LC_17_12_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_11_LC_17_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_11_LC_17_12_4  (
            .in0(_gnd_net_),
            .in1(N__72962),
            .in2(N__72909),
            .in3(N__69255),
            .lcout(\pid_side.pid_preregZ0Z_11 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_0_cry_10 ),
            .carryout(\pid_side.un1_pid_prereg_0_cry_11 ),
            .clk(N__87069),
            .ce(N__69897),
            .sr(N__79652));
    defparam \pid_side.pid_prereg_esr_12_LC_17_12_5 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_12_LC_17_12_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_12_LC_17_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_12_LC_17_12_5  (
            .in0(_gnd_net_),
            .in1(N__78828),
            .in2(N__69519),
            .in3(N__69465),
            .lcout(\pid_side.pid_preregZ0Z_12 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_0_cry_11 ),
            .carryout(\pid_side.un1_pid_prereg_0_cry_12 ),
            .clk(N__87069),
            .ce(N__69897),
            .sr(N__79652));
    defparam \pid_side.pid_prereg_esr_13_LC_17_12_6 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_13_LC_17_12_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_13_LC_17_12_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_13_LC_17_12_6  (
            .in0(_gnd_net_),
            .in1(N__78752),
            .in2(N__78738),
            .in3(N__69462),
            .lcout(\pid_side.pid_preregZ0Z_13 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_0_cry_12 ),
            .carryout(\pid_side.un1_pid_prereg_0_cry_13 ),
            .clk(N__87069),
            .ce(N__69897),
            .sr(N__79652));
    defparam \pid_side.un1_pid_prereg_0_cry_13_THRU_LUT4_0_LC_17_12_7 .C_ON=1'b1;
    defparam \pid_side.un1_pid_prereg_0_cry_13_THRU_LUT4_0_LC_17_12_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.un1_pid_prereg_0_cry_13_THRU_LUT4_0_LC_17_12_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.un1_pid_prereg_0_cry_13_THRU_LUT4_0_LC_17_12_7  (
            .in0(_gnd_net_),
            .in1(N__81926),
            .in2(_gnd_net_),
            .in3(N__69450),
            .lcout(\pid_side.un1_pid_prereg_0_cry_13_THRU_CO ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_0_cry_13 ),
            .carryout(\pid_side.un1_pid_prereg_0_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_esr_15_LC_17_13_0 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_15_LC_17_13_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_15_LC_17_13_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_15_LC_17_13_0  (
            .in0(_gnd_net_),
            .in1(N__80091),
            .in2(N__80022),
            .in3(N__69447),
            .lcout(\pid_side.pid_preregZ0Z_15 ),
            .ltout(),
            .carryin(bfn_17_13_0_),
            .carryout(\pid_side.un1_pid_prereg_0_cry_15 ),
            .clk(N__87081),
            .ce(N__69898),
            .sr(N__79661));
    defparam \pid_side.pid_prereg_esr_16_LC_17_13_1 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_16_LC_17_13_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_16_LC_17_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_16_LC_17_13_1  (
            .in0(_gnd_net_),
            .in1(N__78927),
            .in2(N__73359),
            .in3(N__69444),
            .lcout(\pid_side.pid_preregZ0Z_16 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_0_cry_15 ),
            .carryout(\pid_side.un1_pid_prereg_0_cry_16 ),
            .clk(N__87081),
            .ce(N__69898),
            .sr(N__79661));
    defparam \pid_side.pid_prereg_esr_17_LC_17_13_2 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_17_LC_17_13_2 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_17_LC_17_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_17_LC_17_13_2  (
            .in0(_gnd_net_),
            .in1(N__69771),
            .in2(N__69804),
            .in3(N__69441),
            .lcout(\pid_side.pid_preregZ0Z_17 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_0_cry_16 ),
            .carryout(\pid_side.un1_pid_prereg_0_cry_17 ),
            .clk(N__87081),
            .ce(N__69898),
            .sr(N__79661));
    defparam \pid_side.pid_prereg_esr_18_LC_17_13_3 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_18_LC_17_13_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_18_LC_17_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_18_LC_17_13_3  (
            .in0(_gnd_net_),
            .in1(N__70176),
            .in2(N__73449),
            .in3(N__69438),
            .lcout(\pid_side.pid_preregZ0Z_18 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_0_cry_17 ),
            .carryout(\pid_side.un1_pid_prereg_0_cry_18 ),
            .clk(N__87081),
            .ce(N__69898),
            .sr(N__79661));
    defparam \pid_side.pid_prereg_esr_19_LC_17_13_4 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_19_LC_17_13_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_19_LC_17_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_19_LC_17_13_4  (
            .in0(_gnd_net_),
            .in1(N__70122),
            .in2(N__70164),
            .in3(N__69435),
            .lcout(\pid_side.pid_preregZ0Z_19 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_0_cry_18 ),
            .carryout(\pid_side.un1_pid_prereg_0_cry_19 ),
            .clk(N__87081),
            .ce(N__69898),
            .sr(N__79661));
    defparam \pid_side.pid_prereg_esr_20_LC_17_13_5 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_20_LC_17_13_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_20_LC_17_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_20_LC_17_13_5  (
            .in0(_gnd_net_),
            .in1(N__73299),
            .in2(N__70110),
            .in3(N__69420),
            .lcout(\pid_side.pid_preregZ0Z_20 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_0_cry_19 ),
            .carryout(\pid_side.un1_pid_prereg_0_cry_20 ),
            .clk(N__87081),
            .ce(N__69898),
            .sr(N__79661));
    defparam \pid_side.pid_prereg_esr_21_LC_17_13_6 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_21_LC_17_13_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_21_LC_17_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_21_LC_17_13_6  (
            .in0(_gnd_net_),
            .in1(N__73080),
            .in2(N__73710),
            .in3(N__69750),
            .lcout(\pid_side.pid_preregZ0Z_21 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_0_cry_20 ),
            .carryout(\pid_side.un1_pid_prereg_0_cry_21 ),
            .clk(N__87081),
            .ce(N__69898),
            .sr(N__79661));
    defparam \pid_side.pid_prereg_esr_22_LC_17_13_7 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_22_LC_17_13_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_22_LC_17_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_22_LC_17_13_7  (
            .in0(_gnd_net_),
            .in1(N__73488),
            .in2(N__73071),
            .in3(N__69735),
            .lcout(\pid_side.pid_preregZ0Z_22 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_0_cry_21 ),
            .carryout(\pid_side.un1_pid_prereg_0_cry_22 ),
            .clk(N__87081),
            .ce(N__69898),
            .sr(N__79661));
    defparam \pid_side.pid_prereg_esr_23_LC_17_14_0 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_23_LC_17_14_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_23_LC_17_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_23_LC_17_14_0  (
            .in0(_gnd_net_),
            .in1(N__73398),
            .in2(N__69732),
            .in3(N__69702),
            .lcout(\pid_side.pid_preregZ0Z_23 ),
            .ltout(),
            .carryin(bfn_17_14_0_),
            .carryout(\pid_side.un1_pid_prereg_0_cry_23 ),
            .clk(N__87095),
            .ce(N__69899),
            .sr(N__79668));
    defparam \pid_side.pid_prereg_esr_24_LC_17_14_1 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_24_LC_17_14_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_24_LC_17_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_24_LC_17_14_1  (
            .in0(_gnd_net_),
            .in1(N__69699),
            .in2(N__69690),
            .in3(N__69663),
            .lcout(\pid_side.pid_preregZ0Z_24 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_0_cry_23 ),
            .carryout(\pid_side.un1_pid_prereg_0_cry_24 ),
            .clk(N__87095),
            .ce(N__69899),
            .sr(N__79668));
    defparam \pid_side.pid_prereg_esr_25_LC_17_14_2 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_25_LC_17_14_2 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_25_LC_17_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_25_LC_17_14_2  (
            .in0(_gnd_net_),
            .in1(N__69660),
            .in2(N__69651),
            .in3(N__69624),
            .lcout(\pid_side.pid_preregZ0Z_25 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_0_cry_24 ),
            .carryout(\pid_side.un1_pid_prereg_0_cry_25 ),
            .clk(N__87095),
            .ce(N__69899),
            .sr(N__79668));
    defparam \pid_side.pid_prereg_esr_26_LC_17_14_3 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_26_LC_17_14_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_26_LC_17_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_26_LC_17_14_3  (
            .in0(_gnd_net_),
            .in1(N__72834),
            .in2(N__69621),
            .in3(N__69591),
            .lcout(\pid_side.pid_preregZ0Z_26 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_0_cry_25 ),
            .carryout(\pid_side.un1_pid_prereg_0_cry_26 ),
            .clk(N__87095),
            .ce(N__69899),
            .sr(N__79668));
    defparam \pid_side.pid_prereg_esr_27_LC_17_14_4 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_27_LC_17_14_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_27_LC_17_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_27_LC_17_14_4  (
            .in0(_gnd_net_),
            .in1(N__73218),
            .in2(N__69588),
            .in3(N__69558),
            .lcout(\pid_side.pid_preregZ0Z_27 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_0_cry_26 ),
            .carryout(\pid_side.un1_pid_prereg_0_cry_27 ),
            .clk(N__87095),
            .ce(N__69899),
            .sr(N__79668));
    defparam \pid_side.pid_prereg_esr_28_LC_17_14_5 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_28_LC_17_14_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_28_LC_17_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_28_LC_17_14_5  (
            .in0(_gnd_net_),
            .in1(N__69555),
            .in2(N__69546),
            .in3(N__69522),
            .lcout(\pid_side.pid_preregZ0Z_28 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_0_cry_27 ),
            .carryout(\pid_side.un1_pid_prereg_0_cry_28 ),
            .clk(N__87095),
            .ce(N__69899),
            .sr(N__79668));
    defparam \pid_side.pid_prereg_esr_29_LC_17_14_6 .C_ON=1'b1;
    defparam \pid_side.pid_prereg_esr_29_LC_17_14_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_29_LC_17_14_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.pid_prereg_esr_29_LC_17_14_6  (
            .in0(_gnd_net_),
            .in1(N__70062),
            .in2(N__70053),
            .in3(N__70026),
            .lcout(\pid_side.pid_preregZ0Z_29 ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_0_cry_28 ),
            .carryout(\pid_side.un1_pid_prereg_0_cry_29 ),
            .clk(N__87095),
            .ce(N__69899),
            .sr(N__79668));
    defparam \pid_side.pid_prereg_esr_30_LC_17_14_7 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_esr_30_LC_17_14_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_30_LC_17_14_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_side.pid_prereg_esr_30_LC_17_14_7  (
            .in0(_gnd_net_),
            .in1(N__70023),
            .in2(_gnd_net_),
            .in3(N__70014),
            .lcout(\pid_side.pid_preregZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87095),
            .ce(N__69899),
            .sr(N__79668));
    defparam \pid_side.error_d_reg_prev_esr_RNIMN4E2_0_21_LC_17_15_0 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIMN4E2_0_21_LC_17_15_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIMN4E2_0_21_LC_17_15_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIMN4E2_0_21_LC_17_15_0  (
            .in0(N__69852),
            .in1(N__73103),
            .in2(_gnd_net_),
            .in3(N__69826),
            .lcout(\pid_side.un1_pid_prereg_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIFCVC2_0_15_LC_17_15_1 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIFCVC2_0_15_LC_17_15_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIFCVC2_0_15_LC_17_15_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIFCVC2_0_15_LC_17_15_1  (
            .in0(N__78938),
            .in1(N__69787),
            .in2(_gnd_net_),
            .in3(N__82919),
            .lcout(\pid_side.un1_pid_prereg_0_1 ),
            .ltout(\pid_side.un1_pid_prereg_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIMFTP4_14_LC_17_15_2 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIMFTP4_14_LC_17_15_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIMFTP4_14_LC_17_15_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIMFTP4_14_LC_17_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__69807),
            .in3(N__73373),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIMFTP4Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIFF3E2_0_20_LC_17_15_3 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIFF3E2_0_20_LC_17_15_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIFF3E2_0_20_LC_17_15_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIFF3E2_0_20_LC_17_15_3  (
            .in0(N__73059),
            .in1(N__82961),
            .in2(_gnd_net_),
            .in3(N__73030),
            .lcout(\pid_side.un1_pid_prereg_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIFCVC2_15_LC_17_15_4 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIFCVC2_15_LC_17_15_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIFCVC2_15_LC_17_15_4 .LUT_INIT=16'b1110100011101000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIFCVC2_15_LC_17_15_4  (
            .in0(N__69788),
            .in1(N__78939),
            .in2(N__82923),
            .in3(_gnd_net_),
            .lcout(\pid_side.un1_pid_prereg_0_2 ),
            .ltout(\pid_side.un1_pid_prereg_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNISHTJ9_14_LC_17_15_5 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNISHTJ9_14_LC_17_15_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNISHTJ9_14_LC_17_15_5 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNISHTJ9_14_LC_17_15_5  (
            .in0(N__73374),
            .in1(N__73389),
            .in2(N__69774),
            .in3(N__73465),
            .lcout(\pid_side.error_d_reg_prev_esr_RNISHTJ9Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI73UC2_14_LC_17_15_6 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI73UC2_14_LC_17_15_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI73UC2_14_LC_17_15_6 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI73UC2_14_LC_17_15_6  (
            .in0(N__79005),
            .in1(N__78963),
            .in2(_gnd_net_),
            .in3(N__78982),
            .lcout(\pid_side.un1_pid_prereg_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNINL0D2_0_16_LC_17_15_7 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNINL0D2_0_16_LC_17_15_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNINL0D2_0_16_LC_17_15_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNINL0D2_0_16_LC_17_15_7  (
            .in0(N__82650),
            .in1(N__82626),
            .in2(_gnd_net_),
            .in3(N__70091),
            .lcout(\pid_side.un1_pid_prereg_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNISM2K9_15_LC_17_16_0 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNISM2K9_15_LC_17_16_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNISM2K9_15_LC_17_16_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNISM2K9_15_LC_17_16_0  (
            .in0(N__70133),
            .in1(N__73482),
            .in2(N__73470),
            .in3(N__70072),
            .lcout(\pid_side.error_d_reg_prev_esr_RNISM2K9Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIVU1D2_0_17_LC_17_16_1 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIVU1D2_0_17_LC_17_16_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIVU1D2_0_17_LC_17_16_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIVU1D2_0_17_LC_17_16_1  (
            .in0(N__83423),
            .in1(N__83441),
            .in2(_gnd_net_),
            .in3(N__70147),
            .lcout(\pid_side.un1_pid_prereg_0_5 ),
            .ltout(\pid_side.un1_pid_prereg_0_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIMK2Q4_16_LC_17_16_2 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIMK2Q4_16_LC_17_16_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIMK2Q4_16_LC_17_16_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIMK2Q4_16_LC_17_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__70167),
            .in3(N__70073),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIMK2Q4Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIVU1D2_17_LC_17_16_3 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIVU1D2_17_LC_17_16_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIVU1D2_17_LC_17_16_3 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIVU1D2_17_LC_17_16_3  (
            .in0(N__83424),
            .in1(N__83442),
            .in2(_gnd_net_),
            .in3(N__70148),
            .lcout(\pid_side.un1_pid_prereg_0_6 ),
            .ltout(\pid_side.un1_pid_prereg_0_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNISR7K9_16_LC_17_16_4 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNISR7K9_16_LC_17_16_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNISR7K9_16_LC_17_16_4 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNISR7K9_16_LC_17_16_4  (
            .in0(N__70134),
            .in1(N__73325),
            .in2(N__70125),
            .in3(N__70074),
            .lcout(\pid_side.error_d_reg_prev_esr_RNISR7K9Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI783D2_0_18_LC_17_16_5 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI783D2_0_18_LC_17_16_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI783D2_0_18_LC_17_16_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI783D2_0_18_LC_17_16_5  (
            .in0(N__81734),
            .in1(N__83094),
            .in2(_gnd_net_),
            .in3(N__73342),
            .lcout(\pid_side.un1_pid_prereg_0_7 ),
            .ltout(\pid_side.un1_pid_prereg_0_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI675Q4_17_LC_17_16_6 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI675Q4_17_LC_17_16_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI675Q4_17_LC_17_16_6 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI675Q4_17_LC_17_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__70113),
            .in3(N__73313),
            .lcout(\pid_side.error_d_reg_prev_esr_RNI675Q4Z0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNINL0D2_16_LC_17_16_7 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNINL0D2_16_LC_17_16_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNINL0D2_16_LC_17_16_7 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNINL0D2_16_LC_17_16_7  (
            .in0(N__82625),
            .in1(N__82649),
            .in2(_gnd_net_),
            .in3(N__70090),
            .lcout(\pid_side.un1_pid_prereg_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_4_c_RNIMMS12_LC_17_17_0 .C_ON=1'b0;
    defparam \pid_side.error_cry_4_c_RNIMMS12_LC_17_17_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_4_c_RNIMMS12_LC_17_17_0 .LUT_INIT=16'b0010010100101111;
    LogicCell40 \pid_side.error_cry_4_c_RNIMMS12_LC_17_17_0  (
            .in0(N__77892),
            .in1(N__74624),
            .in2(N__75998),
            .in3(N__74547),
            .lcout(\pid_side.m21_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_6_12_LC_17_17_1 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_6_12_LC_17_17_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_6_12_LC_17_17_1 .LUT_INIT=16'b0000110001110111;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_6_12_LC_17_17_1  (
            .in0(N__74548),
            .in1(N__77751),
            .in2(N__74642),
            .in3(N__80780),
            .lcout(),
            .ltout(\pid_side.g0_i_m4_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_2_12_LC_17_17_2 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_2_12_LC_17_17_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_2_12_LC_17_17_2 .LUT_INIT=16'b1111000001010011;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_2_12_LC_17_17_2  (
            .in0(N__74382),
            .in1(N__74481),
            .in2(N__70254),
            .in3(N__77795),
            .lcout(\pid_side.N_8_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_8_c_RNI3TEU1_LC_17_17_3 .C_ON=1'b0;
    defparam \pid_side.error_cry_8_c_RNI3TEU1_LC_17_17_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_8_c_RNI3TEU1_LC_17_17_3 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \pid_side.error_cry_8_c_RNI3TEU1_LC_17_17_3  (
            .in0(N__80779),
            .in1(N__74479),
            .in2(_gnd_net_),
            .in3(N__74381),
            .lcout(\pid_side.N_36_0 ),
            .ltout(\pid_side.N_36_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_2_16_LC_17_17_4 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_2_16_LC_17_17_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_2_16_LC_17_17_4 .LUT_INIT=16'b1000000011110111;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_2_16_LC_17_17_4  (
            .in0(N__80532),
            .in1(N__72053),
            .in2(N__70242),
            .in3(N__74841),
            .lcout(\pid_side.error_i_reg_esr_RNO_2Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_1_24_LC_17_17_5 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_1_24_LC_17_17_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_1_24_LC_17_17_5 .LUT_INIT=16'b1111010100000101;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_1_24_LC_17_17_5  (
            .in0(N__74842),
            .in1(_gnd_net_),
            .in2(N__72062),
            .in3(N__70233),
            .lcout(),
            .ltout(\pid_side.N_57_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_0_24_LC_17_17_6 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_0_24_LC_17_17_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_0_24_LC_17_17_6 .LUT_INIT=16'b1000000011110111;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_0_24_LC_17_17_6  (
            .in0(N__71549),
            .in1(N__76267),
            .in2(N__70227),
            .in3(N__74843),
            .lcout(),
            .ltout(\pid_side.N_59_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_24_LC_17_17_7 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_24_LC_17_17_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_esr_24_LC_17_17_7 .LUT_INIT=16'b1000110000000100;
    LogicCell40 \pid_side.error_i_reg_esr_24_LC_17_17_7  (
            .in0(N__76946),
            .in1(N__76572),
            .in2(N__70224),
            .in3(N__70221),
            .lcout(\pid_side.error_i_regZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87139),
            .ce(N__75356),
            .sr(N__79682));
    defparam \pid_front.error_p_reg_esr_RNITCC61_18_LC_17_18_0 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_esr_RNITCC61_18_LC_17_18_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_p_reg_esr_RNITCC61_18_LC_17_18_0 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_front.error_p_reg_esr_RNITCC61_18_LC_17_18_0  (
            .in0(N__70206),
            .in1(N__70508),
            .in2(_gnd_net_),
            .in3(N__87545),
            .lcout(\pid_front.error_p_reg_esr_RNITCC61Z0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_prev_esr_18_LC_17_18_1 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_prev_esr_18_LC_17_18_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_prev_esr_18_LC_17_18_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_front.error_d_reg_prev_esr_18_LC_17_18_1  (
            .in0(N__87546),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_d_reg_prevZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87158),
            .ce(N__70472),
            .sr(N__70358));
    defparam \pid_side.error_axb_8_l_ofx_LC_17_18_2 .C_ON=1'b0;
    defparam \pid_side.error_axb_8_l_ofx_LC_17_18_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_axb_8_l_ofx_LC_17_18_2 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \pid_side.error_axb_8_l_ofx_LC_17_18_2  (
            .in0(N__70308),
            .in1(N__74093),
            .in2(_gnd_net_),
            .in3(N__73941),
            .lcout(\pid_side.error_axb_8_l_ofxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_axb_7_LC_17_18_3 .C_ON=1'b0;
    defparam \pid_side.error_axb_7_LC_17_18_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_axb_7_LC_17_18_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \pid_side.error_axb_7_LC_17_18_3  (
            .in0(N__73940),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70307),
            .lcout(\pid_side.error_axbZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNIV6RD_12_LC_17_18_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNIV6RD_12_LC_17_18_4 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNIV6RD_12_LC_17_18_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_RNIV6RD_12_LC_17_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__74092),
            .lcout(drone_H_disp_side_i_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_3_c_RNIIVLQ1_LC_17_18_5 .C_ON=1'b0;
    defparam \pid_side.error_cry_3_c_RNIIVLQ1_LC_17_18_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_3_c_RNIIVLQ1_LC_17_18_5 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \pid_side.error_cry_3_c_RNIIVLQ1_LC_17_18_5  (
            .in0(N__75984),
            .in1(N__75007),
            .in2(_gnd_net_),
            .in3(N__75050),
            .lcout(\pid_side.N_9_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_3_13_LC_17_19_0 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_3_13_LC_17_19_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_3_13_LC_17_19_0 .LUT_INIT=16'b0010000001111111;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_3_13_LC_17_19_0  (
            .in0(N__80791),
            .in1(N__74387),
            .in2(N__80980),
            .in3(N__74844),
            .lcout(\pid_side.N_126 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_5_c_RNI5U9G2_LC_17_19_1 .C_ON=1'b0;
    defparam \pid_side.error_cry_5_c_RNI5U9G2_LC_17_19_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_5_c_RNI5U9G2_LC_17_19_1 .LUT_INIT=16'b0000101001110111;
    LogicCell40 \pid_side.error_cry_5_c_RNI5U9G2_LC_17_19_1  (
            .in0(N__77889),
            .in1(N__74152),
            .in2(N__74575),
            .in3(N__78360),
            .lcout(),
            .ltout(\pid_side.m87_0_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_7_c_RNI06H95_LC_17_19_2 .C_ON=1'b0;
    defparam \pid_side.error_cry_7_c_RNI06H95_LC_17_19_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_7_c_RNI06H95_LC_17_19_2 .LUT_INIT=16'b1010000111110001;
    LogicCell40 \pid_side.error_cry_7_c_RNI06H95_LC_17_19_2  (
            .in0(N__80964),
            .in1(N__74038),
            .in2(N__70278),
            .in3(N__74482),
            .lcout(\pid_side.N_88_0 ),
            .ltout(\pid_side.N_88_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_7_c_RNIQ8TL9_LC_17_19_3 .C_ON=1'b0;
    defparam \pid_side.error_cry_7_c_RNIQ8TL9_LC_17_19_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_7_c_RNIQ8TL9_LC_17_19_3 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \pid_side.error_cry_7_c_RNIQ8TL9_LC_17_19_3  (
            .in0(_gnd_net_),
            .in1(N__80611),
            .in2(N__70275),
            .in3(N__70758),
            .lcout(\pid_side.N_90_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_3_0_c_RNI72GR1_LC_17_19_4 .C_ON=1'b0;
    defparam \pid_side.error_cry_3_0_c_RNI72GR1_LC_17_19_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_3_0_c_RNI72GR1_LC_17_19_4 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \pid_side.error_cry_3_0_c_RNI72GR1_LC_17_19_4  (
            .in0(N__78359),
            .in1(N__74630),
            .in2(_gnd_net_),
            .in3(N__74735),
            .lcout(\pid_side.N_48_1 ),
            .ltout(\pid_side.N_48_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_1_0_c_RNILC344_LC_17_19_5 .C_ON=1'b0;
    defparam \pid_side.error_cry_1_0_c_RNILC344_LC_17_19_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_1_0_c_RNILC344_LC_17_19_5 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \pid_side.error_cry_1_0_c_RNILC344_LC_17_19_5  (
            .in0(N__74664),
            .in1(_gnd_net_),
            .in2(N__70761),
            .in3(N__80963),
            .lcout(\pid_side.N_89_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_0_13_LC_17_19_6 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_0_13_LC_17_19_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_0_13_LC_17_19_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_0_13_LC_17_19_6  (
            .in0(N__80612),
            .in1(N__70752),
            .in2(_gnd_net_),
            .in3(N__70746),
            .lcout(),
            .ltout(\pid_side.N_127_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_13_LC_17_19_7 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_13_LC_17_19_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_esr_13_LC_17_19_7 .LUT_INIT=16'b0011111100001100;
    LogicCell40 \pid_side.error_i_reg_esr_13_LC_17_19_7  (
            .in0(_gnd_net_),
            .in1(N__70740),
            .in2(N__70728),
            .in3(N__70545),
            .lcout(\pid_side.error_i_regZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87172),
            .ce(N__75366),
            .sr(N__79691));
    defparam \pid_side.m153_e_4_LC_17_20_1 .C_ON=1'b0;
    defparam \pid_side.m153_e_4_LC_17_20_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.m153_e_4_LC_17_20_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \pid_side.m153_e_4_LC_17_20_1  (
            .in0(N__70703),
            .in1(N__70675),
            .in2(N__70638),
            .in3(N__77392),
            .lcout(pid_side_m153_e_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_5_13_LC_17_20_3 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_5_13_LC_17_20_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_5_13_LC_17_20_3 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_5_13_LC_17_20_3  (
            .in0(N__75669),
            .in1(N__71509),
            .in2(_gnd_net_),
            .in3(N__70579),
            .lcout(\pid_side.m1_2_03 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_3_0_c_RNIJ9LC4_LC_17_20_4 .C_ON=1'b0;
    defparam \pid_side.error_cry_3_0_c_RNIJ9LC4_LC_17_20_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_3_0_c_RNIJ9LC4_LC_17_20_4 .LUT_INIT=16'b1100000111001101;
    LogicCell40 \pid_side.error_cry_3_0_c_RNIJ9LC4_LC_17_20_4  (
            .in0(N__74750),
            .in1(N__75759),
            .in2(N__78098),
            .in3(N__74656),
            .lcout(\pid_side.N_89_0_1 ),
            .ltout(\pid_side.N_89_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_1_13_LC_17_20_5 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_1_13_LC_17_20_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_1_13_LC_17_20_5 .LUT_INIT=16'b0011111100001100;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_1_13_LC_17_20_5  (
            .in0(_gnd_net_),
            .in1(N__71036),
            .in2(N__70548),
            .in3(N__70815),
            .lcout(\pid_side.error_i_reg_9_rn_2_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_5_c_RNITLN73_LC_17_20_6 .C_ON=1'b0;
    defparam \pid_front.error_cry_5_c_RNITLN73_LC_17_20_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_5_c_RNITLN73_LC_17_20_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \pid_front.error_cry_5_c_RNITLN73_LC_17_20_6  (
            .in0(N__78072),
            .in1(N__72203),
            .in2(_gnd_net_),
            .in3(N__72236),
            .lcout(\pid_front.N_49_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.m70_0_LC_17_21_0 .C_ON=1'b0;
    defparam \pid_front.m70_0_LC_17_21_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.m70_0_LC_17_21_0 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \pid_front.m70_0_LC_17_21_0  (
            .in0(N__76986),
            .in1(N__76299),
            .in2(_gnd_net_),
            .in3(N__76631),
            .lcout(pid_side_N_166_mux),
            .ltout(pid_side_N_166_mux_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_1_15_LC_17_21_1 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_1_15_LC_17_21_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_1_15_LC_17_21_1 .LUT_INIT=16'b1111011111110010;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_1_15_LC_17_21_1  (
            .in0(N__71037),
            .in1(N__76060),
            .in2(N__71040),
            .in3(N__76391),
            .lcout(\pid_front.error_i_reg_esr_RNO_1Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_9_rn_sn_15_LC_17_21_2 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_9_rn_sn_15_LC_17_21_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_9_rn_sn_15_LC_17_21_2 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \pid_front.error_i_reg_9_rn_sn_15_LC_17_21_2  (
            .in0(N__77687),
            .in1(N__76985),
            .in2(_gnd_net_),
            .in3(N__76630),
            .lcout(pid_front_error_i_reg_9_rn_sn_15),
            .ltout(pid_front_error_i_reg_9_rn_sn_15_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_2_15_LC_17_21_3 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_2_15_LC_17_21_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_2_15_LC_17_21_3 .LUT_INIT=16'b0001010100010000;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_2_15_LC_17_21_3  (
            .in0(N__70902),
            .in1(N__76061),
            .in2(N__71025),
            .in3(N__76392),
            .lcout(\pid_front.error_i_reg_esr_RNO_2Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_1_LC_17_21_4 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_1_LC_17_21_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_esr_1_LC_17_21_4 .LUT_INIT=16'b1000000011010000;
    LogicCell40 \pid_front.error_i_reg_esr_1_LC_17_21_4  (
            .in0(N__71548),
            .in1(N__71020),
            .in2(N__70928),
            .in3(N__70868),
            .lcout(\pid_front.error_i_regZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87202),
            .ce(N__72423),
            .sr(N__79698));
    defparam \pid_side.error_i_reg_esr_RNO_4_13_LC_17_21_6 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_4_13_LC_17_21_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_4_13_LC_17_21_6 .LUT_INIT=16'b1000000010001010;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_4_13_LC_17_21_6  (
            .in0(N__76553),
            .in1(N__70821),
            .in2(N__77018),
            .in3(N__75222),
            .lcout(\pid_side.error_i_reg_9_rn_rn_2_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_15_LC_17_22_0 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_15_LC_17_22_0 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_esr_15_LC_17_22_0 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \pid_front.error_i_reg_esr_15_LC_17_22_0  (
            .in0(_gnd_net_),
            .in1(N__70779),
            .in2(N__70809),
            .in3(N__70800),
            .lcout(\pid_front.error_i_regZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87220),
            .ce(N__72417),
            .sr(N__79704));
    defparam \pid_front.error_i_reg_esr_RNO_0_15_LC_17_22_1 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_0_15_LC_17_22_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_0_15_LC_17_22_1 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_0_15_LC_17_22_1  (
            .in0(N__71130),
            .in1(N__71552),
            .in2(_gnd_net_),
            .in3(N__71304),
            .lcout(\pid_front.N_134 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_0_23_LC_17_22_2 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_0_23_LC_17_22_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_0_23_LC_17_22_2 .LUT_INIT=16'b0111111101000000;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_0_23_LC_17_22_2  (
            .in0(N__71305),
            .in1(N__76298),
            .in2(N__71562),
            .in3(N__71131),
            .lcout(),
            .ltout(\pid_front.error_i_reg_esr_RNO_0_0_23_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_23_LC_17_22_3 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_23_LC_17_22_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_esr_23_LC_17_22_3 .LUT_INIT=16'b1100100001000000;
    LogicCell40 \pid_front.error_i_reg_esr_23_LC_17_22_3  (
            .in0(N__77025),
            .in1(N__76557),
            .in2(N__71331),
            .in3(N__76017),
            .lcout(\pid_front.error_i_regZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87220),
            .ce(N__72417),
            .sr(N__79704));
    defparam \pid_front.error_cry_9_c_RNICELJ1_LC_17_22_4 .C_ON=1'b0;
    defparam \pid_front.error_cry_9_c_RNICELJ1_LC_17_22_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_9_c_RNICELJ1_LC_17_22_4 .LUT_INIT=16'b1111010011110111;
    LogicCell40 \pid_front.error_cry_9_c_RNICELJ1_LC_17_22_4  (
            .in0(N__72110),
            .in1(N__78330),
            .in2(N__72061),
            .in3(N__71128),
            .lcout(\pid_front.error_cry_9_c_RNICELJZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_9_c_RNICELJ1_0_LC_17_22_5 .C_ON=1'b0;
    defparam \pid_front.error_cry_9_c_RNICELJ1_0_LC_17_22_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_9_c_RNICELJ1_0_LC_17_22_5 .LUT_INIT=16'b0000000100110001;
    LogicCell40 \pid_front.error_cry_9_c_RNICELJ1_0_LC_17_22_5  (
            .in0(N__71129),
            .in1(N__72050),
            .in2(N__78372),
            .in3(N__72111),
            .lcout(),
            .ltout(\pid_front.error_cry_9_c_RNICELJ1Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_9_c_RNIGTAH4_LC_17_22_6 .C_ON=1'b0;
    defparam \pid_front.error_cry_9_c_RNIGTAH4_LC_17_22_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_9_c_RNIGTAH4_LC_17_22_6 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \pid_front.error_cry_9_c_RNIGTAH4_LC_17_22_6  (
            .in0(_gnd_net_),
            .in1(N__72185),
            .in2(N__71316),
            .in3(N__71313),
            .lcout(\pid_front.N_46_1 ),
            .ltout(\pid_front.N_46_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_1_19_LC_17_22_7 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_1_19_LC_17_22_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_1_19_LC_17_22_7 .LUT_INIT=16'b0000010010001100;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_1_19_LC_17_22_7  (
            .in0(N__80610),
            .in1(N__71265),
            .in2(N__71238),
            .in3(N__76068),
            .lcout(\pid_front.error_i_reg_esr_RNO_1Z0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_esr_3_LC_17_23_7 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_3_LC_17_23_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_3_LC_17_23_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_esr_3_LC_17_23_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__71229),
            .lcout(\pid_front.error_d_regZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87234),
            .ce(N__86329),
            .sr(N__86002));
    defparam \pid_front.error_i_reg_esr_RNO_2_17_LC_17_24_0 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_2_17_LC_17_24_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_2_17_LC_17_24_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_2_17_LC_17_24_0  (
            .in0(N__71874),
            .in1(N__72273),
            .in2(_gnd_net_),
            .in3(N__71188),
            .lcout(),
            .ltout(\pid_front.N_131_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_0_17_LC_17_24_1 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_0_17_LC_17_24_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_0_17_LC_17_24_1 .LUT_INIT=16'b1000101000000010;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_0_17_LC_17_24_1  (
            .in0(N__76605),
            .in1(N__77003),
            .in2(N__71055),
            .in3(N__71052),
            .lcout(),
            .ltout(\pid_front.error_i_reg_9_rn_1_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_17_LC_17_24_2 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_17_LC_17_24_2 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_i_reg_esr_17_LC_17_24_2 .LUT_INIT=16'b0011000011111100;
    LogicCell40 \pid_front.error_i_reg_esr_17_LC_17_24_2  (
            .in0(_gnd_net_),
            .in1(N__72447),
            .in2(N__72438),
            .in3(N__72166),
            .lcout(\pid_front.error_i_regZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87246),
            .ce(N__72418),
            .sr(N__79712));
    defparam \pid_front.error_i_reg_esr_RNO_4_17_LC_17_24_3 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_4_17_LC_17_24_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_4_17_LC_17_24_3 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_4_17_LC_17_24_3  (
            .in0(N__72051),
            .in1(N__78347),
            .in2(N__77779),
            .in3(N__72130),
            .lcout(\pid_front.error_i_reg_esr_RNO_4_0_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_1_0_c_RNI7HHJ3_LC_17_24_4 .C_ON=1'b0;
    defparam \pid_front.error_cry_1_0_c_RNI7HHJ3_LC_17_24_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_1_0_c_RNI7HHJ3_LC_17_24_4 .LUT_INIT=16'b0010010101110101;
    LogicCell40 \pid_front.error_cry_1_0_c_RNI7HHJ3_LC_17_24_4  (
            .in0(N__78071),
            .in1(N__72267),
            .in2(N__77410),
            .in3(N__72237),
            .lcout(),
            .ltout(\pid_front.m89_0_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_5_c_RNIM3P96_LC_17_24_5 .C_ON=1'b0;
    defparam \pid_front.error_cry_5_c_RNIM3P96_LC_17_24_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_5_c_RNIM3P96_LC_17_24_5 .LUT_INIT=16'b0101111000001110;
    LogicCell40 \pid_front.error_cry_5_c_RNIM3P96_LC_17_24_5  (
            .in0(N__77747),
            .in1(N__72210),
            .in2(N__72192),
            .in3(N__72189),
            .lcout(\pid_front.N_90_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_5_17_LC_17_24_6 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_5_17_LC_17_24_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_5_17_LC_17_24_6 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_5_17_LC_17_24_6  (
            .in0(N__72131),
            .in1(N__77743),
            .in2(N__78381),
            .in3(N__72052),
            .lcout(\pid_front.error_i_reg_esr_RNO_5_0_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.state_RNICP2N1_0_LC_18_7_7 .C_ON=1'b0;
    defparam \pid_alt.state_RNICP2N1_0_LC_18_7_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.state_RNICP2N1_0_LC_18_7_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \pid_alt.state_RNICP2N1_0_LC_18_7_7  (
            .in0(_gnd_net_),
            .in1(N__71868),
            .in2(_gnd_net_),
            .in3(N__86151),
            .lcout(\pid_alt.N_939_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_esr_RNIKLMT_10_LC_18_10_2 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_esr_RNIKLMT_10_LC_18_10_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_esr_RNIKLMT_10_LC_18_10_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \pid_side.pid_prereg_esr_RNIKLMT_10_LC_18_10_2  (
            .in0(N__71833),
            .in1(N__71797),
            .in2(N__71767),
            .in3(N__71726),
            .lcout(),
            .ltout(\pid_side.source_pid_1_sqmuxa_1_0_a2_1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_esr_RNIS3LQ1_8_LC_18_10_3 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_esr_RNIS3LQ1_8_LC_18_10_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_esr_RNIS3LQ1_8_LC_18_10_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \pid_side.pid_prereg_esr_RNIS3LQ1_8_LC_18_10_3  (
            .in0(N__71701),
            .in1(N__71662),
            .in2(N__71634),
            .in3(N__71623),
            .lcout(\pid_side.N_99 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_esr_RNI6L23_16_LC_18_10_4 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_esr_RNI6L23_16_LC_18_10_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_esr_RNI6L23_16_LC_18_10_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_side.pid_prereg_esr_RNI6L23_16_LC_18_10_4  (
            .in0(N__72777),
            .in1(N__72768),
            .in2(N__72759),
            .in3(N__72744),
            .lcout(\pid_side.un11lto30_i_a2_3_and ),
            .ltout(\pid_side.un11lto30_i_a2_3_and_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_esr_RNIAEHI_15_LC_18_10_5 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_esr_RNIAEHI_15_LC_18_10_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_esr_RNIAEHI_15_LC_18_10_5 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \pid_side.pid_prereg_esr_RNIAEHI_15_LC_18_10_5  (
            .in0(N__72719),
            .in1(_gnd_net_),
            .in2(N__72699),
            .in3(N__72696),
            .lcout(\pid_side.source_pid_1_sqmuxa_1_0_a2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNISSNM4_12_LC_18_11_3 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNISSNM4_12_LC_18_11_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNISSNM4_12_LC_18_11_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNISSNM4_12_LC_18_11_3  (
            .in0(N__81975),
            .in1(N__83016),
            .in2(_gnd_net_),
            .in3(N__82215),
            .lcout(\pid_side.error_d_reg_prev_esr_RNISSNM4Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_acumm_prereg_esr_RNIOG5R_28_LC_18_11_4 .C_ON=1'b0;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIOG5R_28_LC_18_11_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_acumm_prereg_esr_RNIOG5R_28_LC_18_11_4 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \pid_side.error_i_acumm_prereg_esr_RNIOG5R_28_LC_18_11_4  (
            .in0(N__72654),
            .in1(N__72552),
            .in2(_gnd_net_),
            .in3(N__79935),
            .lcout(\pid_side.error_i_acumm_3_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNI5RKP3_5_LC_18_11_6 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNI5RKP3_5_LC_18_11_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNI5RKP3_5_LC_18_11_6 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_side.error_p_reg_esr_RNI5RKP3_5_LC_18_11_6  (
            .in0(N__78471),
            .in1(N__78552),
            .in2(_gnd_net_),
            .in3(N__78540),
            .lcout(\pid_side.error_p_reg_esr_RNI5RKP3Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIM6H42_0_LC_18_11_7 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIM6H42_0_LC_18_11_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIM6H42_0_LC_18_11_7 .LUT_INIT=16'b0101010110011001;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIM6H42_0_LC_18_11_7  (
            .in0(N__82464),
            .in1(N__82110),
            .in2(N__72489),
            .in3(N__82584),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIM6H42Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNITU3P4_0_10_LC_18_12_0 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNITU3P4_0_10_LC_18_12_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNITU3P4_0_10_LC_18_12_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNITU3P4_0_10_LC_18_12_0  (
            .in0(_gnd_net_),
            .in1(N__78874),
            .in2(_gnd_net_),
            .in3(N__78896),
            .lcout(\pid_side.error_d_reg_prev_esr_RNITU3P4_0Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_9_LC_18_12_1 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_9_LC_18_12_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_9_LC_18_12_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_9_LC_18_12_1  (
            .in0(N__81129),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_d_reg_prevZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87082),
            .ce(N__83400),
            .sr(N__83254));
    defparam \pid_side.error_d_reg_prev_esr_RNI20FI_9_LC_18_12_2 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI20FI_9_LC_18_12_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI20FI_9_LC_18_12_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI20FI_9_LC_18_12_2  (
            .in0(_gnd_net_),
            .in1(N__78441),
            .in2(_gnd_net_),
            .in3(N__81127),
            .lcout(\pid_side.N_2380_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNIKGHS6_10_LC_18_12_3 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIKGHS6_10_LC_18_12_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIKGHS6_10_LC_18_12_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_side.error_p_reg_esr_RNIKGHS6_10_LC_18_12_3  (
            .in0(N__72969),
            .in1(N__72950),
            .in2(N__73002),
            .in3(N__72931),
            .lcout(\pid_side.error_p_reg_esr_RNIKGHS6Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_10_LC_18_12_4 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_10_LC_18_12_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_10_LC_18_12_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_10_LC_18_12_4  (
            .in0(N__81309),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_d_reg_prevZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87082),
            .ce(N__83400),
            .sr(N__83254));
    defparam \pid_side.error_d_reg_prev_esr_RNIIARG_10_LC_18_12_5 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIIARG_10_LC_18_12_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIIARG_10_LC_18_12_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIIARG_10_LC_18_12_5  (
            .in0(_gnd_net_),
            .in1(N__78806),
            .in2(_gnd_net_),
            .in3(N__81308),
            .lcout(),
            .ltout(\pid_side.N_2386_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNIRE1B1_10_LC_18_12_6 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIRE1B1_10_LC_18_12_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIRE1B1_10_LC_18_12_6 .LUT_INIT=16'b0101101010010110;
    LogicCell40 \pid_side.error_p_reg_esr_RNIRE1B1_10_LC_18_12_6  (
            .in0(N__81627),
            .in1(N__78442),
            .in2(N__72972),
            .in3(N__81128),
            .lcout(\pid_side.error_p_reg_esr_RNIRE1B1Z0Z_10 ),
            .ltout(\pid_side.error_p_reg_esr_RNIRE1B1Z0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNIV4S38_10_LC_18_12_7 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIV4S38_10_LC_18_12_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIV4S38_10_LC_18_12_7 .LUT_INIT=16'b1111110011000000;
    LogicCell40 \pid_side.error_p_reg_esr_RNIV4S38_10_LC_18_12_7  (
            .in0(N__72963),
            .in1(N__72951),
            .in2(N__72936),
            .in3(N__72932),
            .lcout(\pid_side.error_p_reg_esr_RNIV4S38Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIT8IL1_22_LC_18_13_0 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIT8IL1_22_LC_18_13_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIT8IL1_22_LC_18_13_0 .LUT_INIT=16'b1110111100001000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIT8IL1_22_LC_18_13_0  (
            .in0(N__84630),
            .in1(N__83550),
            .in2(N__73205),
            .in3(N__72900),
            .lcout(\pid_side.un1_pid_prereg_0_20 ),
            .ltout(\pid_side.un1_pid_prereg_0_20_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIK39M6_22_LC_18_13_1 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIK39M6_22_LC_18_13_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIK39M6_22_LC_18_13_1 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIK39M6_22_LC_18_13_1  (
            .in0(N__72870),
            .in1(N__72855),
            .in2(N__72837),
            .in3(N__72788),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIK39M6Z0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIVBJL1_0_22_LC_18_13_2 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIVBJL1_0_22_LC_18_13_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIVBJL1_0_22_LC_18_13_2 .LUT_INIT=16'b0001100011100111;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIVBJL1_0_22_LC_18_13_2  (
            .in0(N__84631),
            .in1(N__83551),
            .in2(N__73206),
            .in3(N__72827),
            .lcout(\pid_side.un1_pid_prereg_0_21 ),
            .ltout(\pid_side.un1_pid_prereg_0_21_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNISK5B3_22_LC_18_13_3 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNISK5B3_22_LC_18_13_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNISK5B3_22_LC_18_13_3 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNISK5B3_22_LC_18_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__73242),
            .in3(N__73229),
            .lcout(\pid_side.error_d_reg_prev_esr_RNISK5B3Z0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_22_LC_18_13_4 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_22_LC_18_13_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_22_LC_18_13_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_22_LC_18_13_4  (
            .in0(N__84632),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_d_reg_prevZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87096),
            .ce(N__83393),
            .sr(N__83261));
    defparam \pid_side.error_d_reg_prev_esr_RNIVNLO_0_21_LC_18_13_5 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIVNLO_0_21_LC_18_13_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIVNLO_0_21_LC_18_13_5 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIVNLO_0_21_LC_18_13_5  (
            .in0(N__83548),
            .in1(N__73112),
            .in2(_gnd_net_),
            .in3(N__84664),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIVNLO_0Z0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_21_LC_18_13_6 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_21_LC_18_13_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_21_LC_18_13_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_21_LC_18_13_6  (
            .in0(N__84666),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_d_reg_prevZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87096),
            .ce(N__83393),
            .sr(N__83261));
    defparam \pid_side.error_d_reg_prev_esr_RNIVNLO_21_LC_18_13_7 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIVNLO_21_LC_18_13_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIVNLO_21_LC_18_13_7 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIVNLO_21_LC_18_13_7  (
            .in0(N__83549),
            .in1(N__73113),
            .in2(_gnd_net_),
            .in3(N__84665),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIVNLOZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNICOLL9_18_LC_18_14_0 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNICOLL9_18_LC_18_14_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNICOLL9_18_LC_18_14_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNICOLL9_18_LC_18_14_0  (
            .in0(N__73257),
            .in1(N__73513),
            .in2(N__73725),
            .in3(N__73499),
            .lcout(\pid_side.error_d_reg_prev_esr_RNICOLL9Z0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIBG7D2_19_LC_18_14_1 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIBG7D2_19_LC_18_14_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIBG7D2_19_LC_18_14_1 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIBG7D2_19_LC_18_14_1  (
            .in0(N__81653),
            .in1(N__81698),
            .in2(_gnd_net_),
            .in3(N__73289),
            .lcout(\pid_side.un1_pid_prereg_0_10 ),
            .ltout(\pid_side.un1_pid_prereg_0_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIQVAR4_19_LC_18_14_2 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIQVAR4_19_LC_18_14_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIQVAR4_19_LC_18_14_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIQVAR4_19_LC_18_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__73074),
            .in3(N__73514),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIQVAR4Z0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIFF3E2_20_LC_18_14_3 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIFF3E2_20_LC_18_14_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIFF3E2_20_LC_18_14_3 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIFF3E2_20_LC_18_14_3  (
            .in0(N__82965),
            .in1(N__73058),
            .in2(_gnd_net_),
            .in3(N__73043),
            .lcout(\pid_side.un1_pid_prereg_0_12 ),
            .ltout(\pid_side.un1_pid_prereg_0_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIV6JN9_19_LC_18_14_4 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIV6JN9_19_LC_18_14_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIV6JN9_19_LC_18_14_4 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIV6JN9_19_LC_18_14_4  (
            .in0(N__73515),
            .in1(N__73500),
            .in2(N__73491),
            .in3(N__73412),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIV6JN9Z0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI620Q4_15_LC_18_14_5 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI620Q4_15_LC_18_14_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI620Q4_15_LC_18_14_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI620Q4_15_LC_18_14_5  (
            .in0(_gnd_net_),
            .in1(N__73481),
            .in2(_gnd_net_),
            .in3(N__73466),
            .lcout(\pid_side.error_d_reg_prev_esr_RNI620Q4Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI578S4_20_LC_18_14_6 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI578S4_20_LC_18_14_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI578S4_20_LC_18_14_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI578S4_20_LC_18_14_6  (
            .in0(_gnd_net_),
            .in1(N__73430),
            .in2(_gnd_net_),
            .in3(N__73411),
            .lcout(\pid_side.error_d_reg_prev_esr_RNI578S4Z0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI1OK5F_12_LC_18_14_7 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI1OK5F_12_LC_18_14_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI1OK5F_12_LC_18_14_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI1OK5F_12_LC_18_14_7  (
            .in0(N__80115),
            .in1(N__73385),
            .in2(N__80067),
            .in3(N__73372),
            .lcout(\pid_side.error_d_reg_prev_esr_RNI1OK5FZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_1_LC_18_15_2 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_1_LC_18_15_2 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_1_LC_18_15_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_1_LC_18_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__83052),
            .lcout(\pid_side.error_d_reg_prevZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87125),
            .ce(N__83397),
            .sr(N__83219));
    defparam \pid_side.error_d_reg_prev_esr_RNI783D2_18_LC_18_15_3 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI783D2_18_LC_18_15_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI783D2_18_LC_18_15_3 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI783D2_18_LC_18_15_3  (
            .in0(N__81735),
            .in1(N__83093),
            .in2(_gnd_net_),
            .in3(N__73349),
            .lcout(\pid_side.un1_pid_prereg_0_8 ),
            .ltout(\pid_side.un1_pid_prereg_0_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIOVFK9_17_LC_18_15_4 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIOVFK9_17_LC_18_15_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIOVFK9_17_LC_18_15_4 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIOVFK9_17_LC_18_15_4  (
            .in0(N__73326),
            .in1(N__73314),
            .in2(N__73302),
            .in3(N__73253),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIOVFK9Z0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIBG7D2_0_19_LC_18_15_5 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIBG7D2_0_19_LC_18_15_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIBG7D2_0_19_LC_18_15_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIBG7D2_0_19_LC_18_15_5  (
            .in0(N__81657),
            .in1(N__81702),
            .in2(_gnd_net_),
            .in3(N__73285),
            .lcout(\pid_side.un1_pid_prereg_0_9 ),
            .ltout(\pid_side.un1_pid_prereg_0_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIIOAQ4_18_LC_18_15_6 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIIOAQ4_18_LC_18_15_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIIOAQ4_18_LC_18_15_6 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIIOAQ4_18_LC_18_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__73728),
            .in3(N__73721),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIIOAQ4Z0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIQ8P41_0_LC_18_15_7 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIQ8P41_0_LC_18_15_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIQ8P41_0_LC_18_15_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIQ8P41_0_LC_18_15_7  (
            .in0(N__73695),
            .in1(N__82109),
            .in2(_gnd_net_),
            .in3(N__82583),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIQ8P41Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_CH2data_esr_0_LC_18_16_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH2data_esr_0_LC_18_16_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH2data_esr_0_LC_18_16_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH2data_esr_0_LC_18_16_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__83837),
            .lcout(side_command_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87140),
            .ce(N__73929),
            .sr(N__79683));
    defparam \Commands_frame_decoder.source_CH2data_esr_1_LC_18_16_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH2data_esr_1_LC_18_16_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH2data_esr_1_LC_18_16_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH2data_esr_1_LC_18_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84214),
            .lcout(side_command_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87140),
            .ce(N__73929),
            .sr(N__79683));
    defparam \Commands_frame_decoder.source_CH2data_esr_2_LC_18_16_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH2data_esr_2_LC_18_16_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH2data_esr_2_LC_18_16_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Commands_frame_decoder.source_CH2data_esr_2_LC_18_16_2  (
            .in0(N__77586),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(side_command_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87140),
            .ce(N__73929),
            .sr(N__79683));
    defparam \Commands_frame_decoder.source_CH2data_esr_3_LC_18_16_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH2data_esr_3_LC_18_16_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH2data_esr_3_LC_18_16_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH2data_esr_3_LC_18_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84030),
            .lcout(side_command_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87140),
            .ce(N__73929),
            .sr(N__79683));
    defparam \Commands_frame_decoder.source_CH2data_esr_4_LC_18_16_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH2data_esr_4_LC_18_16_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH2data_esr_4_LC_18_16_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH2data_esr_4_LC_18_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85028),
            .lcout(side_command_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87140),
            .ce(N__73929),
            .sr(N__79683));
    defparam \Commands_frame_decoder.source_CH2data_esr_5_LC_18_16_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH2data_esr_5_LC_18_16_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH2data_esr_5_LC_18_16_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH2data_esr_5_LC_18_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85214),
            .lcout(side_command_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87140),
            .ce(N__73929),
            .sr(N__79683));
    defparam \Commands_frame_decoder.source_CH2data_esr_6_LC_18_16_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH2data_esr_6_LC_18_16_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH2data_esr_6_LC_18_16_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH2data_esr_6_LC_18_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73656),
            .lcout(side_command_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87140),
            .ce(N__73929),
            .sr(N__79683));
    defparam \Commands_frame_decoder.source_CH2data_ess_7_LC_18_16_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH2data_ess_7_LC_18_16_7 .SEQ_MODE=4'b1001;
    defparam \Commands_frame_decoder.source_CH2data_ess_7_LC_18_16_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Commands_frame_decoder.source_CH2data_ess_7_LC_18_16_7  (
            .in0(N__85396),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(side_command_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87140),
            .ce(N__73929),
            .sr(N__79683));
    defparam \pid_side.error_cry_0_c_inv_LC_18_17_0 .C_ON=1'b1;
    defparam \pid_side.error_cry_0_c_inv_LC_18_17_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_0_c_inv_LC_18_17_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_side.error_cry_0_c_inv_LC_18_17_0  (
            .in0(_gnd_net_),
            .in1(N__73902),
            .in2(_gnd_net_),
            .in3(N__73911),
            .lcout(\pid_side.error_axb_0 ),
            .ltout(),
            .carryin(bfn_18_17_0_),
            .carryout(\pid_side.error_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_0_c_RNI43F5_LC_18_17_1 .C_ON=1'b1;
    defparam \pid_side.error_cry_0_c_RNI43F5_LC_18_17_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_0_c_RNI43F5_LC_18_17_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_side.error_cry_0_c_RNI43F5_LC_18_17_1  (
            .in0(_gnd_net_),
            .in1(N__73896),
            .in2(_gnd_net_),
            .in3(N__73818),
            .lcout(\pid_side.error_1 ),
            .ltout(),
            .carryin(\pid_side.error_cry_0 ),
            .carryout(\pid_side.error_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_1_c_RNI66G5_LC_18_17_2 .C_ON=1'b1;
    defparam \pid_side.error_cry_1_c_RNI66G5_LC_18_17_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_1_c_RNI66G5_LC_18_17_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_side.error_cry_1_c_RNI66G5_LC_18_17_2  (
            .in0(_gnd_net_),
            .in1(N__73815),
            .in2(_gnd_net_),
            .in3(N__73806),
            .lcout(\pid_side.error_2 ),
            .ltout(),
            .carryin(\pid_side.error_cry_1 ),
            .carryout(\pid_side.error_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_2_c_RNI89H5_LC_18_17_3 .C_ON=1'b1;
    defparam \pid_side.error_cry_2_c_RNI89H5_LC_18_17_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_2_c_RNI89H5_LC_18_17_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_side.error_cry_2_c_RNI89H5_LC_18_17_3  (
            .in0(_gnd_net_),
            .in1(N__73803),
            .in2(_gnd_net_),
            .in3(N__73794),
            .lcout(\pid_side.error_3 ),
            .ltout(),
            .carryin(\pid_side.error_cry_2 ),
            .carryout(\pid_side.error_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_3_c_RNI1SDJ_LC_18_17_4 .C_ON=1'b1;
    defparam \pid_side.error_cry_3_c_RNI1SDJ_LC_18_17_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_3_c_RNI1SDJ_LC_18_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_cry_3_c_RNI1SDJ_LC_18_17_4  (
            .in0(_gnd_net_),
            .in1(N__73791),
            .in2(N__73782),
            .in3(N__73773),
            .lcout(\pid_side.error_4 ),
            .ltout(),
            .carryin(\pid_side.error_cry_3 ),
            .carryout(\pid_side.error_cry_0_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_0_0_c_RNIF3ET_LC_18_17_5 .C_ON=1'b1;
    defparam \pid_side.error_cry_0_0_c_RNIF3ET_LC_18_17_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_0_0_c_RNIF3ET_LC_18_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_cry_0_0_c_RNIF3ET_LC_18_17_5  (
            .in0(_gnd_net_),
            .in1(N__73770),
            .in2(N__73761),
            .in3(N__73752),
            .lcout(\pid_side.error_5 ),
            .ltout(),
            .carryin(\pid_side.error_cry_0_0 ),
            .carryout(\pid_side.error_cry_1_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_1_0_c_RNII9K11_LC_18_17_6 .C_ON=1'b1;
    defparam \pid_side.error_cry_1_0_c_RNII9K11_LC_18_17_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_1_0_c_RNII9K11_LC_18_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_cry_1_0_c_RNII9K11_LC_18_17_6  (
            .in0(_gnd_net_),
            .in1(N__73749),
            .in2(N__73743),
            .in3(N__73731),
            .lcout(\pid_side.error_6 ),
            .ltout(),
            .carryin(\pid_side.error_cry_1_0 ),
            .carryout(\pid_side.error_cry_2_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_2_0_c_RNILFQL_LC_18_17_7 .C_ON=1'b1;
    defparam \pid_side.error_cry_2_0_c_RNILFQL_LC_18_17_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_2_0_c_RNILFQL_LC_18_17_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_cry_2_0_c_RNILFQL_LC_18_17_7  (
            .in0(_gnd_net_),
            .in1(N__74310),
            .in2(N__74304),
            .in3(N__74292),
            .lcout(\pid_side.error_7 ),
            .ltout(),
            .carryin(\pid_side.error_cry_2_0 ),
            .carryout(\pid_side.error_cry_3_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_3_0_c_RNIOL0Q_LC_18_18_0 .C_ON=1'b1;
    defparam \pid_side.error_cry_3_0_c_RNIOL0Q_LC_18_18_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_3_0_c_RNIOL0Q_LC_18_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_cry_3_0_c_RNIOL0Q_LC_18_18_0  (
            .in0(_gnd_net_),
            .in1(N__74289),
            .in2(N__74274),
            .in3(N__74262),
            .lcout(\pid_side.error_8 ),
            .ltout(),
            .carryin(bfn_18_18_0_),
            .carryout(\pid_side.error_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_4_c_RNIC8FJ_LC_18_18_1 .C_ON=1'b1;
    defparam \pid_side.error_cry_4_c_RNIC8FJ_LC_18_18_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_4_c_RNIC8FJ_LC_18_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_cry_4_c_RNIC8FJ_LC_18_18_1  (
            .in0(_gnd_net_),
            .in1(N__74259),
            .in2(N__74244),
            .in3(N__74232),
            .lcout(\pid_side.error_9 ),
            .ltout(),
            .carryin(\pid_side.error_cry_4 ),
            .carryout(\pid_side.error_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_5_c_RNIM4IS_LC_18_18_2 .C_ON=1'b1;
    defparam \pid_side.error_cry_5_c_RNIM4IS_LC_18_18_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_5_c_RNIM4IS_LC_18_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_cry_5_c_RNIM4IS_LC_18_18_2  (
            .in0(_gnd_net_),
            .in1(N__74229),
            .in2(N__74214),
            .in3(N__74202),
            .lcout(\pid_side.error_10 ),
            .ltout(),
            .carryin(\pid_side.error_cry_5 ),
            .carryout(\pid_side.error_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_6_c_RNIQBMT_LC_18_18_3 .C_ON=1'b1;
    defparam \pid_side.error_cry_6_c_RNIQBMT_LC_18_18_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_6_c_RNIQBMT_LC_18_18_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_side.error_cry_6_c_RNIQBMT_LC_18_18_3  (
            .in0(_gnd_net_),
            .in1(N__74199),
            .in2(_gnd_net_),
            .in3(N__74109),
            .lcout(\pid_side.error_11 ),
            .ltout(),
            .carryin(\pid_side.error_cry_6 ),
            .carryout(\pid_side.error_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_7_c_RNIPRDP1_LC_18_18_4 .C_ON=1'b1;
    defparam \pid_side.error_cry_7_c_RNIPRDP1_LC_18_18_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_7_c_RNIPRDP1_LC_18_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_cry_7_c_RNIPRDP1_LC_18_18_4  (
            .in0(_gnd_net_),
            .in1(N__74106),
            .in2(N__74100),
            .in3(N__73989),
            .lcout(\pid_side.error_12 ),
            .ltout(),
            .carryin(\pid_side.error_cry_7 ),
            .carryout(\pid_side.error_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_8_c_RNIUUKS_LC_18_18_5 .C_ON=1'b1;
    defparam \pid_side.error_cry_8_c_RNIUUKS_LC_18_18_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_8_c_RNIUUKS_LC_18_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_cry_8_c_RNIUUKS_LC_18_18_5  (
            .in0(_gnd_net_),
            .in1(N__73986),
            .in2(N__73980),
            .in3(N__73956),
            .lcout(\pid_side.error_13 ),
            .ltout(),
            .carryin(\pid_side.error_cry_8 ),
            .carryout(\pid_side.error_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_9_c_RNI13MS_LC_18_18_6 .C_ON=1'b1;
    defparam \pid_side.error_cry_9_c_RNI13MS_LC_18_18_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_9_c_RNI13MS_LC_18_18_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_cry_9_c_RNI13MS_LC_18_18_6  (
            .in0(_gnd_net_),
            .in1(N__73953),
            .in2(N__74949),
            .in3(N__73944),
            .lcout(\pid_side.error_14 ),
            .ltout(),
            .carryin(\pid_side.error_cry_9 ),
            .carryout(\pid_side.error_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_10_c_RNIBCT11_LC_18_18_7 .C_ON=1'b0;
    defparam \pid_side.error_cry_10_c_RNIBCT11_LC_18_18_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_10_c_RNIBCT11_LC_18_18_7 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_side.error_cry_10_c_RNIBCT11_LC_18_18_7  (
            .in0(N__74958),
            .in1(N__74948),
            .in2(_gnd_net_),
            .in3(N__74934),
            .lcout(\pid_side.error_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_1_0_c_RNI9P812_LC_18_19_0 .C_ON=1'b0;
    defparam \pid_side.error_cry_1_0_c_RNI9P812_LC_18_19_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_1_0_c_RNI9P812_LC_18_19_0 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \pid_side.error_cry_1_0_c_RNI9P812_LC_18_19_0  (
            .in0(N__75968),
            .in1(N__75879),
            .in2(_gnd_net_),
            .in3(N__75821),
            .lcout(\pid_side.N_51_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_3_0_c_RNIL6HL1_LC_18_19_1 .C_ON=1'b0;
    defparam \pid_side.error_cry_3_0_c_RNIL6HL1_LC_18_19_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_3_0_c_RNIL6HL1_LC_18_19_1 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \pid_side.error_cry_3_0_c_RNIL6HL1_LC_18_19_1  (
            .in0(N__78209),
            .in1(N__74734),
            .in2(_gnd_net_),
            .in3(N__74628),
            .lcout(\pid_side.N_48_1_0 ),
            .ltout(\pid_side.N_48_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_10_21_LC_18_19_2 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_10_21_LC_18_19_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_10_21_LC_18_19_2 .LUT_INIT=16'b1111111010111010;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_10_21_LC_18_19_2  (
            .in0(N__77698),
            .in1(N__78041),
            .in2(N__74703),
            .in3(N__74699),
            .lcout(\pid_side.error_i_reg_esr_RNO_10Z0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_9_21_LC_18_19_3 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_9_21_LC_18_19_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_9_21_LC_18_19_3 .LUT_INIT=16'b0010001100100000;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_9_21_LC_18_19_3  (
            .in0(N__74700),
            .in1(N__77699),
            .in2(N__78085),
            .in3(N__74691),
            .lcout(),
            .ltout(\pid_side.error_i_reg_esr_RNO_9Z0Z_21_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_5_21_LC_18_19_4 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_5_21_LC_18_19_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_5_21_LC_18_19_4 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_5_21_LC_18_19_4  (
            .in0(_gnd_net_),
            .in1(N__74964),
            .in2(N__74685),
            .in3(N__74682),
            .lcout(\pid_side.N_116_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_1_0_c_RNIATE52_LC_18_19_5 .C_ON=1'b0;
    defparam \pid_side.error_cry_1_0_c_RNIATE52_LC_18_19_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_1_0_c_RNIATE52_LC_18_19_5 .LUT_INIT=16'b0000111101010101;
    LogicCell40 \pid_side.error_cry_1_0_c_RNIATE52_LC_18_19_5  (
            .in0(N__75822),
            .in1(_gnd_net_),
            .in2(N__75896),
            .in3(N__78334),
            .lcout(\pid_side.N_51_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_6_20_LC_18_19_6 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_6_20_LC_18_19_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_6_20_LC_18_19_6 .LUT_INIT=16'b0100001101001111;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_6_20_LC_18_19_6  (
            .in0(N__74629),
            .in1(N__77401),
            .in2(N__78373),
            .in3(N__74557),
            .lcout(),
            .ltout(\pid_side.G_5_0_m4_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_3_20_LC_18_19_7 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_3_20_LC_18_19_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_3_20_LC_18_19_7 .LUT_INIT=16'b0101111000001110;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_3_20_LC_18_19_7  (
            .in0(N__77402),
            .in1(N__74480),
            .in2(N__74424),
            .in3(N__74383),
            .lcout(\pid_side.N_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_1_0_c_RNIC27G2_LC_18_20_0 .C_ON=1'b0;
    defparam \pid_side.error_cry_1_0_c_RNIC27G2_LC_18_20_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_1_0_c_RNIC27G2_LC_18_20_0 .LUT_INIT=16'b0010010101110101;
    LogicCell40 \pid_side.error_cry_1_0_c_RNIC27G2_LC_18_20_0  (
            .in0(N__75964),
            .in1(N__75883),
            .in2(N__78084),
            .in3(N__75823),
            .lcout(\pid_side.g0_7_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_5_LC_18_20_2 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_5_LC_18_20_2 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_i_reg_esr_5_LC_18_20_2 .LUT_INIT=16'b1000000011010000;
    LogicCell40 \pid_side.error_i_reg_esr_5_LC_18_20_2  (
            .in0(N__75740),
            .in1(N__75546),
            .in2(N__75528),
            .in3(N__75207),
            .lcout(\pid_side.error_i_regZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87203),
            .ce(N__75367),
            .sr(N__79699));
    defparam \pid_side.error_cry_1_c_RNIJOP31_LC_18_20_3 .C_ON=1'b0;
    defparam \pid_side.error_cry_1_c_RNIJOP31_LC_18_20_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_1_c_RNIJOP31_LC_18_20_3 .LUT_INIT=16'b0010010101110101;
    LogicCell40 \pid_side.error_cry_1_c_RNIJOP31_LC_18_20_3  (
            .in0(N__75962),
            .in1(N__75118),
            .in2(N__78083),
            .in3(N__75184),
            .lcout(),
            .ltout(\pid_side.g0_6_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_3_c_RNI61K33_LC_18_20_4 .C_ON=1'b0;
    defparam \pid_side.error_cry_3_c_RNI61K33_LC_18_20_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_3_c_RNI61K33_LC_18_20_4 .LUT_INIT=16'b1010000111110001;
    LogicCell40 \pid_side.error_cry_3_c_RNI61K33_LC_18_20_4  (
            .in0(N__78039),
            .in1(N__75015),
            .in2(N__75225),
            .in3(N__75068),
            .lcout(\pid_side.N_12_1_1 ),
            .ltout(\pid_side.N_12_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_0_5_LC_18_20_5 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_0_5_LC_18_20_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_0_5_LC_18_20_5 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_0_5_LC_18_20_5  (
            .in0(_gnd_net_),
            .in1(N__77704),
            .in2(N__75216),
            .in3(N__75213),
            .lcout(\pid_side.N_116_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_12_21_LC_18_20_6 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_12_21_LC_18_20_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_12_21_LC_18_20_6 .LUT_INIT=16'b0000110001110111;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_12_21_LC_18_20_6  (
            .in0(N__75185),
            .in1(N__78035),
            .in2(N__75130),
            .in3(N__75963),
            .lcout(),
            .ltout(\pid_side.g0_10_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_8_21_LC_18_20_7 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_8_21_LC_18_20_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_8_21_LC_18_20_7 .LUT_INIT=16'b1111000001010011;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_8_21_LC_18_20_7  (
            .in0(N__75069),
            .in1(N__75014),
            .in2(N__74967),
            .in3(N__78040),
            .lcout(\pid_side.N_12_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_3_23_LC_18_21_0 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_3_23_LC_18_21_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_3_23_LC_18_21_0 .LUT_INIT=16'b1111001000000010;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_3_23_LC_18_21_0  (
            .in0(N__77703),
            .in1(N__76097),
            .in2(N__76310),
            .in3(N__76337),
            .lcout(\pid_front.error_i_reg_esr_RNO_3Z0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_0_c_RNIVSLV_LC_18_21_1 .C_ON=1'b0;
    defparam \pid_front.error_cry_0_c_RNIVSLV_LC_18_21_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_0_c_RNIVSLV_LC_18_21_1 .LUT_INIT=16'b0010010101110101;
    LogicCell40 \pid_front.error_cry_0_c_RNIVSLV_LC_18_21_1  (
            .in0(N__78166),
            .in1(N__77258),
            .in2(N__77849),
            .in3(N__77175),
            .lcout(),
            .ltout(\pid_front.m14_0_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_1_c_RNI0UV52_LC_18_21_2 .C_ON=1'b0;
    defparam \pid_front.error_cry_1_c_RNI0UV52_LC_18_21_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_1_c_RNI0UV52_LC_18_21_2 .LUT_INIT=16'b1010000111110001;
    LogicCell40 \pid_front.error_cry_1_c_RNI0UV52_LC_18_21_2  (
            .in0(N__77947),
            .in1(N__77125),
            .in2(N__77094),
            .in3(N__77071),
            .lcout(\pid_front.N_15_1 ),
            .ltout(\pid_front.N_15_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_1_c_RNI9B9J2_LC_18_21_3 .C_ON=1'b0;
    defparam \pid_front.error_cry_1_c_RNI9B9J2_LC_18_21_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_1_c_RNI9B9J2_LC_18_21_3 .LUT_INIT=16'b0000000000000101;
    LogicCell40 \pid_front.error_cry_1_c_RNI9B9J2_LC_18_21_3  (
            .in0(N__77682),
            .in1(_gnd_net_),
            .in2(N__77034),
            .in3(N__80304),
            .lcout(),
            .ltout(\pid_front.m3_2_03_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_1_c_RNISFH18_LC_18_21_4 .C_ON=1'b0;
    defparam \pid_front.error_cry_1_c_RNISFH18_LC_18_21_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_1_c_RNISFH18_LC_18_21_4 .LUT_INIT=16'b1000000011000100;
    LogicCell40 \pid_front.error_cry_1_c_RNISFH18_LC_18_21_4  (
            .in0(N__76990),
            .in1(N__76629),
            .in2(N__76395),
            .in3(N__76096),
            .lcout(\pid_front.error_i_reg_9_rn_rn_2_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_1_c_RNI4G2A2_LC_18_21_5 .C_ON=1'b0;
    defparam \pid_front.error_cry_1_c_RNI4G2A2_LC_18_21_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_1_c_RNI4G2A2_LC_18_21_5 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \pid_front.error_cry_1_c_RNI4G2A2_LC_18_21_5  (
            .in0(N__77681),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__76362),
            .lcout(\pid_front.N_104 ),
            .ltout(\pid_front.N_104_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_2_23_LC_18_21_6 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_2_23_LC_18_21_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_2_23_LC_18_21_6 .LUT_INIT=16'b1011000111110101;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_2_23_LC_18_21_6  (
            .in0(N__76286),
            .in1(N__77683),
            .in2(N__76101),
            .in3(N__76098),
            .lcout(),
            .ltout(\pid_front.error_i_reg_esr_RNO_2Z0Z_23_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_i_reg_esr_RNO_1_23_LC_18_21_7 .C_ON=1'b0;
    defparam \pid_front.error_i_reg_esr_RNO_1_23_LC_18_21_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_i_reg_esr_RNO_1_23_LC_18_21_7 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \pid_front.error_i_reg_esr_RNO_1_23_LC_18_21_7  (
            .in0(_gnd_net_),
            .in1(N__76062),
            .in2(N__76026),
            .in3(N__76023),
            .lcout(\pid_front.error_i_reg_esr_RNO_1_0_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_xy_ki_0_rep1_esr_LC_18_22_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_ki_0_rep1_esr_LC_18_22_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_ki_0_rep1_esr_LC_18_22_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_xy_ki_0_rep1_esr_LC_18_22_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__83848),
            .lcout(xy_ki_0_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87235),
            .ce(N__78711),
            .sr(N__79709));
    defparam \Commands_frame_decoder.source_xy_ki_0_rep2_esr_LC_18_22_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_ki_0_rep2_esr_LC_18_22_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_ki_0_rep2_esr_LC_18_22_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Commands_frame_decoder.source_xy_ki_0_rep2_esr_LC_18_22_1  (
            .in0(N__83849),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(xy_ki_0_rep2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87235),
            .ce(N__78711),
            .sr(N__79709));
    defparam \Commands_frame_decoder.source_xy_ki_fast_esr_0_LC_18_22_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_ki_fast_esr_0_LC_18_22_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_ki_fast_esr_0_LC_18_22_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_xy_ki_fast_esr_0_LC_18_22_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__83850),
            .lcout(xy_ki_fast_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87235),
            .ce(N__78711),
            .sr(N__79709));
    defparam \Commands_frame_decoder.source_xy_ki_1_rep1_esr_LC_18_22_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_ki_1_rep1_esr_LC_18_22_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_ki_1_rep1_esr_LC_18_22_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_xy_ki_1_rep1_esr_LC_18_22_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84221),
            .lcout(xy_ki_1_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87235),
            .ce(N__78711),
            .sr(N__79709));
    defparam \Commands_frame_decoder.source_xy_ki_fast_esr_1_LC_18_22_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_ki_fast_esr_1_LC_18_22_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_ki_fast_esr_1_LC_18_22_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Commands_frame_decoder.source_xy_ki_fast_esr_1_LC_18_22_4  (
            .in0(N__84222),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(xy_ki_fast_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87235),
            .ce(N__78711),
            .sr(N__79709));
    defparam \Commands_frame_decoder.source_xy_ki_2_rep1_esr_LC_18_22_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_ki_2_rep1_esr_LC_18_22_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_ki_2_rep1_esr_LC_18_22_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Commands_frame_decoder.source_xy_ki_2_rep1_esr_LC_18_22_5  (
            .in0(N__77572),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(xy_ki_2_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87235),
            .ce(N__78711),
            .sr(N__79709));
    defparam \Commands_frame_decoder.source_xy_ki_fast_esr_2_LC_18_22_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_ki_fast_esr_2_LC_18_22_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_ki_fast_esr_2_LC_18_22_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_xy_ki_fast_esr_2_LC_18_22_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__77571),
            .lcout(xy_ki_fast_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87235),
            .ce(N__78711),
            .sr(N__79709));
    defparam \Commands_frame_decoder.source_xy_ki_3_rep1_esr_LC_18_22_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_ki_3_rep1_esr_LC_18_22_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_ki_3_rep1_esr_LC_18_22_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_xy_ki_3_rep1_esr_LC_18_22_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84000),
            .lcout(xy_ki_3_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87235),
            .ce(N__78711),
            .sr(N__79709));
    defparam \pid_side.error_p_reg_esr_6_LC_20_10_4 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_6_LC_20_10_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_6_LC_20_10_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_p_reg_esr_6_LC_20_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__77292),
            .lcout(\pid_side.error_p_regZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87084),
            .ce(N__85746),
            .sr(N__86019));
    defparam \pid_side.error_p_reg_esr_RNIG7MC2_0_5_LC_20_11_0 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIG7MC2_0_5_LC_20_11_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIG7MC2_0_5_LC_20_11_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_side.error_p_reg_esr_RNIG7MC2_0_5_LC_20_11_0  (
            .in0(_gnd_net_),
            .in1(N__78485),
            .in2(_gnd_net_),
            .in3(N__78510),
            .lcout(\pid_side.error_p_reg_esr_RNIG7MC2_0Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNI76TK1_0_5_LC_20_11_1 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNI76TK1_0_5_LC_20_11_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNI76TK1_0_5_LC_20_11_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \pid_side.error_p_reg_esr_RNI76TK1_0_5_LC_20_11_1  (
            .in0(N__78611),
            .in1(N__81366),
            .in2(N__80127),
            .in3(N__78621),
            .lcout(\pid_side.error_p_reg_esr_RNI76TK1_0Z0Z_5 ),
            .ltout(\pid_side.error_p_reg_esr_RNI76TK1_0Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNIG7MC2_5_LC_20_11_2 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIG7MC2_5_LC_20_11_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIG7MC2_5_LC_20_11_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \pid_side.error_p_reg_esr_RNIG7MC2_5_LC_20_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__78636),
            .in3(N__78511),
            .lcout(\pid_side.error_p_reg_esr_RNIG7MC2Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNIIHEQ_4_LC_20_11_3 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIIHEQ_4_LC_20_11_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIIHEQ_4_LC_20_11_3 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_side.error_p_reg_esr_RNIIHEQ_4_LC_20_11_3  (
            .in0(N__81563),
            .in1(N__81548),
            .in2(_gnd_net_),
            .in3(N__81524),
            .lcout(\pid_side.error_p_reg_esr_RNIIHEQZ0Z_4 ),
            .ltout(\pid_side.error_p_reg_esr_RNIIHEQZ0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNI76TK1_5_LC_20_11_4 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNI76TK1_5_LC_20_11_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNI76TK1_5_LC_20_11_4 .LUT_INIT=16'b1101010011101000;
    LogicCell40 \pid_side.error_p_reg_esr_RNI76TK1_5_LC_20_11_4  (
            .in0(N__81367),
            .in1(N__80126),
            .in2(N__78615),
            .in3(N__78612),
            .lcout(\pid_side.error_p_reg_esr_RNI76TK1Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNIIFTC1_0_6_LC_20_11_5 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIIFTC1_0_6_LC_20_11_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIIFTC1_0_6_LC_20_11_5 .LUT_INIT=16'b0010110111010010;
    LogicCell40 \pid_side.error_p_reg_esr_RNIIFTC1_0_6_LC_20_11_5  (
            .in0(N__78610),
            .in1(N__81365),
            .in2(N__78584),
            .in3(N__78567),
            .lcout(\pid_side.error_p_reg_esr_RNIIFTC1_0Z0Z_6 ),
            .ltout(\pid_side.error_p_reg_esr_RNIIFTC1_0Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNIUKN42_6_LC_20_11_6 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIUKN42_6_LC_20_11_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIUKN42_6_LC_20_11_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \pid_side.error_p_reg_esr_RNIUKN42_6_LC_20_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__78543),
            .in3(N__78539),
            .lcout(),
            .ltout(\pid_side.un1_pid_prereg_66_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNIL2B66_5_LC_20_11_7 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIL2B66_5_LC_20_11_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIL2B66_5_LC_20_11_7 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \pid_side.error_p_reg_esr_RNIL2B66_5_LC_20_11_7  (
            .in0(N__78512),
            .in1(N__78486),
            .in2(N__78474),
            .in3(N__78467),
            .lcout(\pid_side.error_p_reg_esr_RNIL2B66Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNI4O091_10_LC_20_12_0 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNI4O091_10_LC_20_12_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNI4O091_10_LC_20_12_0 .LUT_INIT=16'b1110111110001100;
    LogicCell40 \pid_side.error_p_reg_esr_RNI4O091_10_LC_20_12_0  (
            .in0(N__81118),
            .in1(N__81619),
            .in2(N__78447),
            .in3(N__81299),
            .lcout(\pid_side.error_p_reg_esr_RNI4O091Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNI4O091_0_10_LC_20_12_1 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNI4O091_0_10_LC_20_12_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNI4O091_0_10_LC_20_12_1 .LUT_INIT=16'b1111010101110001;
    LogicCell40 \pid_side.error_p_reg_esr_RNI4O091_0_10_LC_20_12_1  (
            .in0(N__81300),
            .in1(N__78446),
            .in2(N__81626),
            .in3(N__81119),
            .lcout(),
            .ltout(\pid_side.error_p_reg_esr_RNI4O091_0Z0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIV62K2_10_LC_20_12_2 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIV62K2_10_LC_20_12_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIV62K2_10_LC_20_12_2 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIV62K2_10_LC_20_12_2  (
            .in0(N__78814),
            .in1(_gnd_net_),
            .in2(N__78915),
            .in3(N__78912),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIV62K2Z0Z_10 ),
            .ltout(\pid_side.error_d_reg_prev_esr_RNIV62K2Z0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNID3GT3_0_10_LC_20_12_3 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNID3GT3_0_10_LC_20_12_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNID3GT3_0_10_LC_20_12_3 .LUT_INIT=16'b1011010001001011;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNID3GT3_0_10_LC_20_12_3  (
            .in0(N__81301),
            .in1(N__78815),
            .in2(N__78906),
            .in3(N__81671),
            .lcout(\pid_side.error_d_reg_prev_esr_RNID3GT3_0Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNI80KL2_12_LC_20_12_4 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNI80KL2_12_LC_20_12_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNI80KL2_12_LC_20_12_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \pid_side.error_p_reg_esr_RNI80KL2_12_LC_20_12_4  (
            .in0(N__81842),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78781),
            .lcout(),
            .ltout(\pid_side.un1_pid_prereg_153_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNII28CB_10_LC_20_12_5 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNII28CB_10_LC_20_12_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNII28CB_10_LC_20_12_5 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNII28CB_10_LC_20_12_5  (
            .in0(N__78895),
            .in1(N__78876),
            .in2(N__78831),
            .in3(N__78789),
            .lcout(\pid_side.error_d_reg_prev_esr_RNII28CBZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNID3GT3_10_LC_20_12_6 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNID3GT3_10_LC_20_12_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNID3GT3_10_LC_20_12_6 .LUT_INIT=16'b1110111110001010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNID3GT3_10_LC_20_12_6  (
            .in0(N__81672),
            .in1(N__81302),
            .in2(N__78819),
            .in3(N__78795),
            .lcout(\pid_side.error_d_reg_prev_esr_RNID3GT3Z0Z_10 ),
            .ltout(\pid_side.error_d_reg_prev_esr_RNID3GT3Z0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIH0S9B_10_LC_20_12_7 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIH0S9B_10_LC_20_12_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIH0S9B_10_LC_20_12_7 .LUT_INIT=16'b1111101010100000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIH0S9B_10_LC_20_12_7  (
            .in0(N__78782),
            .in1(N__78759),
            .in2(N__78741),
            .in3(N__81843),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIH0S9BZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_esr_4_LC_20_13_1 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_4_LC_20_13_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_4_LC_20_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_esr_4_LC_20_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__78726),
            .lcout(\pid_side.error_d_regZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87127),
            .ce(N__85723),
            .sr(N__86012));
    defparam \Commands_frame_decoder.source_xy_ki_1_rep2_esr_LC_20_14_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_ki_1_rep2_esr_LC_20_14_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_ki_1_rep2_esr_LC_20_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_xy_ki_1_rep2_esr_LC_20_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84208),
            .lcout(xy_ki_1_rep2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87142),
            .ce(N__78710),
            .sr(N__79684));
    defparam \pid_side.error_d_reg_prev_esr_RNI5RIO_0_14_LC_20_15_0 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI5RIO_0_14_LC_20_15_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI5RIO_0_14_LC_20_15_0 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI5RIO_0_14_LC_20_15_0  (
            .in0(N__84456),
            .in1(N__84252),
            .in2(_gnd_net_),
            .in3(N__85809),
            .lcout(\pid_side.error_d_reg_prev_esr_RNI5RIO_0Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_14_LC_20_15_1 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_14_LC_20_15_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_14_LC_20_15_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_14_LC_20_15_1  (
            .in0(N__85811),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_d_reg_prevZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87160),
            .ce(N__83402),
            .sr(N__83228));
    defparam \pid_side.error_d_reg_prev_esr_RNI5RIO_14_LC_20_15_2 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI5RIO_14_LC_20_15_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI5RIO_14_LC_20_15_2 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI5RIO_14_LC_20_15_2  (
            .in0(N__84457),
            .in1(N__84253),
            .in2(_gnd_net_),
            .in3(N__85810),
            .lcout(\pid_side.error_d_reg_prev_esr_RNI5RIOZ0Z_14 ),
            .ltout(\pid_side.error_d_reg_prev_esr_RNI5RIOZ0Z_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI73UC2_0_14_LC_20_15_3 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI73UC2_0_14_LC_20_15_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI73UC2_0_14_LC_20_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI73UC2_0_14_LC_20_15_3  (
            .in0(_gnd_net_),
            .in1(N__78959),
            .in2(N__78993),
            .in3(N__78989),
            .lcout(\pid_side.error_d_reg_prev_esr_RNI73UC2_0Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI8UIO_0_15_LC_20_15_4 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI8UIO_0_15_LC_20_15_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI8UIO_0_15_LC_20_15_4 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI8UIO_0_15_LC_20_15_4  (
            .in0(N__84329),
            .in1(N__78947),
            .in2(_gnd_net_),
            .in3(N__82297),
            .lcout(\pid_side.error_d_reg_prev_esr_RNI8UIO_0Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_15_LC_20_15_5 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_15_LC_20_15_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_15_LC_20_15_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_15_LC_20_15_5  (
            .in0(N__82299),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_d_reg_prevZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87160),
            .ce(N__83402),
            .sr(N__83228));
    defparam \pid_side.error_d_reg_prev_esr_RNI8UIO_15_LC_20_15_6 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI8UIO_15_LC_20_15_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI8UIO_15_LC_20_15_6 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI8UIO_15_LC_20_15_6  (
            .in0(N__84330),
            .in1(N__78948),
            .in2(_gnd_net_),
            .in3(N__82298),
            .lcout(\pid_side.error_d_reg_prev_esr_RNI8UIOZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_fast_esr_RNIPEC11_12_LC_20_16_0 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_fast_esr_RNIPEC11_12_LC_20_16_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_fast_esr_RNIPEC11_12_LC_20_16_0 .LUT_INIT=16'b1111011001100000;
    LogicCell40 \pid_side.error_d_reg_fast_esr_RNIPEC11_12_LC_20_16_0  (
            .in0(N__81900),
            .in1(N__81864),
            .in2(N__84807),
            .in3(N__82051),
            .lcout(\pid_side.error_d_reg_fast_esr_RNIPEC11Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_fast_esr_RNIPHKN_12_LC_20_16_1 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_fast_esr_RNIPHKN_12_LC_20_16_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_fast_esr_RNIPHKN_12_LC_20_16_1 .LUT_INIT=16'b1101110111101110;
    LogicCell40 \pid_side.error_d_reg_fast_esr_RNIPHKN_12_LC_20_16_1  (
            .in0(N__81865),
            .in1(N__84804),
            .in2(_gnd_net_),
            .in3(N__81901),
            .lcout(\pid_side.error_d_reg_fast_esr_RNIPHKNZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIB8NBA_12_LC_20_16_2 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIB8NBA_12_LC_20_16_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIB8NBA_12_LC_20_16_2 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIB8NBA_12_LC_20_16_2  (
            .in0(N__80057),
            .in1(_gnd_net_),
            .in2(N__80111),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIB8NBAZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI0UI8J_12_LC_20_16_3 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI0UI8J_12_LC_20_16_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI0UI8J_12_LC_20_16_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI0UI8J_12_LC_20_16_3  (
            .in0(N__80015),
            .in1(N__80104),
            .in2(_gnd_net_),
            .in3(N__80056),
            .lcout(\pid_side.error_d_reg_prev_esr_RNI0UI8JZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIGA6A3_13_LC_20_16_4 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIGA6A3_13_LC_20_16_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIGA6A3_13_LC_20_16_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIGA6A3_13_LC_20_16_4  (
            .in0(_gnd_net_),
            .in1(N__83011),
            .in2(_gnd_net_),
            .in3(N__82226),
            .lcout(),
            .ltout(\pid_side.un1_pid_prereg_97_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI45PU7_12_LC_20_16_5 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI45PU7_12_LC_20_16_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI45PU7_12_LC_20_16_5 .LUT_INIT=16'b1110111011101000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI45PU7_12_LC_20_16_5  (
            .in0(N__85443),
            .in1(N__80079),
            .in2(N__80070),
            .in3(N__81798),
            .lcout(\pid_side.error_d_reg_prev_esr_RNI45PU7Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_fast_esr_RNIEIJH2_12_LC_20_16_6 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_fast_esr_RNIEIJH2_12_LC_20_16_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_fast_esr_RNIEIJH2_12_LC_20_16_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \pid_side.error_d_reg_fast_esr_RNIEIJH2_12_LC_20_16_6  (
            .in0(N__82074),
            .in1(N__80043),
            .in2(_gnd_net_),
            .in3(N__80037),
            .lcout(\pid_side.error_d_reg_fast_esr_RNIEIJH2Z0Z_12 ),
            .ltout(\pid_side.error_d_reg_fast_esr_RNIEIJH2Z0Z_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI6P1R3_12_LC_20_16_7 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI6P1R3_12_LC_20_16_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI6P1R3_12_LC_20_16_7 .LUT_INIT=16'b1010010101101001;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI6P1R3_12_LC_20_16_7  (
            .in0(N__83012),
            .in1(N__82271),
            .in2(N__80031),
            .in3(N__82850),
            .lcout(\pid_side.error_d_reg_prev_esr_RNI6P1R3Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIMERG_1_12_LC_20_17_0 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIMERG_1_12_LC_20_17_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIMERG_1_12_LC_20_17_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIMERG_1_12_LC_20_17_0  (
            .in0(_gnd_net_),
            .in1(N__82270),
            .in2(_gnd_net_),
            .in3(N__82851),
            .lcout(),
            .ltout(\pid_side.g1_2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNIDALP2_12_LC_20_17_1 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIDALP2_12_LC_20_17_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIDALP2_12_LC_20_17_1 .LUT_INIT=16'b1100100110010011;
    LogicCell40 \pid_side.error_p_reg_esr_RNIDALP2_12_LC_20_17_1  (
            .in0(N__81684),
            .in1(N__81879),
            .in2(N__80028),
            .in3(N__84800),
            .lcout(),
            .ltout(\pid_side.g1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNILLRS8_12_LC_20_17_2 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNILLRS8_12_LC_20_17_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNILLRS8_12_LC_20_17_2 .LUT_INIT=16'b1000000011101010;
    LogicCell40 \pid_side.error_p_reg_esr_RNILLRS8_12_LC_20_17_2  (
            .in0(N__82023),
            .in1(N__81982),
            .in2(N__80025),
            .in3(N__81087),
            .lcout(\pid_side.error_p_reg_esr_RNILLRS8Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI2OIO_0_13_LC_20_17_3 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI2OIO_0_13_LC_20_17_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI2OIO_0_13_LC_20_17_3 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI2OIO_0_13_LC_20_17_3  (
            .in0(N__85504),
            .in1(N__85548),
            .in2(_gnd_net_),
            .in3(N__85608),
            .lcout(),
            .ltout(\pid_side.N_2405_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI7J5H1_0_14_LC_20_17_4 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI7J5H1_0_14_LC_20_17_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI7J5H1_0_14_LC_20_17_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI7J5H1_0_14_LC_20_17_4  (
            .in0(N__85815),
            .in1(N__84462),
            .in2(N__81093),
            .in3(N__84264),
            .lcout(),
            .ltout(\pid_side.g0_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIQ0PB4_12_LC_20_17_5 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIQ0PB4_12_LC_20_17_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIQ0PB4_12_LC_20_17_5 .LUT_INIT=16'b1101001001001011;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIQ0PB4_12_LC_20_17_5  (
            .in0(N__82284),
            .in1(N__81081),
            .in2(N__81090),
            .in3(N__81783),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIQ0PB4Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI2OIO_3_13_LC_20_17_6 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI2OIO_3_13_LC_20_17_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI2OIO_3_13_LC_20_17_6 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI2OIO_3_13_LC_20_17_6  (
            .in0(N__85609),
            .in1(_gnd_net_),
            .in2(N__85556),
            .in3(N__85505),
            .lcout(\pid_side.N_4_1_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.m12_1_LC_20_18_6 .C_ON=1'b0;
    defparam \pid_side.m12_1_LC_20_18_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.m12_1_LC_20_18_6 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \pid_side.m12_1_LC_20_18_6  (
            .in0(N__81071),
            .in1(N__80857),
            .in2(_gnd_net_),
            .in3(N__80765),
            .lcout(\pid_side.m0_0_03 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_i_reg_esr_RNO_5_12_LC_20_19_7 .C_ON=1'b0;
    defparam \pid_side.error_i_reg_esr_RNO_5_12_LC_20_19_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_i_reg_esr_RNO_5_12_LC_20_19_7 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \pid_side.error_i_reg_esr_RNO_5_12_LC_20_19_7  (
            .in0(N__80608),
            .in1(N__80339),
            .in2(_gnd_net_),
            .in3(N__80201),
            .lcout(\pid_side.m0_2_03 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_4_LC_21_10_0 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_4_LC_21_10_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_4_LC_21_10_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_p_reg_esr_4_LC_21_10_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80178),
            .lcout(\pid_side.error_p_regZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87098),
            .ce(N__85754),
            .sr(N__86023));
    defparam \pid_side.error_p_reg_esr_9_LC_21_10_1 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_9_LC_21_10_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_9_LC_21_10_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_p_reg_esr_9_LC_21_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80169),
            .lcout(\pid_side.error_p_regZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87098),
            .ce(N__85754),
            .sr(N__86023));
    defparam \pid_side.error_p_reg_esr_5_LC_21_10_6 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_5_LC_21_10_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_5_LC_21_10_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_p_reg_esr_5_LC_21_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__80139),
            .lcout(\pid_side.error_p_regZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87098),
            .ce(N__85754),
            .sr(N__86023));
    defparam \pid_side.error_d_reg_esr_5_LC_21_11_1 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_5_LC_21_11_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_5_LC_21_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_esr_5_LC_21_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81396),
            .lcout(\pid_side.error_d_regZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87113),
            .ce(N__85747),
            .sr(N__86020));
    defparam \pid_side.error_p_reg_esr_3_LC_21_11_5 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_3_LC_21_11_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_3_LC_21_11_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_p_reg_esr_3_LC_21_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81345),
            .lcout(\pid_side.error_p_regZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87113),
            .ce(N__85747),
            .sr(N__86020));
    defparam \pid_side.error_d_reg_esr_2_LC_21_11_6 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_2_LC_21_11_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_2_LC_21_11_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_esr_2_LC_21_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81333),
            .lcout(\pid_side.error_d_regZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87113),
            .ce(N__85747),
            .sr(N__86020));
    defparam \pid_side.error_d_reg_esr_10_LC_21_12_0 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_10_LC_21_12_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_10_LC_21_12_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_esr_10_LC_21_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81321),
            .lcout(\pid_side.error_d_regZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87128),
            .ce(N__85710),
            .sr(N__86016));
    defparam \pid_side.error_d_reg_esr_6_LC_21_12_1 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_6_LC_21_12_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_6_LC_21_12_1 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \pid_side.error_d_reg_esr_6_LC_21_12_1  (
            .in0(_gnd_net_),
            .in1(N__81282),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_d_regZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87128),
            .ce(N__85710),
            .sr(N__86016));
    defparam \pid_side.error_d_reg_esr_7_LC_21_12_2 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_7_LC_21_12_2 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_7_LC_21_12_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_esr_7_LC_21_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81246),
            .lcout(\pid_side.error_d_regZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87128),
            .ce(N__85710),
            .sr(N__86016));
    defparam \pid_side.error_d_reg_esr_8_LC_21_12_3 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_8_LC_21_12_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_8_LC_21_12_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_esr_8_LC_21_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81183),
            .lcout(\pid_side.error_d_regZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87128),
            .ce(N__85710),
            .sr(N__86016));
    defparam \pid_side.error_d_reg_esr_9_LC_21_12_4 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_9_LC_21_12_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_9_LC_21_12_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_esr_9_LC_21_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81141),
            .lcout(\pid_side.error_d_regZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87128),
            .ce(N__85710),
            .sr(N__86016));
    defparam \pid_side.error_p_reg_esr_1_LC_21_12_6 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_1_LC_21_12_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_1_LC_21_12_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_p_reg_esr_1_LC_21_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__81105),
            .lcout(\pid_side.error_p_regZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87128),
            .ce(N__85710),
            .sr(N__86016));
    defparam \pid_side.error_p_reg_esr_10_LC_21_12_7 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_10_LC_21_12_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_10_LC_21_12_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_side.error_p_reg_esr_10_LC_21_12_7  (
            .in0(N__81639),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_p_regZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87128),
            .ce(N__85710),
            .sr(N__86016));
    defparam \pid_side.error_d_reg_prev_esr_3_LC_21_13_0 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_3_LC_21_13_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_3_LC_21_13_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_3_LC_21_13_0  (
            .in0(N__82536),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_d_reg_prevZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87143),
            .ce(N__83392),
            .sr(N__83257));
    defparam \pid_side.error_p_reg_esr_RNIFEEQ_3_LC_21_13_1 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIFEEQ_3_LC_21_13_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIFEEQ_3_LC_21_13_1 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_side.error_p_reg_esr_RNIFEEQ_3_LC_21_13_1  (
            .in0(N__81413),
            .in1(N__81422),
            .in2(_gnd_net_),
            .in3(N__82534),
            .lcout(\pid_side.error_p_reg_esr_RNIFEEQZ0Z_3 ),
            .ltout(\pid_side.error_p_reg_esr_RNIFEEQZ0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNIN4BP4_3_LC_21_13_2 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIN4BP4_3_LC_21_13_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIN4BP4_3_LC_21_13_2 .LUT_INIT=16'b1111101010100000;
    LogicCell40 \pid_side.error_p_reg_esr_RNIN4BP4_3_LC_21_13_2  (
            .in0(N__81501),
            .in1(N__81606),
            .in2(N__81588),
            .in3(N__81482),
            .lcout(\pid_side.error_p_reg_esr_RNIN4BP4Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNIIHEQ_0_4_LC_21_13_3 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIIHEQ_0_4_LC_21_13_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIIHEQ_0_4_LC_21_13_3 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_side.error_p_reg_esr_RNIIHEQ_0_4_LC_21_13_3  (
            .in0(N__81567),
            .in1(N__81552),
            .in2(_gnd_net_),
            .in3(N__81520),
            .lcout(\pid_side.error_p_reg_esr_RNIIHEQ_0Z0Z_4 ),
            .ltout(\pid_side.error_p_reg_esr_RNIIHEQ_0Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNI5G8P4_3_LC_21_13_4 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNI5G8P4_3_LC_21_13_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNI5G8P4_3_LC_21_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_p_reg_esr_RNI5G8P4_3_LC_21_13_4  (
            .in0(N__81440),
            .in1(N__81492),
            .in2(N__81486),
            .in3(N__81481),
            .lcout(\pid_side.error_p_reg_esr_RNI5G8P4Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNIUIJC2_2_LC_21_13_5 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIUIJC2_2_LC_21_13_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIUIJC2_2_LC_21_13_5 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_side.error_p_reg_esr_RNIUIJC2_2_LC_21_13_5  (
            .in0(N__82377),
            .in1(N__81402),
            .in2(_gnd_net_),
            .in3(N__81777),
            .lcout(\pid_side.error_p_reg_esr_RNIUIJC2Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNIFEEQ_0_3_LC_21_13_6 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIFEEQ_0_3_LC_21_13_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIFEEQ_0_3_LC_21_13_6 .LUT_INIT=16'b0101101010100101;
    LogicCell40 \pid_side.error_p_reg_esr_RNIFEEQ_0_3_LC_21_13_6  (
            .in0(N__82535),
            .in1(_gnd_net_),
            .in2(N__81426),
            .in3(N__81414),
            .lcout(\pid_side.error_p_reg_esr_RNIFEEQ_0Z0Z_3 ),
            .ltout(\pid_side.error_p_reg_esr_RNIFEEQ_0Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNI7U286_2_LC_21_13_7 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNI7U286_2_LC_21_13_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNI7U286_2_LC_21_13_7 .LUT_INIT=16'b1001011010010110;
    LogicCell40 \pid_side.error_p_reg_esr_RNI7U286_2_LC_21_13_7  (
            .in0(N__82376),
            .in1(N__81776),
            .in2(N__81753),
            .in3(N__82200),
            .lcout(\pid_side.error_p_reg_esr_RNI7U286Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIKAJO_0_19_LC_21_14_0 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIKAJO_0_19_LC_21_14_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIKAJO_0_19_LC_21_14_0 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIKAJO_0_19_LC_21_14_0  (
            .in0(N__84691),
            .in1(N__83597),
            .in2(_gnd_net_),
            .in3(N__81710),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIKAJO_0Z0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_19_LC_21_14_1 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_19_LC_21_14_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_19_LC_21_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_19_LC_21_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84693),
            .lcout(\pid_side.error_d_reg_prevZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87161),
            .ce(N__83405),
            .sr(N__83256));
    defparam \pid_side.error_d_reg_prev_esr_RNIKAJO_19_LC_21_14_2 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIKAJO_19_LC_21_14_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIKAJO_19_LC_21_14_2 .LUT_INIT=16'b1000100011101110;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIKAJO_19_LC_21_14_2  (
            .in0(N__84692),
            .in1(N__83598),
            .in2(_gnd_net_),
            .in3(N__81711),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIKAJOZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNISHIO_11_LC_21_14_3 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNISHIO_11_LC_21_14_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNISHIO_11_LC_21_14_3 .LUT_INIT=16'b1111010101010000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNISHIO_11_LC_21_14_3  (
            .in0(N__81831),
            .in1(_gnd_net_),
            .in2(N__82341),
            .in3(N__82893),
            .lcout(\pid_side.g0_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNISHIO_2_11_LC_21_14_4 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNISHIO_2_11_LC_21_14_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNISHIO_2_11_LC_21_14_4 .LUT_INIT=16'b0100010011011101;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNISHIO_2_11_LC_21_14_4  (
            .in0(N__82891),
            .in1(N__81829),
            .in2(_gnd_net_),
            .in3(N__82332),
            .lcout(\pid_side.g0_19_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNISHIO_1_11_LC_21_14_5 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNISHIO_1_11_LC_21_14_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNISHIO_1_11_LC_21_14_5 .LUT_INIT=16'b0101101010100101;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNISHIO_1_11_LC_21_14_5  (
            .in0(N__81830),
            .in1(_gnd_net_),
            .in2(N__82340),
            .in3(N__82892),
            .lcout(\pid_side.error_d_reg_prev_esr_RNISHIO_1Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNISKLO_0_20_LC_21_14_6 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNISKLO_0_20_LC_21_14_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNISKLO_0_20_LC_21_14_6 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNISKLO_0_20_LC_21_14_6  (
            .in0(N__84536),
            .in1(N__84284),
            .in2(_gnd_net_),
            .in3(N__82976),
            .lcout(\pid_side.error_d_reg_prev_esr_RNISKLO_0Z0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_20_LC_21_14_7 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_20_LC_21_14_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_20_LC_21_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_20_LC_21_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84537),
            .lcout(\pid_side.error_d_reg_prevZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87161),
            .ce(N__83405),
            .sr(N__83256));
    defparam \pid_side.error_d_reg_prev_esr_RNISHIO_0_11_LC_21_15_0 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNISHIO_0_11_LC_21_15_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNISHIO_0_11_LC_21_15_0 .LUT_INIT=16'b1111010100000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNISHIO_0_11_LC_21_15_0  (
            .in0(N__81828),
            .in1(_gnd_net_),
            .in2(N__82339),
            .in3(N__82889),
            .lcout(\pid_side.un1_pid_prereg_135_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_11_LC_21_15_1 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_11_LC_21_15_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_11_LC_21_15_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_11_LC_21_15_1  (
            .in0(N__82890),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_d_reg_prevZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87174),
            .ce(N__83403),
            .sr(N__83240));
    defparam \pid_side.error_d_reg_fast_esr_RNIGBTF_0_12_LC_21_15_2 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_fast_esr_RNIGBTF_0_12_LC_21_15_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_fast_esr_RNIGBTF_0_12_LC_21_15_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \pid_side.error_d_reg_fast_esr_RNIGBTF_0_12_LC_21_15_2  (
            .in0(_gnd_net_),
            .in1(N__81902),
            .in2(_gnd_net_),
            .in3(N__81870),
            .lcout(\pid_side.N_2398_i ),
            .ltout(\pid_side.N_2398_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNIL0VP1_12_LC_21_15_3 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIL0VP1_12_LC_21_15_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIL0VP1_12_LC_21_15_3 .LUT_INIT=16'b0011110001101001;
    LogicCell40 \pid_side.error_p_reg_esr_RNIL0VP1_12_LC_21_15_3  (
            .in0(N__82076),
            .in1(N__84799),
            .in2(N__81846),
            .in3(N__82052),
            .lcout(\pid_side.error_p_reg_esr_RNIL0VP1Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_fast_esr_12_LC_21_15_4 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_fast_esr_12_LC_21_15_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_fast_esr_12_LC_21_15_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_side.error_d_reg_prev_fast_esr_12_LC_21_15_4  (
            .in0(N__82834),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_d_reg_prev_fastZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87174),
            .ce(N__83403),
            .sr(N__83240));
    defparam \pid_side.error_d_reg_prev_esr_RNI0TN9_11_LC_21_15_5 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI0TN9_11_LC_21_15_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI0TN9_11_LC_21_15_5 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI0TN9_11_LC_21_15_5  (
            .in0(_gnd_net_),
            .in1(N__82328),
            .in2(_gnd_net_),
            .in3(N__81827),
            .lcout(\pid_side.un1_pid_prereg_79 ),
            .ltout(\pid_side.un1_pid_prereg_79_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNIL0VP1_0_12_LC_21_15_6 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIL0VP1_0_12_LC_21_15_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIL0VP1_0_12_LC_21_15_6 .LUT_INIT=16'b0100010001001101;
    LogicCell40 \pid_side.error_p_reg_esr_RNIL0VP1_0_12_LC_21_15_6  (
            .in0(N__84798),
            .in1(N__81810),
            .in2(N__81804),
            .in3(N__82075),
            .lcout(),
            .ltout(\pid_side.un1_pid_prereg_167_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNID7D33_12_LC_21_15_7 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNID7D33_12_LC_21_15_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNID7D33_12_LC_21_15_7 .LUT_INIT=16'b1100111101000101;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNID7D33_12_LC_21_15_7  (
            .in0(N__82277),
            .in1(N__83002),
            .in2(N__81801),
            .in3(N__82833),
            .lcout(\pid_side.un1_pid_prereg_167_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_12_LC_21_16_0 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_12_LC_21_16_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_12_LC_21_16_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_12_LC_21_16_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82832),
            .lcout(\pid_side.error_d_reg_prevZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87188),
            .ce(N__83401),
            .sr(N__83244));
    defparam \pid_side.error_p_reg_esr_RNIR65H1_12_LC_21_16_1 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIR65H1_12_LC_21_16_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIR65H1_12_LC_21_16_1 .LUT_INIT=16'b1101010001001101;
    LogicCell40 \pid_side.error_p_reg_esr_RNIR65H1_12_LC_21_16_1  (
            .in0(N__84806),
            .in1(N__81792),
            .in2(N__82843),
            .in3(N__82269),
            .lcout(\pid_side.g0_19_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIMERG_12_LC_21_16_3 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIMERG_12_LC_21_16_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIMERG_12_LC_21_16_3 .LUT_INIT=16'b1010111110101111;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIMERG_12_LC_21_16_3  (
            .in0(N__82827),
            .in1(_gnd_net_),
            .in2(N__82272),
            .in3(_gnd_net_),
            .lcout(\pid_side.N_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIMERG_2_12_LC_21_16_4 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIMERG_2_12_LC_21_16_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIMERG_2_12_LC_21_16_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIMERG_2_12_LC_21_16_4  (
            .in0(_gnd_net_),
            .in1(N__82257),
            .in2(_gnd_net_),
            .in3(N__82831),
            .lcout(),
            .ltout(\pid_side.N_3_i_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNIR3TQ1_12_LC_21_16_5 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIR3TQ1_12_LC_21_16_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIR3TQ1_12_LC_21_16_5 .LUT_INIT=16'b0000010100010111;
    LogicCell40 \pid_side.error_p_reg_esr_RNIR3TQ1_12_LC_21_16_5  (
            .in0(N__84805),
            .in1(N__82077),
            .in2(N__82056),
            .in3(N__82053),
            .lcout(),
            .ltout(\pid_side.N_3_i_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIQTGL4_12_LC_21_16_6 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIQTGL4_12_LC_21_16_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIQTGL4_12_LC_21_16_6 .LUT_INIT=16'b0010101111010100;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIQTGL4_12_LC_21_16_6  (
            .in0(N__82035),
            .in1(N__85620),
            .in2(N__82026),
            .in3(N__84231),
            .lcout(),
            .ltout(\pid_side.error_d_reg_prev_esr_RNIQTGL4Z0Z_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIE108A_12_LC_21_16_7 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIE108A_12_LC_21_16_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIE108A_12_LC_21_16_7 .LUT_INIT=16'b1001011001011010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIE108A_12_LC_21_16_7  (
            .in0(N__82022),
            .in1(N__81984),
            .in2(N__81939),
            .in3(N__81936),
            .lcout(\pid_side.un1_pid_prereg_0_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_fast_esr_RNIGBTF_12_LC_21_17_2 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_fast_esr_RNIGBTF_12_LC_21_17_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_fast_esr_RNIGBTF_12_LC_21_17_2 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \pid_side.error_d_reg_fast_esr_RNIGBTF_12_LC_21_17_2  (
            .in0(_gnd_net_),
            .in1(N__81906),
            .in2(_gnd_net_),
            .in3(N__81869),
            .lcout(),
            .ltout(\pid_side.g1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNII3G81_13_LC_21_17_3 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNII3G81_13_LC_21_17_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNII3G81_13_LC_21_17_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNII3G81_13_LC_21_17_3  (
            .in0(N__85506),
            .in1(N__85610),
            .in2(N__81882),
            .in3(N__85537),
            .lcout(\pid_side.g0_3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_fast_esr_12_LC_21_17_4 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_fast_esr_12_LC_21_17_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_fast_esr_12_LC_21_17_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_fast_esr_12_LC_21_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82872),
            .lcout(\pid_side.error_d_reg_fastZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87205),
            .ce(N__85753),
            .sr(N__86010));
    defparam \pid_side.error_d_reg_prev_esr_RNIMERG_0_12_LC_21_17_6 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIMERG_0_12_LC_21_17_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIMERG_0_12_LC_21_17_6 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIMERG_0_12_LC_21_17_6  (
            .in0(_gnd_net_),
            .in1(N__82273),
            .in2(_gnd_net_),
            .in3(N__82841),
            .lcout(\pid_side.N_5_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI41F23_12_LC_21_17_7 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI41F23_12_LC_21_17_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI41F23_12_LC_21_17_7 .LUT_INIT=16'b0101000010101111;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI41F23_12_LC_21_17_7  (
            .in0(N__82842),
            .in1(_gnd_net_),
            .in2(N__82278),
            .in3(N__82227),
            .lcout(\pid_side.error_d_reg_prev_esr_RNI41F23Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI9BFR3_1_LC_22_11_0 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI9BFR3_1_LC_22_11_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI9BFR3_1_LC_22_11_0 .LUT_INIT=16'b1110111110001100;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI9BFR3_1_LC_22_11_0  (
            .in0(N__83045),
            .in1(N__82608),
            .in2(N__82511),
            .in3(N__82176),
            .lcout(\pid_side.error_d_reg_prev_esr_RNI9BFR3Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNIIQL11_0_1_LC_22_11_1 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIIQL11_0_1_LC_22_11_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIIQL11_0_1_LC_22_11_1 .LUT_INIT=16'b1000110011101111;
    LogicCell40 \pid_side.error_p_reg_esr_RNIIQL11_0_1_LC_22_11_1  (
            .in0(N__82564),
            .in1(N__82480),
            .in2(N__82102),
            .in3(N__83043),
            .lcout(),
            .ltout(\pid_side.error_p_reg_esr_RNIIQL11_0Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIBGIE2_1_LC_22_11_2 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIBGIE2_1_LC_22_11_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIBGIE2_1_LC_22_11_2 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIBGIE2_1_LC_22_11_2  (
            .in0(N__82504),
            .in1(_gnd_net_),
            .in2(N__82179),
            .in3(N__82122),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIBGIE2Z0Z_1 ),
            .ltout(\pid_side.error_d_reg_prev_esr_RNIBGIE2Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI905J4_1_LC_22_11_3 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI905J4_1_LC_22_11_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI905J4_1_LC_22_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI905J4_1_LC_22_11_3  (
            .in0(N__82170),
            .in1(N__82607),
            .in2(N__82134),
            .in3(N__82116),
            .lcout(\pid_side.error_d_reg_prev_esr_RNI905J4Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNIIQL11_1_LC_22_11_4 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNIIQL11_1_LC_22_11_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNIIQL11_1_LC_22_11_4 .LUT_INIT=16'b1110100011111010;
    LogicCell40 \pid_side.error_p_reg_esr_RNIIQL11_1_LC_22_11_4  (
            .in0(N__83042),
            .in1(N__82563),
            .in2(N__82482),
            .in3(N__82092),
            .lcout(\pid_side.error_p_reg_esr_RNIIQL11Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIIFEI_1_LC_22_11_5 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIIFEI_1_LC_22_11_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIIFEI_1_LC_22_11_5 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIIFEI_1_LC_22_11_5  (
            .in0(_gnd_net_),
            .in1(N__82503),
            .in2(_gnd_net_),
            .in3(N__83044),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIIFEIZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_0_LC_22_11_6 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_0_LC_22_11_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_0_LC_22_11_6 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \pid_side.error_d_reg_prev_esr_0_LC_22_11_6  (
            .in0(_gnd_net_),
            .in1(N__82565),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_d_reg_prevZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87129),
            .ce(N__83398),
            .sr(N__83262));
    defparam \pid_side.error_p_reg_esr_RNICBEQ_0_2_LC_22_11_7 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNICBEQ_0_2_LC_22_11_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNICBEQ_0_2_LC_22_11_7 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_side.error_p_reg_esr_RNICBEQ_0_2_LC_22_11_7  (
            .in0(N__82421),
            .in1(N__82406),
            .in2(_gnd_net_),
            .in3(N__82438),
            .lcout(\pid_side.error_p_reg_esr_RNICBEQ_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_esr_0_LC_22_12_1 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_0_LC_22_12_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_0_LC_22_12_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_esr_0_LC_22_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82596),
            .lcout(\pid_side.error_d_regZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87144),
            .ce(N__85708),
            .sr(N__86021));
    defparam \pid_side.error_d_reg_esr_3_LC_22_12_2 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_3_LC_22_12_2 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_3_LC_22_12_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_esr_3_LC_22_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82548),
            .lcout(\pid_side.error_d_regZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87144),
            .ce(N__85708),
            .sr(N__86021));
    defparam \pid_side.error_p_reg_esr_2_LC_22_12_3 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_2_LC_22_12_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_2_LC_22_12_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_p_reg_esr_2_LC_22_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82524),
            .lcout(\pid_side.error_p_regZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87144),
            .ce(N__85708),
            .sr(N__86021));
    defparam \pid_side.error_p_reg_esr_RNI98EQ_1_LC_22_13_1 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNI98EQ_1_LC_22_13_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNI98EQ_1_LC_22_13_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_side.error_p_reg_esr_RNI98EQ_1_LC_22_13_1  (
            .in0(N__82512),
            .in1(N__82481),
            .in2(_gnd_net_),
            .in3(N__83041),
            .lcout(\pid_side.un1_pid_prereg_9_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_RNICBEQ_2_LC_22_13_2 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_RNICBEQ_2_LC_22_13_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_p_reg_esr_RNICBEQ_2_LC_22_13_2 .LUT_INIT=16'b1000100011101110;
    LogicCell40 \pid_side.error_p_reg_esr_RNICBEQ_2_LC_22_13_2  (
            .in0(N__82445),
            .in1(N__82422),
            .in2(_gnd_net_),
            .in3(N__82410),
            .lcout(\pid_side.error_p_reg_esr_RNICBEQZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.state_RNIK1B71_0_LC_22_13_7 .C_ON=1'b0;
    defparam \pid_side.state_RNIK1B71_0_LC_22_13_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.state_RNIK1B71_0_LC_22_13_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \pid_side.state_RNIK1B71_0_LC_22_13_7  (
            .in0(_gnd_net_),
            .in1(N__82368),
            .in2(_gnd_net_),
            .in3(N__86152),
            .lcout(\pid_side.N_873_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_esr_11_LC_22_14_0 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_11_LC_22_14_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_11_LC_22_14_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_p_reg_esr_11_LC_22_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82353),
            .lcout(\pid_side.error_p_regZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87175),
            .ce(N__85709),
            .sr(N__86015));
    defparam \pid_side.error_d_reg_esr_15_LC_22_15_0 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_15_LC_22_15_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_15_LC_22_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_esr_15_LC_22_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82311),
            .lcout(\pid_side.error_d_regZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87189),
            .ce(N__85724),
            .sr(N__86013));
    defparam \pid_side.error_d_reg_esr_11_LC_22_15_2 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_11_LC_22_15_2 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_11_LC_22_15_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_esr_11_LC_22_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82905),
            .lcout(\pid_side.error_d_regZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87189),
            .ce(N__85724),
            .sr(N__86013));
    defparam \pid_side.error_d_reg_esr_12_LC_22_15_7 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_12_LC_22_15_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_12_LC_22_15_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_esr_12_LC_22_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82868),
            .lcout(\pid_side.error_d_regZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87189),
            .ce(N__85724),
            .sr(N__86013));
    defparam \pid_side.error_d_reg_prev_esr_13_LC_22_16_4 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_13_LC_22_16_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_13_LC_22_16_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_13_LC_22_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85611),
            .lcout(\pid_side.error_d_reg_prevZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87206),
            .ce(N__83404),
            .sr(N__83236));
    defparam \pid_front.error_d_reg_esr_14_LC_22_23_3 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_14_LC_22_23_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_14_LC_22_23_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_esr_14_LC_22_23_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__82788),
            .lcout(\pid_front.error_d_regZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87267),
            .ce(N__86339),
            .sr(N__86003));
    defparam \Commands_frame_decoder.source_xy_kp_e_0_1_LC_23_11_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_kp_e_0_1_LC_23_11_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_kp_e_0_1_LC_23_11_7 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_xy_kp_e_0_1_LC_23_11_7  (
            .in0(_gnd_net_),
            .in1(N__84204),
            .in2(_gnd_net_),
            .in3(N__86165),
            .lcout(xy_kp_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87145),
            .ce(N__82692),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIB1JO_16_LC_23_13_0 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIB1JO_16_LC_23_13_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIB1JO_16_LC_23_13_0 .LUT_INIT=16'b1000100011101110;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIB1JO_16_LC_23_13_0  (
            .in0(N__85772),
            .in1(N__84309),
            .in2(_gnd_net_),
            .in3(N__82937),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIB1JOZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_16_LC_23_13_1 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_16_LC_23_13_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_16_LC_23_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_prev_esr_16_LC_23_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85773),
            .lcout(\pid_side.error_d_reg_prevZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87176),
            .ce(N__83406),
            .sr(N__83255));
    defparam \pid_side.error_d_reg_prev_esr_RNIE4JO_0_17_LC_23_13_2 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIE4JO_0_17_LC_23_13_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIE4JO_0_17_LC_23_13_2 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIE4JO_0_17_LC_23_13_2  (
            .in0(N__84350),
            .in1(N__83450),
            .in2(_gnd_net_),
            .in3(N__84736),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIE4JO_0Z0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_17_LC_23_13_3 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_17_LC_23_13_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_17_LC_23_13_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_17_LC_23_13_3  (
            .in0(N__84738),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_d_reg_prevZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87176),
            .ce(N__83406),
            .sr(N__83255));
    defparam \pid_side.error_d_reg_prev_esr_RNIE4JO_17_LC_23_13_4 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIE4JO_17_LC_23_13_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIE4JO_17_LC_23_13_4 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIE4JO_17_LC_23_13_4  (
            .in0(N__84351),
            .in1(N__83451),
            .in2(_gnd_net_),
            .in3(N__84737),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIE4JOZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIH7JO_0_18_LC_23_13_5 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIH7JO_0_18_LC_23_13_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIH7JO_0_18_LC_23_13_5 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIH7JO_0_18_LC_23_13_5  (
            .in0(N__83465),
            .in1(N__83102),
            .in2(_gnd_net_),
            .in3(N__84715),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIH7JO_0Z0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_18_LC_23_13_6 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_18_LC_23_13_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_prev_esr_18_LC_23_13_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_18_LC_23_13_6  (
            .in0(N__84717),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_d_reg_prevZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87176),
            .ce(N__83406),
            .sr(N__83255));
    defparam \pid_side.error_d_reg_prev_esr_RNIH7JO_18_LC_23_13_7 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIH7JO_18_LC_23_13_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIH7JO_18_LC_23_13_7 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIH7JO_18_LC_23_13_7  (
            .in0(N__83466),
            .in1(N__83103),
            .in2(_gnd_net_),
            .in3(N__84716),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIH7JOZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_esr_1_LC_23_14_4 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_1_LC_23_14_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_1_LC_23_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_esr_1_LC_23_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__83064),
            .lcout(\pid_side.error_d_regZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87190),
            .ce(N__85728),
            .sr(N__86017));
    defparam \pid_side.error_d_reg_prev_esr_RNI2OIO_4_13_LC_23_15_2 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI2OIO_4_13_LC_23_15_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI2OIO_4_13_LC_23_15_2 .LUT_INIT=16'b0101101010100101;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI2OIO_4_13_LC_23_15_2  (
            .in0(N__85530),
            .in1(_gnd_net_),
            .in2(N__85503),
            .in3(N__85586),
            .lcout(\pid_side.error_d_reg_prev_esr_RNI2OIO_4Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNISKLO_20_LC_23_15_5 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNISKLO_20_LC_23_15_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNISKLO_20_LC_23_15_5 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNISKLO_20_LC_23_15_5  (
            .in0(N__84285),
            .in1(N__82983),
            .in2(_gnd_net_),
            .in3(N__84535),
            .lcout(\pid_side.error_d_reg_prev_esr_RNISKLOZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNIB1JO_0_16_LC_23_15_7 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNIB1JO_0_16_LC_23_15_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNIB1JO_0_16_LC_23_15_7 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNIB1JO_0_16_LC_23_15_7  (
            .in0(N__84308),
            .in1(N__82938),
            .in2(_gnd_net_),
            .in3(N__85766),
            .lcout(\pid_side.error_d_reg_prev_esr_RNIB1JO_0Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI2OIO_13_LC_23_16_2 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI2OIO_13_LC_23_16_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI2OIO_13_LC_23_16_2 .LUT_INIT=16'b1101110101000100;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI2OIO_13_LC_23_16_2  (
            .in0(N__85529),
            .in1(N__85489),
            .in2(_gnd_net_),
            .in3(N__85585),
            .lcout(),
            .ltout(\pid_side.N_2405_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI7J5H1_14_LC_23_16_3 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI7J5H1_14_LC_23_16_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI7J5H1_14_LC_23_16_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI7J5H1_14_LC_23_16_3  (
            .in0(N__84458),
            .in1(N__84260),
            .in2(N__84234),
            .in3(N__85798),
            .lcout(\pid_side.g0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_xy_kd_1_LC_23_17_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_kd_1_LC_23_17_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_kd_1_LC_23_17_7 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_xy_kd_1_LC_23_17_7  (
            .in0(_gnd_net_),
            .in1(N__84215),
            .in2(_gnd_net_),
            .in3(N__86157),
            .lcout(xy_kd_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87237),
            .ce(N__84866),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_xy_kd_3_LC_23_19_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_kd_3_LC_23_19_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_kd_3_LC_23_19_5 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_xy_kd_3_LC_23_19_5  (
            .in0(_gnd_net_),
            .in1(N__84028),
            .in2(_gnd_net_),
            .in3(N__86154),
            .lcout(xy_kd_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87253),
            .ce(N__84867),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_xy_kd_0_LC_23_21_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_kd_0_LC_23_21_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_kd_0_LC_23_21_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_xy_kd_0_LC_23_21_1  (
            .in0(_gnd_net_),
            .in1(N__83836),
            .in2(_gnd_net_),
            .in3(N__86153),
            .lcout(xy_kd_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87263),
            .ce(N__84873),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_esr_20_LC_23_23_1 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_20_LC_23_23_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_20_LC_23_23_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_esr_20_LC_23_23_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__83655),
            .lcout(\pid_front.error_d_regZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87271),
            .ce(N__86340),
            .sr(N__86004));
    defparam \pid_side.error_p_reg_esr_19_LC_24_10_0 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_19_LC_24_10_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_19_LC_24_10_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_side.error_p_reg_esr_19_LC_24_10_0  (
            .in0(N__83607),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_p_regZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87146),
            .ce(N__85745),
            .sr(N__86028));
    defparam \pid_side.error_p_reg_esr_21_LC_24_10_2 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_21_LC_24_10_2 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_21_LC_24_10_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_p_reg_esr_21_LC_24_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__83583),
            .lcout(\pid_side.error_p_regZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87146),
            .ce(N__85745),
            .sr(N__86028));
    defparam \pid_side.error_p_reg_esr_18_LC_24_10_4 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_18_LC_24_10_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_18_LC_24_10_4 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \pid_side.error_p_reg_esr_18_LC_24_10_4  (
            .in0(_gnd_net_),
            .in1(N__83475),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_p_regZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87146),
            .ce(N__85745),
            .sr(N__86028));
    defparam \pid_side.error_p_reg_esr_14_LC_24_10_5 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_14_LC_24_10_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_14_LC_24_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_p_reg_esr_14_LC_24_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84471),
            .lcout(\pid_side.error_p_regZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87146),
            .ce(N__85745),
            .sr(N__86028));
    defparam \pid_side.error_p_reg_esr_7_LC_24_10_7 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_7_LC_24_10_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_7_LC_24_10_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_p_reg_esr_7_LC_24_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84423),
            .lcout(\pid_side.error_p_regZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87146),
            .ce(N__85745),
            .sr(N__86028));
    defparam \pid_side.error_p_reg_esr_8_LC_24_11_0 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_8_LC_24_11_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_8_LC_24_11_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_p_reg_esr_8_LC_24_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84390),
            .lcout(\pid_side.error_p_regZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87162),
            .ce(N__85751),
            .sr(N__86025));
    defparam \pid_side.error_p_reg_esr_13_LC_24_11_2 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_13_LC_24_11_2 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_13_LC_24_11_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_p_reg_esr_13_LC_24_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84363),
            .lcout(\pid_side.error_p_regZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87162),
            .ce(N__85751),
            .sr(N__86025));
    defparam \pid_side.error_p_reg_esr_17_LC_24_11_3 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_17_LC_24_11_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_17_LC_24_11_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_p_reg_esr_17_LC_24_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84357),
            .lcout(\pid_side.error_p_regZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87162),
            .ce(N__85751),
            .sr(N__86025));
    defparam \pid_side.error_p_reg_esr_15_LC_24_11_4 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_15_LC_24_11_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_15_LC_24_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_p_reg_esr_15_LC_24_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84336),
            .lcout(\pid_side.error_p_regZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87162),
            .ce(N__85751),
            .sr(N__86025));
    defparam \pid_side.error_p_reg_esr_16_LC_24_11_5 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_16_LC_24_11_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_16_LC_24_11_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_p_reg_esr_16_LC_24_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84315),
            .lcout(\pid_side.error_p_regZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87162),
            .ce(N__85751),
            .sr(N__86025));
    defparam \pid_side.error_p_reg_esr_20_LC_24_11_6 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_20_LC_24_11_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_20_LC_24_11_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_p_reg_esr_20_LC_24_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84291),
            .lcout(\pid_side.error_p_regZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87162),
            .ce(N__85751),
            .sr(N__86025));
    defparam \pid_side.error_p_reg_esr_12_LC_24_12_0 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_12_LC_24_12_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_12_LC_24_12_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_p_reg_esr_12_LC_24_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84813),
            .lcout(\pid_side.error_p_regZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87177),
            .ce(N__85755),
            .sr(N__86024));
    defparam \pid_side.error_d_reg_esr_17_LC_24_14_0 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_17_LC_24_14_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_17_LC_24_14_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_esr_17_LC_24_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84750),
            .lcout(\pid_side.error_d_regZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87207),
            .ce(N__85741),
            .sr(N__86022));
    defparam \pid_side.error_d_reg_esr_18_LC_24_14_1 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_18_LC_24_14_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_18_LC_24_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_esr_18_LC_24_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84726),
            .lcout(\pid_side.error_d_regZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87207),
            .ce(N__85741),
            .sr(N__86022));
    defparam \pid_side.error_d_reg_esr_19_LC_24_14_2 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_19_LC_24_14_2 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_19_LC_24_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_esr_19_LC_24_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84705),
            .lcout(\pid_side.error_d_regZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87207),
            .ce(N__85741),
            .sr(N__86022));
    defparam \pid_side.error_d_reg_esr_21_LC_24_14_4 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_21_LC_24_14_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_21_LC_24_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_esr_21_LC_24_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84678),
            .lcout(\pid_side.error_d_regZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87207),
            .ce(N__85741),
            .sr(N__86022));
    defparam \pid_side.error_d_reg_esr_22_LC_24_14_5 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_22_LC_24_14_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_22_LC_24_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_esr_22_LC_24_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84645),
            .lcout(\pid_side.error_d_regZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87207),
            .ce(N__85741),
            .sr(N__86022));
    defparam \pid_side.error_d_reg_esr_20_LC_24_15_1 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_20_LC_24_15_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_20_LC_24_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_esr_20_LC_24_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84546),
            .lcout(\pid_side.error_d_regZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87222),
            .ce(N__85752),
            .sr(N__86018));
    defparam \pid_side.error_p_reg_esr_0_LC_24_15_2 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_esr_0_LC_24_15_2 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_esr_0_LC_24_15_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_p_reg_esr_0_LC_24_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84516),
            .lcout(\pid_side.error_p_regZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87222),
            .ce(N__85752),
            .sr(N__86018));
    defparam \pid_side.error_d_reg_esr_13_LC_24_15_4 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_13_LC_24_15_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_13_LC_24_15_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_esr_13_LC_24_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__84477),
            .lcout(\pid_side.error_d_regZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87222),
            .ce(N__85752),
            .sr(N__86018));
    defparam \pid_side.error_d_reg_esr_14_LC_24_15_5 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_14_LC_24_15_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_14_LC_24_15_5 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \pid_side.error_d_reg_esr_14_LC_24_15_5  (
            .in0(_gnd_net_),
            .in1(N__85824),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_d_regZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87222),
            .ce(N__85752),
            .sr(N__86018));
    defparam \pid_side.error_d_reg_esr_16_LC_24_15_7 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_esr_16_LC_24_15_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_d_reg_esr_16_LC_24_15_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.error_d_reg_esr_16_LC_24_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85782),
            .lcout(\pid_side.error_d_regZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87222),
            .ce(N__85752),
            .sr(N__86018));
    defparam \pid_side.error_d_reg_prev_esr_RNI2OIO_2_13_LC_24_16_3 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI2OIO_2_13_LC_24_16_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI2OIO_2_13_LC_24_16_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI2OIO_2_13_LC_24_16_3  (
            .in0(N__85490),
            .in1(N__85552),
            .in2(_gnd_net_),
            .in3(N__85592),
            .lcout(\pid_side.N_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_d_reg_prev_esr_RNI2OIO_1_13_LC_24_16_6 .C_ON=1'b0;
    defparam \pid_side.error_d_reg_prev_esr_RNI2OIO_1_13_LC_24_16_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_d_reg_prev_esr_RNI2OIO_1_13_LC_24_16_6 .LUT_INIT=16'b1010111100001010;
    LogicCell40 \pid_side.error_d_reg_prev_esr_RNI2OIO_1_13_LC_24_16_6  (
            .in0(N__85593),
            .in1(_gnd_net_),
            .in2(N__85557),
            .in3(N__85491),
            .lcout(\pid_side.error_d_reg_prev_esr_RNI2OIO_1Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_esr_2_LC_24_17_1 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_2_LC_24_17_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_2_LC_24_17_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_esr_2_LC_24_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85434),
            .lcout(\pid_front.error_d_regZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87248),
            .ce(N__86319),
            .sr(N__86014));
    defparam \Commands_frame_decoder.source_xy_kd_7_LC_24_18_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_kd_7_LC_24_18_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_kd_7_LC_24_18_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_xy_kd_7_LC_24_18_2  (
            .in0(_gnd_net_),
            .in1(N__85404),
            .in2(_gnd_net_),
            .in3(N__86160),
            .lcout(xy_kd_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87254),
            .ce(N__84869),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_xy_kd_5_LC_24_19_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_kd_5_LC_24_19_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_kd_5_LC_24_19_2 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Commands_frame_decoder.source_xy_kd_5_LC_24_19_2  (
            .in0(N__86156),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__85215),
            .lcout(xy_kd_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87259),
            .ce(N__84868),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_xy_kd_4_LC_24_19_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_kd_4_LC_24_19_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_kd_4_LC_24_19_7 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_xy_kd_4_LC_24_19_7  (
            .in0(_gnd_net_),
            .in1(N__85040),
            .in2(_gnd_net_),
            .in3(N__86155),
            .lcout(xy_kd_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87259),
            .ce(N__84868),
            .sr(_gnd_net_));
    defparam \pid_front.error_d_reg_esr_17_LC_24_22_0 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_17_LC_24_22_0 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_17_LC_24_22_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_front.error_d_reg_esr_17_LC_24_22_0  (
            .in0(N__87588),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_d_regZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87272),
            .ce(N__86336),
            .sr(N__86008));
    defparam \pid_front.error_d_reg_esr_18_LC_24_22_1 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_18_LC_24_22_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_18_LC_24_22_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_esr_18_LC_24_22_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__87555),
            .lcout(\pid_front.error_d_regZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87272),
            .ce(N__86336),
            .sr(N__86008));
    defparam \pid_front.error_d_reg_esr_19_LC_24_22_2 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_19_LC_24_22_2 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_19_LC_24_22_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_front.error_d_reg_esr_19_LC_24_22_2  (
            .in0(N__87516),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_d_regZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87272),
            .ce(N__86336),
            .sr(N__86008));
    defparam \pid_front.error_d_reg_esr_21_LC_24_22_5 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_21_LC_24_22_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_21_LC_24_22_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_esr_21_LC_24_22_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__87477),
            .lcout(\pid_front.error_d_regZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87272),
            .ce(N__86336),
            .sr(N__86008));
    defparam \pid_front.error_d_reg_esr_22_LC_24_22_6 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_22_LC_24_22_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_22_LC_24_22_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_esr_22_LC_24_22_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__87441),
            .lcout(\pid_front.error_d_regZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87272),
            .ce(N__86336),
            .sr(N__86008));
    defparam \pid_front.error_d_reg_esr_15_LC_24_23_1 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_15_LC_24_23_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_15_LC_24_23_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_front.error_d_reg_esr_15_LC_24_23_1  (
            .in0(N__87333),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_d_regZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87276),
            .ce(N__86338),
            .sr(N__86006));
    defparam \pid_front.error_d_reg_esr_16_LC_24_24_5 .C_ON=1'b0;
    defparam \pid_front.error_d_reg_esr_16_LC_24_24_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_d_reg_esr_16_LC_24_24_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.error_d_reg_esr_16_LC_24_24_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__87303),
            .lcout(\pid_front.error_d_regZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__87279),
            .ce(N__86337),
            .sr(N__86005));
endmodule // Pc2drone
