-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 11 2017 17:29:57

-- File Generated:     May 16 2019 21:18:00

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "Pc2Drone" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of Pc2Drone
entity Pc2Drone is
port (
    ppm_output : out std_logic;
    uart_input_debug : out std_logic;
    uart_input : in std_logic;
    frame_decoder_dv : out std_logic;
    clk_system : in std_logic);
end Pc2Drone;

-- Architecture of Pc2Drone
-- View name is \INTERFACE\
architecture \INTERFACE\ of Pc2Drone is

signal \N__24858\ : std_logic;
signal \N__24857\ : std_logic;
signal \N__24856\ : std_logic;
signal \N__24847\ : std_logic;
signal \N__24846\ : std_logic;
signal \N__24845\ : std_logic;
signal \N__24838\ : std_logic;
signal \N__24837\ : std_logic;
signal \N__24836\ : std_logic;
signal \N__24829\ : std_logic;
signal \N__24828\ : std_logic;
signal \N__24827\ : std_logic;
signal \N__24820\ : std_logic;
signal \N__24819\ : std_logic;
signal \N__24818\ : std_logic;
signal \N__24801\ : std_logic;
signal \N__24798\ : std_logic;
signal \N__24795\ : std_logic;
signal \N__24792\ : std_logic;
signal \N__24789\ : std_logic;
signal \N__24786\ : std_logic;
signal \N__24783\ : std_logic;
signal \N__24780\ : std_logic;
signal \N__24777\ : std_logic;
signal \N__24774\ : std_logic;
signal \N__24771\ : std_logic;
signal \N__24770\ : std_logic;
signal \N__24769\ : std_logic;
signal \N__24768\ : std_logic;
signal \N__24767\ : std_logic;
signal \N__24764\ : std_logic;
signal \N__24761\ : std_logic;
signal \N__24758\ : std_logic;
signal \N__24757\ : std_logic;
signal \N__24754\ : std_logic;
signal \N__24751\ : std_logic;
signal \N__24750\ : std_logic;
signal \N__24749\ : std_logic;
signal \N__24748\ : std_logic;
signal \N__24747\ : std_logic;
signal \N__24746\ : std_logic;
signal \N__24745\ : std_logic;
signal \N__24744\ : std_logic;
signal \N__24743\ : std_logic;
signal \N__24742\ : std_logic;
signal \N__24741\ : std_logic;
signal \N__24738\ : std_logic;
signal \N__24735\ : std_logic;
signal \N__24732\ : std_logic;
signal \N__24729\ : std_logic;
signal \N__24726\ : std_logic;
signal \N__24723\ : std_logic;
signal \N__24720\ : std_logic;
signal \N__24717\ : std_logic;
signal \N__24716\ : std_logic;
signal \N__24713\ : std_logic;
signal \N__24712\ : std_logic;
signal \N__24709\ : std_logic;
signal \N__24706\ : std_logic;
signal \N__24703\ : std_logic;
signal \N__24700\ : std_logic;
signal \N__24697\ : std_logic;
signal \N__24694\ : std_logic;
signal \N__24691\ : std_logic;
signal \N__24690\ : std_logic;
signal \N__24687\ : std_logic;
signal \N__24682\ : std_logic;
signal \N__24679\ : std_logic;
signal \N__24674\ : std_logic;
signal \N__24671\ : std_logic;
signal \N__24668\ : std_logic;
signal \N__24665\ : std_logic;
signal \N__24660\ : std_logic;
signal \N__24651\ : std_logic;
signal \N__24644\ : std_logic;
signal \N__24641\ : std_logic;
signal \N__24634\ : std_logic;
signal \N__24629\ : std_logic;
signal \N__24624\ : std_logic;
signal \N__24617\ : std_logic;
signal \N__24614\ : std_logic;
signal \N__24611\ : std_logic;
signal \N__24608\ : std_logic;
signal \N__24605\ : std_logic;
signal \N__24602\ : std_logic;
signal \N__24599\ : std_logic;
signal \N__24596\ : std_logic;
signal \N__24587\ : std_logic;
signal \N__24582\ : std_logic;
signal \N__24579\ : std_logic;
signal \N__24578\ : std_logic;
signal \N__24577\ : std_logic;
signal \N__24570\ : std_logic;
signal \N__24569\ : std_logic;
signal \N__24566\ : std_logic;
signal \N__24563\ : std_logic;
signal \N__24558\ : std_logic;
signal \N__24555\ : std_logic;
signal \N__24554\ : std_logic;
signal \N__24551\ : std_logic;
signal \N__24550\ : std_logic;
signal \N__24547\ : std_logic;
signal \N__24544\ : std_logic;
signal \N__24541\ : std_logic;
signal \N__24534\ : std_logic;
signal \N__24533\ : std_logic;
signal \N__24530\ : std_logic;
signal \N__24529\ : std_logic;
signal \N__24528\ : std_logic;
signal \N__24525\ : std_logic;
signal \N__24524\ : std_logic;
signal \N__24517\ : std_logic;
signal \N__24514\ : std_logic;
signal \N__24511\ : std_logic;
signal \N__24508\ : std_logic;
signal \N__24507\ : std_logic;
signal \N__24504\ : std_logic;
signal \N__24501\ : std_logic;
signal \N__24500\ : std_logic;
signal \N__24497\ : std_logic;
signal \N__24494\ : std_logic;
signal \N__24491\ : std_logic;
signal \N__24488\ : std_logic;
signal \N__24487\ : std_logic;
signal \N__24486\ : std_logic;
signal \N__24483\ : std_logic;
signal \N__24480\ : std_logic;
signal \N__24477\ : std_logic;
signal \N__24474\ : std_logic;
signal \N__24471\ : std_logic;
signal \N__24468\ : std_logic;
signal \N__24467\ : std_logic;
signal \N__24464\ : std_logic;
signal \N__24463\ : std_logic;
signal \N__24462\ : std_logic;
signal \N__24457\ : std_logic;
signal \N__24452\ : std_logic;
signal \N__24449\ : std_logic;
signal \N__24446\ : std_logic;
signal \N__24443\ : std_logic;
signal \N__24440\ : std_logic;
signal \N__24435\ : std_logic;
signal \N__24432\ : std_logic;
signal \N__24429\ : std_logic;
signal \N__24426\ : std_logic;
signal \N__24411\ : std_logic;
signal \N__24408\ : std_logic;
signal \N__24407\ : std_logic;
signal \N__24406\ : std_logic;
signal \N__24405\ : std_logic;
signal \N__24402\ : std_logic;
signal \N__24401\ : std_logic;
signal \N__24398\ : std_logic;
signal \N__24395\ : std_logic;
signal \N__24394\ : std_logic;
signal \N__24393\ : std_logic;
signal \N__24390\ : std_logic;
signal \N__24387\ : std_logic;
signal \N__24384\ : std_logic;
signal \N__24379\ : std_logic;
signal \N__24374\ : std_logic;
signal \N__24371\ : std_logic;
signal \N__24360\ : std_logic;
signal \N__24357\ : std_logic;
signal \N__24354\ : std_logic;
signal \N__24351\ : std_logic;
signal \N__24348\ : std_logic;
signal \N__24347\ : std_logic;
signal \N__24346\ : std_logic;
signal \N__24345\ : std_logic;
signal \N__24342\ : std_logic;
signal \N__24339\ : std_logic;
signal \N__24336\ : std_logic;
signal \N__24333\ : std_logic;
signal \N__24330\ : std_logic;
signal \N__24321\ : std_logic;
signal \N__24318\ : std_logic;
signal \N__24315\ : std_logic;
signal \N__24312\ : std_logic;
signal \N__24309\ : std_logic;
signal \N__24306\ : std_logic;
signal \N__24303\ : std_logic;
signal \N__24300\ : std_logic;
signal \N__24299\ : std_logic;
signal \N__24298\ : std_logic;
signal \N__24295\ : std_logic;
signal \N__24292\ : std_logic;
signal \N__24289\ : std_logic;
signal \N__24286\ : std_logic;
signal \N__24279\ : std_logic;
signal \N__24276\ : std_logic;
signal \N__24273\ : std_logic;
signal \N__24270\ : std_logic;
signal \N__24267\ : std_logic;
signal \N__24264\ : std_logic;
signal \N__24261\ : std_logic;
signal \N__24260\ : std_logic;
signal \N__24259\ : std_logic;
signal \N__24258\ : std_logic;
signal \N__24257\ : std_logic;
signal \N__24256\ : std_logic;
signal \N__24255\ : std_logic;
signal \N__24254\ : std_logic;
signal \N__24253\ : std_logic;
signal \N__24250\ : std_logic;
signal \N__24247\ : std_logic;
signal \N__24240\ : std_logic;
signal \N__24237\ : std_logic;
signal \N__24236\ : std_logic;
signal \N__24235\ : std_logic;
signal \N__24232\ : std_logic;
signal \N__24229\ : std_logic;
signal \N__24226\ : std_logic;
signal \N__24225\ : std_logic;
signal \N__24222\ : std_logic;
signal \N__24219\ : std_logic;
signal \N__24216\ : std_logic;
signal \N__24213\ : std_logic;
signal \N__24208\ : std_logic;
signal \N__24203\ : std_logic;
signal \N__24200\ : std_logic;
signal \N__24197\ : std_logic;
signal \N__24194\ : std_logic;
signal \N__24191\ : std_logic;
signal \N__24188\ : std_logic;
signal \N__24185\ : std_logic;
signal \N__24178\ : std_logic;
signal \N__24165\ : std_logic;
signal \N__24162\ : std_logic;
signal \N__24161\ : std_logic;
signal \N__24158\ : std_logic;
signal \N__24157\ : std_logic;
signal \N__24154\ : std_logic;
signal \N__24151\ : std_logic;
signal \N__24148\ : std_logic;
signal \N__24147\ : std_logic;
signal \N__24144\ : std_logic;
signal \N__24139\ : std_logic;
signal \N__24136\ : std_logic;
signal \N__24131\ : std_logic;
signal \N__24126\ : std_logic;
signal \N__24125\ : std_logic;
signal \N__24122\ : std_logic;
signal \N__24119\ : std_logic;
signal \N__24118\ : std_logic;
signal \N__24117\ : std_logic;
signal \N__24116\ : std_logic;
signal \N__24113\ : std_logic;
signal \N__24108\ : std_logic;
signal \N__24103\ : std_logic;
signal \N__24096\ : std_logic;
signal \N__24093\ : std_logic;
signal \N__24090\ : std_logic;
signal \N__24089\ : std_logic;
signal \N__24088\ : std_logic;
signal \N__24087\ : std_logic;
signal \N__24086\ : std_logic;
signal \N__24085\ : std_logic;
signal \N__24082\ : std_logic;
signal \N__24079\ : std_logic;
signal \N__24078\ : std_logic;
signal \N__24077\ : std_logic;
signal \N__24074\ : std_logic;
signal \N__24073\ : std_logic;
signal \N__24070\ : std_logic;
signal \N__24069\ : std_logic;
signal \N__24068\ : std_logic;
signal \N__24067\ : std_logic;
signal \N__24066\ : std_logic;
signal \N__24063\ : std_logic;
signal \N__24060\ : std_logic;
signal \N__24057\ : std_logic;
signal \N__24056\ : std_logic;
signal \N__24053\ : std_logic;
signal \N__24050\ : std_logic;
signal \N__24041\ : std_logic;
signal \N__24032\ : std_logic;
signal \N__24029\ : std_logic;
signal \N__24026\ : std_logic;
signal \N__24025\ : std_logic;
signal \N__24024\ : std_logic;
signal \N__24021\ : std_logic;
signal \N__24018\ : std_logic;
signal \N__24017\ : std_logic;
signal \N__24014\ : std_logic;
signal \N__24011\ : std_logic;
signal \N__24006\ : std_logic;
signal \N__24005\ : std_logic;
signal \N__24004\ : std_logic;
signal \N__24003\ : std_logic;
signal \N__24002\ : std_logic;
signal \N__23999\ : std_logic;
signal \N__23996\ : std_logic;
signal \N__23991\ : std_logic;
signal \N__23986\ : std_logic;
signal \N__23983\ : std_logic;
signal \N__23982\ : std_logic;
signal \N__23981\ : std_logic;
signal \N__23980\ : std_logic;
signal \N__23977\ : std_logic;
signal \N__23972\ : std_logic;
signal \N__23969\ : std_logic;
signal \N__23966\ : std_logic;
signal \N__23963\ : std_logic;
signal \N__23962\ : std_logic;
signal \N__23961\ : std_logic;
signal \N__23960\ : std_logic;
signal \N__23959\ : std_logic;
signal \N__23956\ : std_logic;
signal \N__23947\ : std_logic;
signal \N__23944\ : std_logic;
signal \N__23937\ : std_logic;
signal \N__23934\ : std_logic;
signal \N__23931\ : std_logic;
signal \N__23928\ : std_logic;
signal \N__23925\ : std_logic;
signal \N__23920\ : std_logic;
signal \N__23911\ : std_logic;
signal \N__23908\ : std_logic;
signal \N__23889\ : std_logic;
signal \N__23886\ : std_logic;
signal \N__23883\ : std_logic;
signal \N__23882\ : std_logic;
signal \N__23881\ : std_logic;
signal \N__23880\ : std_logic;
signal \N__23879\ : std_logic;
signal \N__23878\ : std_logic;
signal \N__23877\ : std_logic;
signal \N__23876\ : std_logic;
signal \N__23875\ : std_logic;
signal \N__23874\ : std_logic;
signal \N__23873\ : std_logic;
signal \N__23872\ : std_logic;
signal \N__23871\ : std_logic;
signal \N__23870\ : std_logic;
signal \N__23869\ : std_logic;
signal \N__23868\ : std_logic;
signal \N__23867\ : std_logic;
signal \N__23866\ : std_logic;
signal \N__23865\ : std_logic;
signal \N__23864\ : std_logic;
signal \N__23863\ : std_logic;
signal \N__23862\ : std_logic;
signal \N__23861\ : std_logic;
signal \N__23860\ : std_logic;
signal \N__23859\ : std_logic;
signal \N__23858\ : std_logic;
signal \N__23857\ : std_logic;
signal \N__23856\ : std_logic;
signal \N__23855\ : std_logic;
signal \N__23854\ : std_logic;
signal \N__23853\ : std_logic;
signal \N__23852\ : std_logic;
signal \N__23851\ : std_logic;
signal \N__23850\ : std_logic;
signal \N__23849\ : std_logic;
signal \N__23848\ : std_logic;
signal \N__23847\ : std_logic;
signal \N__23846\ : std_logic;
signal \N__23845\ : std_logic;
signal \N__23844\ : std_logic;
signal \N__23843\ : std_logic;
signal \N__23842\ : std_logic;
signal \N__23841\ : std_logic;
signal \N__23840\ : std_logic;
signal \N__23839\ : std_logic;
signal \N__23838\ : std_logic;
signal \N__23837\ : std_logic;
signal \N__23836\ : std_logic;
signal \N__23835\ : std_logic;
signal \N__23834\ : std_logic;
signal \N__23833\ : std_logic;
signal \N__23832\ : std_logic;
signal \N__23831\ : std_logic;
signal \N__23830\ : std_logic;
signal \N__23829\ : std_logic;
signal \N__23828\ : std_logic;
signal \N__23827\ : std_logic;
signal \N__23826\ : std_logic;
signal \N__23825\ : std_logic;
signal \N__23824\ : std_logic;
signal \N__23823\ : std_logic;
signal \N__23822\ : std_logic;
signal \N__23821\ : std_logic;
signal \N__23820\ : std_logic;
signal \N__23819\ : std_logic;
signal \N__23818\ : std_logic;
signal \N__23817\ : std_logic;
signal \N__23816\ : std_logic;
signal \N__23815\ : std_logic;
signal \N__23814\ : std_logic;
signal \N__23813\ : std_logic;
signal \N__23812\ : std_logic;
signal \N__23811\ : std_logic;
signal \N__23810\ : std_logic;
signal \N__23809\ : std_logic;
signal \N__23808\ : std_logic;
signal \N__23807\ : std_logic;
signal \N__23806\ : std_logic;
signal \N__23805\ : std_logic;
signal \N__23804\ : std_logic;
signal \N__23803\ : std_logic;
signal \N__23802\ : std_logic;
signal \N__23801\ : std_logic;
signal \N__23800\ : std_logic;
signal \N__23799\ : std_logic;
signal \N__23798\ : std_logic;
signal \N__23797\ : std_logic;
signal \N__23796\ : std_logic;
signal \N__23795\ : std_logic;
signal \N__23794\ : std_logic;
signal \N__23793\ : std_logic;
signal \N__23792\ : std_logic;
signal \N__23791\ : std_logic;
signal \N__23790\ : std_logic;
signal \N__23789\ : std_logic;
signal \N__23788\ : std_logic;
signal \N__23787\ : std_logic;
signal \N__23786\ : std_logic;
signal \N__23785\ : std_logic;
signal \N__23784\ : std_logic;
signal \N__23783\ : std_logic;
signal \N__23782\ : std_logic;
signal \N__23577\ : std_logic;
signal \N__23574\ : std_logic;
signal \N__23571\ : std_logic;
signal \N__23570\ : std_logic;
signal \N__23569\ : std_logic;
signal \N__23568\ : std_logic;
signal \N__23567\ : std_logic;
signal \N__23566\ : std_logic;
signal \N__23565\ : std_logic;
signal \N__23564\ : std_logic;
signal \N__23563\ : std_logic;
signal \N__23562\ : std_logic;
signal \N__23541\ : std_logic;
signal \N__23538\ : std_logic;
signal \N__23535\ : std_logic;
signal \N__23534\ : std_logic;
signal \N__23533\ : std_logic;
signal \N__23532\ : std_logic;
signal \N__23531\ : std_logic;
signal \N__23530\ : std_logic;
signal \N__23527\ : std_logic;
signal \N__23524\ : std_logic;
signal \N__23523\ : std_logic;
signal \N__23522\ : std_logic;
signal \N__23521\ : std_logic;
signal \N__23520\ : std_logic;
signal \N__23517\ : std_logic;
signal \N__23514\ : std_logic;
signal \N__23513\ : std_logic;
signal \N__23512\ : std_logic;
signal \N__23511\ : std_logic;
signal \N__23508\ : std_logic;
signal \N__23507\ : std_logic;
signal \N__23506\ : std_logic;
signal \N__23505\ : std_logic;
signal \N__23504\ : std_logic;
signal \N__23503\ : std_logic;
signal \N__23502\ : std_logic;
signal \N__23501\ : std_logic;
signal \N__23500\ : std_logic;
signal \N__23499\ : std_logic;
signal \N__23498\ : std_logic;
signal \N__23497\ : std_logic;
signal \N__23496\ : std_logic;
signal \N__23495\ : std_logic;
signal \N__23494\ : std_logic;
signal \N__23493\ : std_logic;
signal \N__23492\ : std_logic;
signal \N__23491\ : std_logic;
signal \N__23490\ : std_logic;
signal \N__23487\ : std_logic;
signal \N__23482\ : std_logic;
signal \N__23479\ : std_logic;
signal \N__23476\ : std_logic;
signal \N__23473\ : std_logic;
signal \N__23470\ : std_logic;
signal \N__23463\ : std_logic;
signal \N__23460\ : std_logic;
signal \N__23457\ : std_logic;
signal \N__23450\ : std_logic;
signal \N__23445\ : std_logic;
signal \N__23442\ : std_logic;
signal \N__23439\ : std_logic;
signal \N__23436\ : std_logic;
signal \N__23433\ : std_logic;
signal \N__23428\ : std_logic;
signal \N__23425\ : std_logic;
signal \N__23422\ : std_logic;
signal \N__23415\ : std_logic;
signal \N__23412\ : std_logic;
signal \N__23409\ : std_logic;
signal \N__23406\ : std_logic;
signal \N__23405\ : std_logic;
signal \N__23404\ : std_logic;
signal \N__23403\ : std_logic;
signal \N__23402\ : std_logic;
signal \N__23401\ : std_logic;
signal \N__23400\ : std_logic;
signal \N__23399\ : std_logic;
signal \N__23398\ : std_logic;
signal \N__23397\ : std_logic;
signal \N__23396\ : std_logic;
signal \N__23395\ : std_logic;
signal \N__23394\ : std_logic;
signal \N__23393\ : std_logic;
signal \N__23392\ : std_logic;
signal \N__23391\ : std_logic;
signal \N__23390\ : std_logic;
signal \N__23389\ : std_logic;
signal \N__23388\ : std_logic;
signal \N__23387\ : std_logic;
signal \N__23386\ : std_logic;
signal \N__23385\ : std_logic;
signal \N__23384\ : std_logic;
signal \N__23383\ : std_logic;
signal \N__23382\ : std_logic;
signal \N__23381\ : std_logic;
signal \N__23380\ : std_logic;
signal \N__23379\ : std_logic;
signal \N__23378\ : std_logic;
signal \N__23377\ : std_logic;
signal \N__23376\ : std_logic;
signal \N__23375\ : std_logic;
signal \N__23374\ : std_logic;
signal \N__23373\ : std_logic;
signal \N__23372\ : std_logic;
signal \N__23371\ : std_logic;
signal \N__23370\ : std_logic;
signal \N__23369\ : std_logic;
signal \N__23368\ : std_logic;
signal \N__23367\ : std_logic;
signal \N__23366\ : std_logic;
signal \N__23365\ : std_logic;
signal \N__23364\ : std_logic;
signal \N__23363\ : std_logic;
signal \N__23362\ : std_logic;
signal \N__23361\ : std_logic;
signal \N__23360\ : std_logic;
signal \N__23359\ : std_logic;
signal \N__23358\ : std_logic;
signal \N__23357\ : std_logic;
signal \N__23356\ : std_logic;
signal \N__23355\ : std_logic;
signal \N__23354\ : std_logic;
signal \N__23353\ : std_logic;
signal \N__23352\ : std_logic;
signal \N__23351\ : std_logic;
signal \N__23350\ : std_logic;
signal \N__23349\ : std_logic;
signal \N__23348\ : std_logic;
signal \N__23347\ : std_logic;
signal \N__23346\ : std_logic;
signal \N__23345\ : std_logic;
signal \N__23344\ : std_logic;
signal \N__23343\ : std_logic;
signal \N__23342\ : std_logic;
signal \N__23341\ : std_logic;
signal \N__23338\ : std_logic;
signal \N__23335\ : std_logic;
signal \N__23332\ : std_logic;
signal \N__23329\ : std_logic;
signal \N__23326\ : std_logic;
signal \N__23323\ : std_logic;
signal \N__23320\ : std_logic;
signal \N__23317\ : std_logic;
signal \N__23314\ : std_logic;
signal \N__23311\ : std_logic;
signal \N__23308\ : std_logic;
signal \N__23305\ : std_logic;
signal \N__23302\ : std_logic;
signal \N__23299\ : std_logic;
signal \N__23296\ : std_logic;
signal \N__23293\ : std_logic;
signal \N__23290\ : std_logic;
signal \N__23287\ : std_logic;
signal \N__23284\ : std_logic;
signal \N__23281\ : std_logic;
signal \N__23278\ : std_logic;
signal \N__23275\ : std_logic;
signal \N__23100\ : std_logic;
signal \N__23097\ : std_logic;
signal \N__23094\ : std_logic;
signal \N__23091\ : std_logic;
signal \N__23088\ : std_logic;
signal \N__23085\ : std_logic;
signal \N__23082\ : std_logic;
signal \N__23079\ : std_logic;
signal \N__23076\ : std_logic;
signal \N__23073\ : std_logic;
signal \N__23070\ : std_logic;
signal \N__23067\ : std_logic;
signal \N__23064\ : std_logic;
signal \N__23061\ : std_logic;
signal \N__23058\ : std_logic;
signal \N__23055\ : std_logic;
signal \N__23052\ : std_logic;
signal \N__23049\ : std_logic;
signal \N__23046\ : std_logic;
signal \N__23043\ : std_logic;
signal \N__23040\ : std_logic;
signal \N__23037\ : std_logic;
signal \N__23034\ : std_logic;
signal \N__23031\ : std_logic;
signal \N__23028\ : std_logic;
signal \N__23025\ : std_logic;
signal \N__23022\ : std_logic;
signal \N__23019\ : std_logic;
signal \N__23018\ : std_logic;
signal \N__23017\ : std_logic;
signal \N__23014\ : std_logic;
signal \N__23009\ : std_logic;
signal \N__23004\ : std_logic;
signal \N__23001\ : std_logic;
signal \N__22998\ : std_logic;
signal \N__22995\ : std_logic;
signal \N__22994\ : std_logic;
signal \N__22991\ : std_logic;
signal \N__22990\ : std_logic;
signal \N__22987\ : std_logic;
signal \N__22984\ : std_logic;
signal \N__22981\ : std_logic;
signal \N__22974\ : std_logic;
signal \N__22971\ : std_logic;
signal \N__22968\ : std_logic;
signal \N__22967\ : std_logic;
signal \N__22966\ : std_logic;
signal \N__22963\ : std_logic;
signal \N__22960\ : std_logic;
signal \N__22957\ : std_logic;
signal \N__22950\ : std_logic;
signal \N__22947\ : std_logic;
signal \N__22944\ : std_logic;
signal \N__22941\ : std_logic;
signal \N__22938\ : std_logic;
signal \N__22937\ : std_logic;
signal \N__22936\ : std_logic;
signal \N__22933\ : std_logic;
signal \N__22930\ : std_logic;
signal \N__22927\ : std_logic;
signal \N__22920\ : std_logic;
signal \N__22917\ : std_logic;
signal \N__22914\ : std_logic;
signal \N__22911\ : std_logic;
signal \N__22908\ : std_logic;
signal \N__22905\ : std_logic;
signal \N__22902\ : std_logic;
signal \N__22899\ : std_logic;
signal \N__22896\ : std_logic;
signal \N__22895\ : std_logic;
signal \N__22892\ : std_logic;
signal \N__22889\ : std_logic;
signal \N__22886\ : std_logic;
signal \N__22883\ : std_logic;
signal \N__22880\ : std_logic;
signal \N__22877\ : std_logic;
signal \N__22872\ : std_logic;
signal \N__22869\ : std_logic;
signal \N__22868\ : std_logic;
signal \N__22863\ : std_logic;
signal \N__22862\ : std_logic;
signal \N__22859\ : std_logic;
signal \N__22856\ : std_logic;
signal \N__22851\ : std_logic;
signal \N__22848\ : std_logic;
signal \N__22845\ : std_logic;
signal \N__22842\ : std_logic;
signal \N__22841\ : std_logic;
signal \N__22840\ : std_logic;
signal \N__22839\ : std_logic;
signal \N__22838\ : std_logic;
signal \N__22837\ : std_logic;
signal \N__22836\ : std_logic;
signal \N__22835\ : std_logic;
signal \N__22832\ : std_logic;
signal \N__22825\ : std_logic;
signal \N__22822\ : std_logic;
signal \N__22819\ : std_logic;
signal \N__22814\ : std_logic;
signal \N__22803\ : std_logic;
signal \N__22800\ : std_logic;
signal \N__22797\ : std_logic;
signal \N__22794\ : std_logic;
signal \N__22791\ : std_logic;
signal \N__22788\ : std_logic;
signal \N__22787\ : std_logic;
signal \N__22784\ : std_logic;
signal \N__22781\ : std_logic;
signal \N__22776\ : std_logic;
signal \N__22773\ : std_logic;
signal \N__22770\ : std_logic;
signal \N__22767\ : std_logic;
signal \N__22766\ : std_logic;
signal \N__22763\ : std_logic;
signal \N__22762\ : std_logic;
signal \N__22759\ : std_logic;
signal \N__22756\ : std_logic;
signal \N__22753\ : std_logic;
signal \N__22746\ : std_logic;
signal \N__22743\ : std_logic;
signal \N__22740\ : std_logic;
signal \N__22737\ : std_logic;
signal \N__22734\ : std_logic;
signal \N__22733\ : std_logic;
signal \N__22732\ : std_logic;
signal \N__22729\ : std_logic;
signal \N__22726\ : std_logic;
signal \N__22723\ : std_logic;
signal \N__22716\ : std_logic;
signal \N__22713\ : std_logic;
signal \N__22710\ : std_logic;
signal \N__22707\ : std_logic;
signal \N__22704\ : std_logic;
signal \N__22703\ : std_logic;
signal \N__22702\ : std_logic;
signal \N__22699\ : std_logic;
signal \N__22696\ : std_logic;
signal \N__22693\ : std_logic;
signal \N__22692\ : std_logic;
signal \N__22689\ : std_logic;
signal \N__22684\ : std_logic;
signal \N__22681\ : std_logic;
signal \N__22676\ : std_logic;
signal \N__22673\ : std_logic;
signal \N__22670\ : std_logic;
signal \N__22667\ : std_logic;
signal \N__22664\ : std_logic;
signal \N__22661\ : std_logic;
signal \N__22656\ : std_logic;
signal \N__22653\ : std_logic;
signal \N__22650\ : std_logic;
signal \N__22647\ : std_logic;
signal \N__22644\ : std_logic;
signal \N__22641\ : std_logic;
signal \N__22640\ : std_logic;
signal \N__22639\ : std_logic;
signal \N__22636\ : std_logic;
signal \N__22633\ : std_logic;
signal \N__22632\ : std_logic;
signal \N__22629\ : std_logic;
signal \N__22626\ : std_logic;
signal \N__22623\ : std_logic;
signal \N__22620\ : std_logic;
signal \N__22617\ : std_logic;
signal \N__22608\ : std_logic;
signal \N__22605\ : std_logic;
signal \N__22602\ : std_logic;
signal \N__22599\ : std_logic;
signal \N__22596\ : std_logic;
signal \N__22593\ : std_logic;
signal \N__22590\ : std_logic;
signal \N__22587\ : std_logic;
signal \N__22584\ : std_logic;
signal \N__22581\ : std_logic;
signal \N__22578\ : std_logic;
signal \N__22577\ : std_logic;
signal \N__22576\ : std_logic;
signal \N__22573\ : std_logic;
signal \N__22570\ : std_logic;
signal \N__22569\ : std_logic;
signal \N__22566\ : std_logic;
signal \N__22563\ : std_logic;
signal \N__22560\ : std_logic;
signal \N__22557\ : std_logic;
signal \N__22554\ : std_logic;
signal \N__22549\ : std_logic;
signal \N__22544\ : std_logic;
signal \N__22539\ : std_logic;
signal \N__22536\ : std_logic;
signal \N__22533\ : std_logic;
signal \N__22530\ : std_logic;
signal \N__22527\ : std_logic;
signal \N__22526\ : std_logic;
signal \N__22525\ : std_logic;
signal \N__22522\ : std_logic;
signal \N__22519\ : std_logic;
signal \N__22516\ : std_logic;
signal \N__22513\ : std_logic;
signal \N__22512\ : std_logic;
signal \N__22509\ : std_logic;
signal \N__22506\ : std_logic;
signal \N__22503\ : std_logic;
signal \N__22500\ : std_logic;
signal \N__22495\ : std_logic;
signal \N__22488\ : std_logic;
signal \N__22485\ : std_logic;
signal \N__22482\ : std_logic;
signal \N__22479\ : std_logic;
signal \N__22476\ : std_logic;
signal \N__22473\ : std_logic;
signal \N__22470\ : std_logic;
signal \N__22469\ : std_logic;
signal \N__22468\ : std_logic;
signal \N__22465\ : std_logic;
signal \N__22462\ : std_logic;
signal \N__22461\ : std_logic;
signal \N__22458\ : std_logic;
signal \N__22455\ : std_logic;
signal \N__22452\ : std_logic;
signal \N__22449\ : std_logic;
signal \N__22440\ : std_logic;
signal \N__22437\ : std_logic;
signal \N__22434\ : std_logic;
signal \N__22431\ : std_logic;
signal \N__22428\ : std_logic;
signal \N__22427\ : std_logic;
signal \N__22424\ : std_logic;
signal \N__22423\ : std_logic;
signal \N__22420\ : std_logic;
signal \N__22417\ : std_logic;
signal \N__22414\ : std_logic;
signal \N__22407\ : std_logic;
signal \N__22404\ : std_logic;
signal \N__22401\ : std_logic;
signal \N__22398\ : std_logic;
signal \N__22395\ : std_logic;
signal \N__22392\ : std_logic;
signal \N__22389\ : std_logic;
signal \N__22386\ : std_logic;
signal \N__22385\ : std_logic;
signal \N__22384\ : std_logic;
signal \N__22381\ : std_logic;
signal \N__22378\ : std_logic;
signal \N__22375\ : std_logic;
signal \N__22368\ : std_logic;
signal \N__22367\ : std_logic;
signal \N__22366\ : std_logic;
signal \N__22363\ : std_logic;
signal \N__22360\ : std_logic;
signal \N__22357\ : std_logic;
signal \N__22350\ : std_logic;
signal \N__22349\ : std_logic;
signal \N__22346\ : std_logic;
signal \N__22345\ : std_logic;
signal \N__22342\ : std_logic;
signal \N__22339\ : std_logic;
signal \N__22336\ : std_logic;
signal \N__22329\ : std_logic;
signal \N__22328\ : std_logic;
signal \N__22327\ : std_logic;
signal \N__22324\ : std_logic;
signal \N__22321\ : std_logic;
signal \N__22318\ : std_logic;
signal \N__22311\ : std_logic;
signal \N__22310\ : std_logic;
signal \N__22307\ : std_logic;
signal \N__22304\ : std_logic;
signal \N__22303\ : std_logic;
signal \N__22300\ : std_logic;
signal \N__22297\ : std_logic;
signal \N__22294\ : std_logic;
signal \N__22287\ : std_logic;
signal \N__22284\ : std_logic;
signal \N__22283\ : std_logic;
signal \N__22280\ : std_logic;
signal \N__22279\ : std_logic;
signal \N__22276\ : std_logic;
signal \N__22273\ : std_logic;
signal \N__22270\ : std_logic;
signal \N__22269\ : std_logic;
signal \N__22266\ : std_logic;
signal \N__22263\ : std_logic;
signal \N__22258\ : std_logic;
signal \N__22251\ : std_logic;
signal \N__22248\ : std_logic;
signal \N__22245\ : std_logic;
signal \N__22242\ : std_logic;
signal \N__22239\ : std_logic;
signal \N__22236\ : std_logic;
signal \N__22235\ : std_logic;
signal \N__22232\ : std_logic;
signal \N__22231\ : std_logic;
signal \N__22228\ : std_logic;
signal \N__22225\ : std_logic;
signal \N__22222\ : std_logic;
signal \N__22219\ : std_logic;
signal \N__22216\ : std_logic;
signal \N__22213\ : std_logic;
signal \N__22210\ : std_logic;
signal \N__22207\ : std_logic;
signal \N__22204\ : std_logic;
signal \N__22201\ : std_logic;
signal \N__22194\ : std_logic;
signal \N__22191\ : std_logic;
signal \N__22188\ : std_logic;
signal \N__22187\ : std_logic;
signal \N__22186\ : std_logic;
signal \N__22185\ : std_logic;
signal \N__22182\ : std_logic;
signal \N__22179\ : std_logic;
signal \N__22176\ : std_logic;
signal \N__22173\ : std_logic;
signal \N__22164\ : std_logic;
signal \N__22161\ : std_logic;
signal \N__22158\ : std_logic;
signal \N__22155\ : std_logic;
signal \N__22154\ : std_logic;
signal \N__22151\ : std_logic;
signal \N__22150\ : std_logic;
signal \N__22147\ : std_logic;
signal \N__22144\ : std_logic;
signal \N__22141\ : std_logic;
signal \N__22134\ : std_logic;
signal \N__22133\ : std_logic;
signal \N__22132\ : std_logic;
signal \N__22129\ : std_logic;
signal \N__22126\ : std_logic;
signal \N__22125\ : std_logic;
signal \N__22124\ : std_logic;
signal \N__22123\ : std_logic;
signal \N__22122\ : std_logic;
signal \N__22121\ : std_logic;
signal \N__22120\ : std_logic;
signal \N__22119\ : std_logic;
signal \N__22118\ : std_logic;
signal \N__22117\ : std_logic;
signal \N__22116\ : std_logic;
signal \N__22111\ : std_logic;
signal \N__22110\ : std_logic;
signal \N__22105\ : std_logic;
signal \N__22102\ : std_logic;
signal \N__22099\ : std_logic;
signal \N__22098\ : std_logic;
signal \N__22097\ : std_logic;
signal \N__22096\ : std_logic;
signal \N__22091\ : std_logic;
signal \N__22084\ : std_logic;
signal \N__22079\ : std_logic;
signal \N__22076\ : std_logic;
signal \N__22073\ : std_logic;
signal \N__22072\ : std_logic;
signal \N__22069\ : std_logic;
signal \N__22068\ : std_logic;
signal \N__22063\ : std_logic;
signal \N__22060\ : std_logic;
signal \N__22059\ : std_logic;
signal \N__22058\ : std_logic;
signal \N__22053\ : std_logic;
signal \N__22050\ : std_logic;
signal \N__22045\ : std_logic;
signal \N__22042\ : std_logic;
signal \N__22039\ : std_logic;
signal \N__22036\ : std_logic;
signal \N__22033\ : std_logic;
signal \N__22030\ : std_logic;
signal \N__22027\ : std_logic;
signal \N__22020\ : std_logic;
signal \N__22015\ : std_logic;
signal \N__22008\ : std_logic;
signal \N__21993\ : std_logic;
signal \N__21992\ : std_logic;
signal \N__21991\ : std_logic;
signal \N__21990\ : std_logic;
signal \N__21989\ : std_logic;
signal \N__21982\ : std_logic;
signal \N__21981\ : std_logic;
signal \N__21980\ : std_logic;
signal \N__21979\ : std_logic;
signal \N__21978\ : std_logic;
signal \N__21977\ : std_logic;
signal \N__21976\ : std_logic;
signal \N__21975\ : std_logic;
signal \N__21974\ : std_logic;
signal \N__21973\ : std_logic;
signal \N__21968\ : std_logic;
signal \N__21967\ : std_logic;
signal \N__21966\ : std_logic;
signal \N__21965\ : std_logic;
signal \N__21964\ : std_logic;
signal \N__21961\ : std_logic;
signal \N__21954\ : std_logic;
signal \N__21951\ : std_logic;
signal \N__21948\ : std_logic;
signal \N__21943\ : std_logic;
signal \N__21942\ : std_logic;
signal \N__21939\ : std_logic;
signal \N__21936\ : std_logic;
signal \N__21933\ : std_logic;
signal \N__21930\ : std_logic;
signal \N__21929\ : std_logic;
signal \N__21928\ : std_logic;
signal \N__21925\ : std_logic;
signal \N__21920\ : std_logic;
signal \N__21915\ : std_logic;
signal \N__21908\ : std_logic;
signal \N__21907\ : std_logic;
signal \N__21904\ : std_logic;
signal \N__21901\ : std_logic;
signal \N__21896\ : std_logic;
signal \N__21893\ : std_logic;
signal \N__21888\ : std_logic;
signal \N__21883\ : std_logic;
signal \N__21882\ : std_logic;
signal \N__21881\ : std_logic;
signal \N__21880\ : std_logic;
signal \N__21875\ : std_logic;
signal \N__21872\ : std_logic;
signal \N__21869\ : std_logic;
signal \N__21864\ : std_logic;
signal \N__21861\ : std_logic;
signal \N__21856\ : std_logic;
signal \N__21849\ : std_logic;
signal \N__21844\ : std_logic;
signal \N__21831\ : std_logic;
signal \N__21830\ : std_logic;
signal \N__21827\ : std_logic;
signal \N__21824\ : std_logic;
signal \N__21821\ : std_logic;
signal \N__21818\ : std_logic;
signal \N__21817\ : std_logic;
signal \N__21814\ : std_logic;
signal \N__21813\ : std_logic;
signal \N__21810\ : std_logic;
signal \N__21807\ : std_logic;
signal \N__21804\ : std_logic;
signal \N__21801\ : std_logic;
signal \N__21798\ : std_logic;
signal \N__21795\ : std_logic;
signal \N__21786\ : std_logic;
signal \N__21785\ : std_logic;
signal \N__21782\ : std_logic;
signal \N__21781\ : std_logic;
signal \N__21780\ : std_logic;
signal \N__21779\ : std_logic;
signal \N__21778\ : std_logic;
signal \N__21777\ : std_logic;
signal \N__21776\ : std_logic;
signal \N__21775\ : std_logic;
signal \N__21774\ : std_logic;
signal \N__21773\ : std_logic;
signal \N__21772\ : std_logic;
signal \N__21769\ : std_logic;
signal \N__21766\ : std_logic;
signal \N__21763\ : std_logic;
signal \N__21762\ : std_logic;
signal \N__21761\ : std_logic;
signal \N__21760\ : std_logic;
signal \N__21753\ : std_logic;
signal \N__21744\ : std_logic;
signal \N__21741\ : std_logic;
signal \N__21738\ : std_logic;
signal \N__21735\ : std_logic;
signal \N__21734\ : std_logic;
signal \N__21733\ : std_logic;
signal \N__21730\ : std_logic;
signal \N__21727\ : std_logic;
signal \N__21722\ : std_logic;
signal \N__21719\ : std_logic;
signal \N__21716\ : std_logic;
signal \N__21713\ : std_logic;
signal \N__21710\ : std_logic;
signal \N__21707\ : std_logic;
signal \N__21704\ : std_logic;
signal \N__21703\ : std_logic;
signal \N__21702\ : std_logic;
signal \N__21699\ : std_logic;
signal \N__21696\ : std_logic;
signal \N__21691\ : std_logic;
signal \N__21688\ : std_logic;
signal \N__21687\ : std_logic;
signal \N__21686\ : std_logic;
signal \N__21685\ : std_logic;
signal \N__21684\ : std_logic;
signal \N__21679\ : std_logic;
signal \N__21676\ : std_logic;
signal \N__21669\ : std_logic;
signal \N__21666\ : std_logic;
signal \N__21659\ : std_logic;
signal \N__21654\ : std_logic;
signal \N__21651\ : std_logic;
signal \N__21644\ : std_logic;
signal \N__21637\ : std_logic;
signal \N__21624\ : std_logic;
signal \N__21623\ : std_logic;
signal \N__21622\ : std_logic;
signal \N__21621\ : std_logic;
signal \N__21620\ : std_logic;
signal \N__21619\ : std_logic;
signal \N__21618\ : std_logic;
signal \N__21615\ : std_logic;
signal \N__21614\ : std_logic;
signal \N__21611\ : std_logic;
signal \N__21610\ : std_logic;
signal \N__21609\ : std_logic;
signal \N__21606\ : std_logic;
signal \N__21603\ : std_logic;
signal \N__21602\ : std_logic;
signal \N__21599\ : std_logic;
signal \N__21594\ : std_logic;
signal \N__21585\ : std_logic;
signal \N__21582\ : std_logic;
signal \N__21579\ : std_logic;
signal \N__21576\ : std_logic;
signal \N__21571\ : std_logic;
signal \N__21566\ : std_logic;
signal \N__21563\ : std_logic;
signal \N__21558\ : std_logic;
signal \N__21555\ : std_logic;
signal \N__21552\ : std_logic;
signal \N__21545\ : std_logic;
signal \N__21540\ : std_logic;
signal \N__21539\ : std_logic;
signal \N__21536\ : std_logic;
signal \N__21533\ : std_logic;
signal \N__21530\ : std_logic;
signal \N__21527\ : std_logic;
signal \N__21524\ : std_logic;
signal \N__21521\ : std_logic;
signal \N__21518\ : std_logic;
signal \N__21513\ : std_logic;
signal \N__21512\ : std_logic;
signal \N__21511\ : std_logic;
signal \N__21508\ : std_logic;
signal \N__21507\ : std_logic;
signal \N__21504\ : std_logic;
signal \N__21501\ : std_logic;
signal \N__21498\ : std_logic;
signal \N__21495\ : std_logic;
signal \N__21492\ : std_logic;
signal \N__21489\ : std_logic;
signal \N__21484\ : std_logic;
signal \N__21481\ : std_logic;
signal \N__21476\ : std_logic;
signal \N__21471\ : std_logic;
signal \N__21468\ : std_logic;
signal \N__21465\ : std_logic;
signal \N__21462\ : std_logic;
signal \N__21461\ : std_logic;
signal \N__21458\ : std_logic;
signal \N__21455\ : std_logic;
signal \N__21450\ : std_logic;
signal \N__21449\ : std_logic;
signal \N__21446\ : std_logic;
signal \N__21445\ : std_logic;
signal \N__21442\ : std_logic;
signal \N__21439\ : std_logic;
signal \N__21436\ : std_logic;
signal \N__21429\ : std_logic;
signal \N__21426\ : std_logic;
signal \N__21423\ : std_logic;
signal \N__21422\ : std_logic;
signal \N__21421\ : std_logic;
signal \N__21414\ : std_logic;
signal \N__21411\ : std_logic;
signal \N__21408\ : std_logic;
signal \N__21407\ : std_logic;
signal \N__21404\ : std_logic;
signal \N__21401\ : std_logic;
signal \N__21398\ : std_logic;
signal \N__21395\ : std_logic;
signal \N__21394\ : std_logic;
signal \N__21389\ : std_logic;
signal \N__21386\ : std_logic;
signal \N__21381\ : std_logic;
signal \N__21378\ : std_logic;
signal \N__21375\ : std_logic;
signal \N__21372\ : std_logic;
signal \N__21369\ : std_logic;
signal \N__21366\ : std_logic;
signal \N__21363\ : std_logic;
signal \N__21360\ : std_logic;
signal \N__21357\ : std_logic;
signal \N__21354\ : std_logic;
signal \N__21351\ : std_logic;
signal \N__21350\ : std_logic;
signal \N__21349\ : std_logic;
signal \N__21346\ : std_logic;
signal \N__21343\ : std_logic;
signal \N__21340\ : std_logic;
signal \N__21337\ : std_logic;
signal \N__21336\ : std_logic;
signal \N__21333\ : std_logic;
signal \N__21330\ : std_logic;
signal \N__21327\ : std_logic;
signal \N__21324\ : std_logic;
signal \N__21321\ : std_logic;
signal \N__21318\ : std_logic;
signal \N__21315\ : std_logic;
signal \N__21312\ : std_logic;
signal \N__21303\ : std_logic;
signal \N__21300\ : std_logic;
signal \N__21297\ : std_logic;
signal \N__21294\ : std_logic;
signal \N__21291\ : std_logic;
signal \N__21288\ : std_logic;
signal \N__21287\ : std_logic;
signal \N__21284\ : std_logic;
signal \N__21281\ : std_logic;
signal \N__21276\ : std_logic;
signal \N__21273\ : std_logic;
signal \N__21272\ : std_logic;
signal \N__21271\ : std_logic;
signal \N__21268\ : std_logic;
signal \N__21265\ : std_logic;
signal \N__21262\ : std_logic;
signal \N__21259\ : std_logic;
signal \N__21256\ : std_logic;
signal \N__21253\ : std_logic;
signal \N__21248\ : std_logic;
signal \N__21245\ : std_logic;
signal \N__21242\ : std_logic;
signal \N__21239\ : std_logic;
signal \N__21234\ : std_logic;
signal \N__21233\ : std_logic;
signal \N__21232\ : std_logic;
signal \N__21231\ : std_logic;
signal \N__21230\ : std_logic;
signal \N__21229\ : std_logic;
signal \N__21228\ : std_logic;
signal \N__21227\ : std_logic;
signal \N__21224\ : std_logic;
signal \N__21223\ : std_logic;
signal \N__21222\ : std_logic;
signal \N__21221\ : std_logic;
signal \N__21220\ : std_logic;
signal \N__21219\ : std_logic;
signal \N__21218\ : std_logic;
signal \N__21217\ : std_logic;
signal \N__21216\ : std_logic;
signal \N__21215\ : std_logic;
signal \N__21214\ : std_logic;
signal \N__21213\ : std_logic;
signal \N__21212\ : std_logic;
signal \N__21211\ : std_logic;
signal \N__21210\ : std_logic;
signal \N__21209\ : std_logic;
signal \N__21208\ : std_logic;
signal \N__21207\ : std_logic;
signal \N__21206\ : std_logic;
signal \N__21205\ : std_logic;
signal \N__21204\ : std_logic;
signal \N__21203\ : std_logic;
signal \N__21202\ : std_logic;
signal \N__21201\ : std_logic;
signal \N__21192\ : std_logic;
signal \N__21187\ : std_logic;
signal \N__21184\ : std_logic;
signal \N__21181\ : std_logic;
signal \N__21178\ : std_logic;
signal \N__21173\ : std_logic;
signal \N__21170\ : std_logic;
signal \N__21169\ : std_logic;
signal \N__21168\ : std_logic;
signal \N__21167\ : std_logic;
signal \N__21164\ : std_logic;
signal \N__21155\ : std_logic;
signal \N__21146\ : std_logic;
signal \N__21145\ : std_logic;
signal \N__21140\ : std_logic;
signal \N__21131\ : std_logic;
signal \N__21130\ : std_logic;
signal \N__21123\ : std_logic;
signal \N__21120\ : std_logic;
signal \N__21115\ : std_logic;
signal \N__21112\ : std_logic;
signal \N__21109\ : std_logic;
signal \N__21106\ : std_logic;
signal \N__21101\ : std_logic;
signal \N__21100\ : std_logic;
signal \N__21099\ : std_logic;
signal \N__21098\ : std_logic;
signal \N__21097\ : std_logic;
signal \N__21094\ : std_logic;
signal \N__21091\ : std_logic;
signal \N__21090\ : std_logic;
signal \N__21089\ : std_logic;
signal \N__21088\ : std_logic;
signal \N__21087\ : std_logic;
signal \N__21086\ : std_logic;
signal \N__21085\ : std_logic;
signal \N__21084\ : std_logic;
signal \N__21083\ : std_logic;
signal \N__21080\ : std_logic;
signal \N__21073\ : std_logic;
signal \N__21070\ : std_logic;
signal \N__21065\ : std_logic;
signal \N__21064\ : std_logic;
signal \N__21063\ : std_logic;
signal \N__21062\ : std_logic;
signal \N__21061\ : std_logic;
signal \N__21060\ : std_logic;
signal \N__21057\ : std_logic;
signal \N__21056\ : std_logic;
signal \N__21055\ : std_logic;
signal \N__21054\ : std_logic;
signal \N__21053\ : std_logic;
signal \N__21044\ : std_logic;
signal \N__21041\ : std_logic;
signal \N__21038\ : std_logic;
signal \N__21035\ : std_logic;
signal \N__21032\ : std_logic;
signal \N__21021\ : std_logic;
signal \N__21010\ : std_logic;
signal \N__21005\ : std_logic;
signal \N__21002\ : std_logic;
signal \N__20993\ : std_logic;
signal \N__20984\ : std_logic;
signal \N__20979\ : std_logic;
signal \N__20970\ : std_logic;
signal \N__20943\ : std_logic;
signal \N__20940\ : std_logic;
signal \N__20937\ : std_logic;
signal \N__20934\ : std_logic;
signal \N__20931\ : std_logic;
signal \N__20930\ : std_logic;
signal \N__20927\ : std_logic;
signal \N__20926\ : std_logic;
signal \N__20923\ : std_logic;
signal \N__20920\ : std_logic;
signal \N__20917\ : std_logic;
signal \N__20914\ : std_logic;
signal \N__20911\ : std_logic;
signal \N__20908\ : std_logic;
signal \N__20905\ : std_logic;
signal \N__20902\ : std_logic;
signal \N__20899\ : std_logic;
signal \N__20894\ : std_logic;
signal \N__20889\ : std_logic;
signal \N__20886\ : std_logic;
signal \N__20885\ : std_logic;
signal \N__20882\ : std_logic;
signal \N__20879\ : std_logic;
signal \N__20876\ : std_logic;
signal \N__20875\ : std_logic;
signal \N__20872\ : std_logic;
signal \N__20869\ : std_logic;
signal \N__20866\ : std_logic;
signal \N__20863\ : std_logic;
signal \N__20856\ : std_logic;
signal \N__20853\ : std_logic;
signal \N__20850\ : std_logic;
signal \N__20847\ : std_logic;
signal \N__20844\ : std_logic;
signal \N__20841\ : std_logic;
signal \N__20838\ : std_logic;
signal \N__20835\ : std_logic;
signal \N__20832\ : std_logic;
signal \N__20829\ : std_logic;
signal \N__20828\ : std_logic;
signal \N__20825\ : std_logic;
signal \N__20822\ : std_logic;
signal \N__20817\ : std_logic;
signal \N__20816\ : std_logic;
signal \N__20815\ : std_logic;
signal \N__20812\ : std_logic;
signal \N__20809\ : std_logic;
signal \N__20806\ : std_logic;
signal \N__20801\ : std_logic;
signal \N__20798\ : std_logic;
signal \N__20793\ : std_logic;
signal \N__20790\ : std_logic;
signal \N__20787\ : std_logic;
signal \N__20784\ : std_logic;
signal \N__20781\ : std_logic;
signal \N__20778\ : std_logic;
signal \N__20777\ : std_logic;
signal \N__20772\ : std_logic;
signal \N__20771\ : std_logic;
signal \N__20770\ : std_logic;
signal \N__20767\ : std_logic;
signal \N__20762\ : std_logic;
signal \N__20757\ : std_logic;
signal \N__20754\ : std_logic;
signal \N__20753\ : std_logic;
signal \N__20752\ : std_logic;
signal \N__20749\ : std_logic;
signal \N__20746\ : std_logic;
signal \N__20743\ : std_logic;
signal \N__20736\ : std_logic;
signal \N__20733\ : std_logic;
signal \N__20732\ : std_logic;
signal \N__20731\ : std_logic;
signal \N__20728\ : std_logic;
signal \N__20725\ : std_logic;
signal \N__20722\ : std_logic;
signal \N__20715\ : std_logic;
signal \N__20712\ : std_logic;
signal \N__20709\ : std_logic;
signal \N__20706\ : std_logic;
signal \N__20703\ : std_logic;
signal \N__20700\ : std_logic;
signal \N__20697\ : std_logic;
signal \N__20694\ : std_logic;
signal \N__20691\ : std_logic;
signal \N__20688\ : std_logic;
signal \N__20685\ : std_logic;
signal \N__20682\ : std_logic;
signal \N__20679\ : std_logic;
signal \N__20676\ : std_logic;
signal \N__20675\ : std_logic;
signal \N__20672\ : std_logic;
signal \N__20669\ : std_logic;
signal \N__20664\ : std_logic;
signal \N__20663\ : std_logic;
signal \N__20660\ : std_logic;
signal \N__20659\ : std_logic;
signal \N__20656\ : std_logic;
signal \N__20653\ : std_logic;
signal \N__20650\ : std_logic;
signal \N__20647\ : std_logic;
signal \N__20644\ : std_logic;
signal \N__20641\ : std_logic;
signal \N__20638\ : std_logic;
signal \N__20635\ : std_logic;
signal \N__20632\ : std_logic;
signal \N__20625\ : std_logic;
signal \N__20622\ : std_logic;
signal \N__20619\ : std_logic;
signal \N__20616\ : std_logic;
signal \N__20615\ : std_logic;
signal \N__20614\ : std_logic;
signal \N__20611\ : std_logic;
signal \N__20608\ : std_logic;
signal \N__20605\ : std_logic;
signal \N__20602\ : std_logic;
signal \N__20599\ : std_logic;
signal \N__20592\ : std_logic;
signal \N__20591\ : std_logic;
signal \N__20588\ : std_logic;
signal \N__20587\ : std_logic;
signal \N__20586\ : std_logic;
signal \N__20583\ : std_logic;
signal \N__20580\ : std_logic;
signal \N__20577\ : std_logic;
signal \N__20574\ : std_logic;
signal \N__20571\ : std_logic;
signal \N__20562\ : std_logic;
signal \N__20559\ : std_logic;
signal \N__20556\ : std_logic;
signal \N__20553\ : std_logic;
signal \N__20550\ : std_logic;
signal \N__20547\ : std_logic;
signal \N__20544\ : std_logic;
signal \N__20541\ : std_logic;
signal \N__20540\ : std_logic;
signal \N__20539\ : std_logic;
signal \N__20536\ : std_logic;
signal \N__20533\ : std_logic;
signal \N__20532\ : std_logic;
signal \N__20531\ : std_logic;
signal \N__20528\ : std_logic;
signal \N__20525\ : std_logic;
signal \N__20522\ : std_logic;
signal \N__20515\ : std_logic;
signal \N__20512\ : std_logic;
signal \N__20507\ : std_logic;
signal \N__20502\ : std_logic;
signal \N__20501\ : std_logic;
signal \N__20498\ : std_logic;
signal \N__20495\ : std_logic;
signal \N__20492\ : std_logic;
signal \N__20487\ : std_logic;
signal \N__20484\ : std_logic;
signal \N__20481\ : std_logic;
signal \N__20478\ : std_logic;
signal \N__20475\ : std_logic;
signal \N__20472\ : std_logic;
signal \N__20469\ : std_logic;
signal \N__20466\ : std_logic;
signal \N__20463\ : std_logic;
signal \N__20460\ : std_logic;
signal \N__20459\ : std_logic;
signal \N__20458\ : std_logic;
signal \N__20455\ : std_logic;
signal \N__20450\ : std_logic;
signal \N__20449\ : std_logic;
signal \N__20444\ : std_logic;
signal \N__20441\ : std_logic;
signal \N__20440\ : std_logic;
signal \N__20435\ : std_logic;
signal \N__20432\ : std_logic;
signal \N__20429\ : std_logic;
signal \N__20426\ : std_logic;
signal \N__20421\ : std_logic;
signal \N__20420\ : std_logic;
signal \N__20419\ : std_logic;
signal \N__20418\ : std_logic;
signal \N__20415\ : std_logic;
signal \N__20414\ : std_logic;
signal \N__20409\ : std_logic;
signal \N__20408\ : std_logic;
signal \N__20407\ : std_logic;
signal \N__20406\ : std_logic;
signal \N__20403\ : std_logic;
signal \N__20400\ : std_logic;
signal \N__20399\ : std_logic;
signal \N__20398\ : std_logic;
signal \N__20397\ : std_logic;
signal \N__20396\ : std_logic;
signal \N__20395\ : std_logic;
signal \N__20392\ : std_logic;
signal \N__20391\ : std_logic;
signal \N__20388\ : std_logic;
signal \N__20381\ : std_logic;
signal \N__20376\ : std_logic;
signal \N__20371\ : std_logic;
signal \N__20368\ : std_logic;
signal \N__20363\ : std_logic;
signal \N__20362\ : std_logic;
signal \N__20359\ : std_logic;
signal \N__20356\ : std_logic;
signal \N__20351\ : std_logic;
signal \N__20350\ : std_logic;
signal \N__20349\ : std_logic;
signal \N__20348\ : std_logic;
signal \N__20347\ : std_logic;
signal \N__20346\ : std_logic;
signal \N__20345\ : std_logic;
signal \N__20344\ : std_logic;
signal \N__20343\ : std_logic;
signal \N__20342\ : std_logic;
signal \N__20337\ : std_logic;
signal \N__20334\ : std_logic;
signal \N__20331\ : std_logic;
signal \N__20328\ : std_logic;
signal \N__20321\ : std_logic;
signal \N__20316\ : std_logic;
signal \N__20311\ : std_logic;
signal \N__20302\ : std_logic;
signal \N__20299\ : std_logic;
signal \N__20294\ : std_logic;
signal \N__20287\ : std_logic;
signal \N__20274\ : std_logic;
signal \N__20273\ : std_logic;
signal \N__20272\ : std_logic;
signal \N__20269\ : std_logic;
signal \N__20266\ : std_logic;
signal \N__20263\ : std_logic;
signal \N__20258\ : std_logic;
signal \N__20257\ : std_logic;
signal \N__20256\ : std_logic;
signal \N__20255\ : std_logic;
signal \N__20250\ : std_logic;
signal \N__20247\ : std_logic;
signal \N__20244\ : std_logic;
signal \N__20243\ : std_logic;
signal \N__20242\ : std_logic;
signal \N__20241\ : std_logic;
signal \N__20240\ : std_logic;
signal \N__20237\ : std_logic;
signal \N__20236\ : std_logic;
signal \N__20235\ : std_logic;
signal \N__20232\ : std_logic;
signal \N__20229\ : std_logic;
signal \N__20226\ : std_logic;
signal \N__20223\ : std_logic;
signal \N__20222\ : std_logic;
signal \N__20219\ : std_logic;
signal \N__20218\ : std_logic;
signal \N__20217\ : std_logic;
signal \N__20214\ : std_logic;
signal \N__20211\ : std_logic;
signal \N__20208\ : std_logic;
signal \N__20203\ : std_logic;
signal \N__20200\ : std_logic;
signal \N__20193\ : std_logic;
signal \N__20190\ : std_logic;
signal \N__20187\ : std_logic;
signal \N__20182\ : std_logic;
signal \N__20177\ : std_logic;
signal \N__20160\ : std_logic;
signal \N__20159\ : std_logic;
signal \N__20158\ : std_logic;
signal \N__20157\ : std_logic;
signal \N__20152\ : std_logic;
signal \N__20151\ : std_logic;
signal \N__20150\ : std_logic;
signal \N__20147\ : std_logic;
signal \N__20144\ : std_logic;
signal \N__20143\ : std_logic;
signal \N__20140\ : std_logic;
signal \N__20137\ : std_logic;
signal \N__20134\ : std_logic;
signal \N__20133\ : std_logic;
signal \N__20132\ : std_logic;
signal \N__20129\ : std_logic;
signal \N__20128\ : std_logic;
signal \N__20127\ : std_logic;
signal \N__20124\ : std_logic;
signal \N__20121\ : std_logic;
signal \N__20120\ : std_logic;
signal \N__20119\ : std_logic;
signal \N__20116\ : std_logic;
signal \N__20115\ : std_logic;
signal \N__20110\ : std_logic;
signal \N__20105\ : std_logic;
signal \N__20104\ : std_logic;
signal \N__20103\ : std_logic;
signal \N__20100\ : std_logic;
signal \N__20097\ : std_logic;
signal \N__20094\ : std_logic;
signal \N__20091\ : std_logic;
signal \N__20088\ : std_logic;
signal \N__20083\ : std_logic;
signal \N__20080\ : std_logic;
signal \N__20077\ : std_logic;
signal \N__20072\ : std_logic;
signal \N__20067\ : std_logic;
signal \N__20060\ : std_logic;
signal \N__20043\ : std_logic;
signal \N__20040\ : std_logic;
signal \N__20039\ : std_logic;
signal \N__20036\ : std_logic;
signal \N__20033\ : std_logic;
signal \N__20032\ : std_logic;
signal \N__20029\ : std_logic;
signal \N__20026\ : std_logic;
signal \N__20023\ : std_logic;
signal \N__20018\ : std_logic;
signal \N__20015\ : std_logic;
signal \N__20014\ : std_logic;
signal \N__20011\ : std_logic;
signal \N__20008\ : std_logic;
signal \N__20005\ : std_logic;
signal \N__20002\ : std_logic;
signal \N__19995\ : std_logic;
signal \N__19992\ : std_logic;
signal \N__19989\ : std_logic;
signal \N__19988\ : std_logic;
signal \N__19985\ : std_logic;
signal \N__19984\ : std_logic;
signal \N__19981\ : std_logic;
signal \N__19978\ : std_logic;
signal \N__19973\ : std_logic;
signal \N__19968\ : std_logic;
signal \N__19965\ : std_logic;
signal \N__19962\ : std_logic;
signal \N__19959\ : std_logic;
signal \N__19958\ : std_logic;
signal \N__19955\ : std_logic;
signal \N__19954\ : std_logic;
signal \N__19951\ : std_logic;
signal \N__19948\ : std_logic;
signal \N__19945\ : std_logic;
signal \N__19942\ : std_logic;
signal \N__19937\ : std_logic;
signal \N__19932\ : std_logic;
signal \N__19931\ : std_logic;
signal \N__19928\ : std_logic;
signal \N__19927\ : std_logic;
signal \N__19924\ : std_logic;
signal \N__19921\ : std_logic;
signal \N__19918\ : std_logic;
signal \N__19915\ : std_logic;
signal \N__19912\ : std_logic;
signal \N__19909\ : std_logic;
signal \N__19902\ : std_logic;
signal \N__19899\ : std_logic;
signal \N__19896\ : std_logic;
signal \N__19893\ : std_logic;
signal \N__19890\ : std_logic;
signal \N__19887\ : std_logic;
signal \N__19884\ : std_logic;
signal \N__19881\ : std_logic;
signal \N__19878\ : std_logic;
signal \N__19877\ : std_logic;
signal \N__19874\ : std_logic;
signal \N__19871\ : std_logic;
signal \N__19866\ : std_logic;
signal \N__19863\ : std_logic;
signal \N__19862\ : std_logic;
signal \N__19861\ : std_logic;
signal \N__19860\ : std_logic;
signal \N__19859\ : std_logic;
signal \N__19858\ : std_logic;
signal \N__19855\ : std_logic;
signal \N__19852\ : std_logic;
signal \N__19849\ : std_logic;
signal \N__19844\ : std_logic;
signal \N__19841\ : std_logic;
signal \N__19830\ : std_logic;
signal \N__19827\ : std_logic;
signal \N__19826\ : std_logic;
signal \N__19823\ : std_logic;
signal \N__19822\ : std_logic;
signal \N__19821\ : std_logic;
signal \N__19820\ : std_logic;
signal \N__19819\ : std_logic;
signal \N__19818\ : std_logic;
signal \N__19817\ : std_logic;
signal \N__19816\ : std_logic;
signal \N__19815\ : std_logic;
signal \N__19812\ : std_logic;
signal \N__19809\ : std_logic;
signal \N__19806\ : std_logic;
signal \N__19801\ : std_logic;
signal \N__19798\ : std_logic;
signal \N__19795\ : std_logic;
signal \N__19790\ : std_logic;
signal \N__19785\ : std_logic;
signal \N__19770\ : std_logic;
signal \N__19769\ : std_logic;
signal \N__19768\ : std_logic;
signal \N__19767\ : std_logic;
signal \N__19766\ : std_logic;
signal \N__19765\ : std_logic;
signal \N__19762\ : std_logic;
signal \N__19759\ : std_logic;
signal \N__19756\ : std_logic;
signal \N__19753\ : std_logic;
signal \N__19750\ : std_logic;
signal \N__19747\ : std_logic;
signal \N__19746\ : std_logic;
signal \N__19745\ : std_logic;
signal \N__19742\ : std_logic;
signal \N__19739\ : std_logic;
signal \N__19730\ : std_logic;
signal \N__19727\ : std_logic;
signal \N__19724\ : std_logic;
signal \N__19715\ : std_logic;
signal \N__19714\ : std_logic;
signal \N__19713\ : std_logic;
signal \N__19710\ : std_logic;
signal \N__19707\ : std_logic;
signal \N__19706\ : std_logic;
signal \N__19705\ : std_logic;
signal \N__19702\ : std_logic;
signal \N__19701\ : std_logic;
signal \N__19698\ : std_logic;
signal \N__19695\ : std_logic;
signal \N__19692\ : std_logic;
signal \N__19691\ : std_logic;
signal \N__19690\ : std_logic;
signal \N__19689\ : std_logic;
signal \N__19688\ : std_logic;
signal \N__19687\ : std_logic;
signal \N__19686\ : std_logic;
signal \N__19683\ : std_logic;
signal \N__19680\ : std_logic;
signal \N__19675\ : std_logic;
signal \N__19672\ : std_logic;
signal \N__19669\ : std_logic;
signal \N__19666\ : std_logic;
signal \N__19655\ : std_logic;
signal \N__19650\ : std_logic;
signal \N__19643\ : std_logic;
signal \N__19632\ : std_logic;
signal \N__19631\ : std_logic;
signal \N__19630\ : std_logic;
signal \N__19627\ : std_logic;
signal \N__19626\ : std_logic;
signal \N__19625\ : std_logic;
signal \N__19624\ : std_logic;
signal \N__19623\ : std_logic;
signal \N__19622\ : std_logic;
signal \N__19621\ : std_logic;
signal \N__19620\ : std_logic;
signal \N__19615\ : std_logic;
signal \N__19610\ : std_logic;
signal \N__19607\ : std_logic;
signal \N__19604\ : std_logic;
signal \N__19603\ : std_logic;
signal \N__19598\ : std_logic;
signal \N__19597\ : std_logic;
signal \N__19594\ : std_logic;
signal \N__19593\ : std_logic;
signal \N__19592\ : std_logic;
signal \N__19591\ : std_logic;
signal \N__19588\ : std_logic;
signal \N__19587\ : std_logic;
signal \N__19582\ : std_logic;
signal \N__19577\ : std_logic;
signal \N__19574\ : std_logic;
signal \N__19571\ : std_logic;
signal \N__19568\ : std_logic;
signal \N__19565\ : std_logic;
signal \N__19558\ : std_logic;
signal \N__19555\ : std_logic;
signal \N__19554\ : std_logic;
signal \N__19553\ : std_logic;
signal \N__19552\ : std_logic;
signal \N__19551\ : std_logic;
signal \N__19548\ : std_logic;
signal \N__19541\ : std_logic;
signal \N__19540\ : std_logic;
signal \N__19539\ : std_logic;
signal \N__19538\ : std_logic;
signal \N__19533\ : std_logic;
signal \N__19526\ : std_logic;
signal \N__19521\ : std_logic;
signal \N__19516\ : std_logic;
signal \N__19513\ : std_logic;
signal \N__19510\ : std_logic;
signal \N__19507\ : std_logic;
signal \N__19502\ : std_logic;
signal \N__19497\ : std_logic;
signal \N__19492\ : std_logic;
signal \N__19479\ : std_logic;
signal \N__19476\ : std_logic;
signal \N__19475\ : std_logic;
signal \N__19472\ : std_logic;
signal \N__19471\ : std_logic;
signal \N__19468\ : std_logic;
signal \N__19467\ : std_logic;
signal \N__19464\ : std_logic;
signal \N__19461\ : std_logic;
signal \N__19458\ : std_logic;
signal \N__19455\ : std_logic;
signal \N__19452\ : std_logic;
signal \N__19449\ : std_logic;
signal \N__19444\ : std_logic;
signal \N__19441\ : std_logic;
signal \N__19436\ : std_logic;
signal \N__19431\ : std_logic;
signal \N__19428\ : std_logic;
signal \N__19425\ : std_logic;
signal \N__19424\ : std_logic;
signal \N__19421\ : std_logic;
signal \N__19418\ : std_logic;
signal \N__19415\ : std_logic;
signal \N__19410\ : std_logic;
signal \N__19407\ : std_logic;
signal \N__19406\ : std_logic;
signal \N__19405\ : std_logic;
signal \N__19402\ : std_logic;
signal \N__19399\ : std_logic;
signal \N__19396\ : std_logic;
signal \N__19393\ : std_logic;
signal \N__19390\ : std_logic;
signal \N__19387\ : std_logic;
signal \N__19384\ : std_logic;
signal \N__19381\ : std_logic;
signal \N__19374\ : std_logic;
signal \N__19373\ : std_logic;
signal \N__19370\ : std_logic;
signal \N__19367\ : std_logic;
signal \N__19364\ : std_logic;
signal \N__19361\ : std_logic;
signal \N__19360\ : std_logic;
signal \N__19357\ : std_logic;
signal \N__19354\ : std_logic;
signal \N__19351\ : std_logic;
signal \N__19348\ : std_logic;
signal \N__19345\ : std_logic;
signal \N__19338\ : std_logic;
signal \N__19337\ : std_logic;
signal \N__19336\ : std_logic;
signal \N__19333\ : std_logic;
signal \N__19330\ : std_logic;
signal \N__19325\ : std_logic;
signal \N__19322\ : std_logic;
signal \N__19319\ : std_logic;
signal \N__19318\ : std_logic;
signal \N__19315\ : std_logic;
signal \N__19312\ : std_logic;
signal \N__19309\ : std_logic;
signal \N__19306\ : std_logic;
signal \N__19303\ : std_logic;
signal \N__19296\ : std_logic;
signal \N__19295\ : std_logic;
signal \N__19292\ : std_logic;
signal \N__19289\ : std_logic;
signal \N__19286\ : std_logic;
signal \N__19283\ : std_logic;
signal \N__19280\ : std_logic;
signal \N__19277\ : std_logic;
signal \N__19274\ : std_logic;
signal \N__19271\ : std_logic;
signal \N__19266\ : std_logic;
signal \N__19263\ : std_logic;
signal \N__19262\ : std_logic;
signal \N__19259\ : std_logic;
signal \N__19256\ : std_logic;
signal \N__19253\ : std_logic;
signal \N__19250\ : std_logic;
signal \N__19247\ : std_logic;
signal \N__19244\ : std_logic;
signal \N__19239\ : std_logic;
signal \N__19236\ : std_logic;
signal \N__19235\ : std_logic;
signal \N__19232\ : std_logic;
signal \N__19231\ : std_logic;
signal \N__19230\ : std_logic;
signal \N__19227\ : std_logic;
signal \N__19224\ : std_logic;
signal \N__19221\ : std_logic;
signal \N__19218\ : std_logic;
signal \N__19209\ : std_logic;
signal \N__19206\ : std_logic;
signal \N__19203\ : std_logic;
signal \N__19200\ : std_logic;
signal \N__19197\ : std_logic;
signal \N__19194\ : std_logic;
signal \N__19191\ : std_logic;
signal \N__19188\ : std_logic;
signal \N__19187\ : std_logic;
signal \N__19184\ : std_logic;
signal \N__19181\ : std_logic;
signal \N__19180\ : std_logic;
signal \N__19177\ : std_logic;
signal \N__19174\ : std_logic;
signal \N__19171\ : std_logic;
signal \N__19170\ : std_logic;
signal \N__19167\ : std_logic;
signal \N__19164\ : std_logic;
signal \N__19159\ : std_logic;
signal \N__19156\ : std_logic;
signal \N__19153\ : std_logic;
signal \N__19150\ : std_logic;
signal \N__19143\ : std_logic;
signal \N__19140\ : std_logic;
signal \N__19137\ : std_logic;
signal \N__19134\ : std_logic;
signal \N__19131\ : std_logic;
signal \N__19128\ : std_logic;
signal \N__19125\ : std_logic;
signal \N__19122\ : std_logic;
signal \N__19119\ : std_logic;
signal \N__19116\ : std_logic;
signal \N__19113\ : std_logic;
signal \N__19110\ : std_logic;
signal \N__19107\ : std_logic;
signal \N__19104\ : std_logic;
signal \N__19101\ : std_logic;
signal \N__19098\ : std_logic;
signal \N__19095\ : std_logic;
signal \N__19092\ : std_logic;
signal \N__19089\ : std_logic;
signal \N__19088\ : std_logic;
signal \N__19085\ : std_logic;
signal \N__19082\ : std_logic;
signal \N__19081\ : std_logic;
signal \N__19078\ : std_logic;
signal \N__19075\ : std_logic;
signal \N__19072\ : std_logic;
signal \N__19069\ : std_logic;
signal \N__19066\ : std_logic;
signal \N__19059\ : std_logic;
signal \N__19056\ : std_logic;
signal \N__19053\ : std_logic;
signal \N__19050\ : std_logic;
signal \N__19047\ : std_logic;
signal \N__19044\ : std_logic;
signal \N__19043\ : std_logic;
signal \N__19040\ : std_logic;
signal \N__19037\ : std_logic;
signal \N__19036\ : std_logic;
signal \N__19033\ : std_logic;
signal \N__19030\ : std_logic;
signal \N__19027\ : std_logic;
signal \N__19024\ : std_logic;
signal \N__19021\ : std_logic;
signal \N__19014\ : std_logic;
signal \N__19011\ : std_logic;
signal \N__19010\ : std_logic;
signal \N__19007\ : std_logic;
signal \N__19004\ : std_logic;
signal \N__19001\ : std_logic;
signal \N__19000\ : std_logic;
signal \N__18997\ : std_logic;
signal \N__18994\ : std_logic;
signal \N__18991\ : std_logic;
signal \N__18984\ : std_logic;
signal \N__18981\ : std_logic;
signal \N__18978\ : std_logic;
signal \N__18975\ : std_logic;
signal \N__18972\ : std_logic;
signal \N__18969\ : std_logic;
signal \N__18966\ : std_logic;
signal \N__18965\ : std_logic;
signal \N__18962\ : std_logic;
signal \N__18959\ : std_logic;
signal \N__18956\ : std_logic;
signal \N__18955\ : std_logic;
signal \N__18952\ : std_logic;
signal \N__18949\ : std_logic;
signal \N__18946\ : std_logic;
signal \N__18939\ : std_logic;
signal \N__18936\ : std_logic;
signal \N__18933\ : std_logic;
signal \N__18932\ : std_logic;
signal \N__18929\ : std_logic;
signal \N__18926\ : std_logic;
signal \N__18921\ : std_logic;
signal \N__18920\ : std_logic;
signal \N__18917\ : std_logic;
signal \N__18914\ : std_logic;
signal \N__18911\ : std_logic;
signal \N__18908\ : std_logic;
signal \N__18903\ : std_logic;
signal \N__18902\ : std_logic;
signal \N__18901\ : std_logic;
signal \N__18900\ : std_logic;
signal \N__18899\ : std_logic;
signal \N__18898\ : std_logic;
signal \N__18897\ : std_logic;
signal \N__18894\ : std_logic;
signal \N__18893\ : std_logic;
signal \N__18890\ : std_logic;
signal \N__18887\ : std_logic;
signal \N__18886\ : std_logic;
signal \N__18885\ : std_logic;
signal \N__18882\ : std_logic;
signal \N__18881\ : std_logic;
signal \N__18878\ : std_logic;
signal \N__18877\ : std_logic;
signal \N__18876\ : std_logic;
signal \N__18871\ : std_logic;
signal \N__18868\ : std_logic;
signal \N__18865\ : std_logic;
signal \N__18860\ : std_logic;
signal \N__18855\ : std_logic;
signal \N__18854\ : std_logic;
signal \N__18851\ : std_logic;
signal \N__18848\ : std_logic;
signal \N__18845\ : std_logic;
signal \N__18842\ : std_logic;
signal \N__18839\ : std_logic;
signal \N__18836\ : std_logic;
signal \N__18827\ : std_logic;
signal \N__18826\ : std_logic;
signal \N__18823\ : std_logic;
signal \N__18820\ : std_logic;
signal \N__18817\ : std_logic;
signal \N__18814\ : std_logic;
signal \N__18805\ : std_logic;
signal \N__18802\ : std_logic;
signal \N__18789\ : std_logic;
signal \N__18788\ : std_logic;
signal \N__18787\ : std_logic;
signal \N__18784\ : std_logic;
signal \N__18783\ : std_logic;
signal \N__18782\ : std_logic;
signal \N__18781\ : std_logic;
signal \N__18780\ : std_logic;
signal \N__18777\ : std_logic;
signal \N__18776\ : std_logic;
signal \N__18775\ : std_logic;
signal \N__18772\ : std_logic;
signal \N__18769\ : std_logic;
signal \N__18764\ : std_logic;
signal \N__18763\ : std_logic;
signal \N__18760\ : std_logic;
signal \N__18759\ : std_logic;
signal \N__18756\ : std_logic;
signal \N__18751\ : std_logic;
signal \N__18748\ : std_logic;
signal \N__18745\ : std_logic;
signal \N__18742\ : std_logic;
signal \N__18741\ : std_logic;
signal \N__18740\ : std_logic;
signal \N__18739\ : std_logic;
signal \N__18736\ : std_logic;
signal \N__18735\ : std_logic;
signal \N__18732\ : std_logic;
signal \N__18727\ : std_logic;
signal \N__18724\ : std_logic;
signal \N__18721\ : std_logic;
signal \N__18716\ : std_logic;
signal \N__18713\ : std_logic;
signal \N__18710\ : std_logic;
signal \N__18707\ : std_logic;
signal \N__18704\ : std_logic;
signal \N__18701\ : std_logic;
signal \N__18698\ : std_logic;
signal \N__18695\ : std_logic;
signal \N__18692\ : std_logic;
signal \N__18687\ : std_logic;
signal \N__18666\ : std_logic;
signal \N__18663\ : std_logic;
signal \N__18660\ : std_logic;
signal \N__18657\ : std_logic;
signal \N__18654\ : std_logic;
signal \N__18653\ : std_logic;
signal \N__18650\ : std_logic;
signal \N__18647\ : std_logic;
signal \N__18644\ : std_logic;
signal \N__18641\ : std_logic;
signal \N__18640\ : std_logic;
signal \N__18637\ : std_logic;
signal \N__18634\ : std_logic;
signal \N__18631\ : std_logic;
signal \N__18628\ : std_logic;
signal \N__18623\ : std_logic;
signal \N__18618\ : std_logic;
signal \N__18615\ : std_logic;
signal \N__18612\ : std_logic;
signal \N__18611\ : std_logic;
signal \N__18608\ : std_logic;
signal \N__18605\ : std_logic;
signal \N__18600\ : std_logic;
signal \N__18597\ : std_logic;
signal \N__18594\ : std_logic;
signal \N__18591\ : std_logic;
signal \N__18590\ : std_logic;
signal \N__18589\ : std_logic;
signal \N__18586\ : std_logic;
signal \N__18581\ : std_logic;
signal \N__18576\ : std_logic;
signal \N__18573\ : std_logic;
signal \N__18572\ : std_logic;
signal \N__18571\ : std_logic;
signal \N__18568\ : std_logic;
signal \N__18563\ : std_logic;
signal \N__18558\ : std_logic;
signal \N__18555\ : std_logic;
signal \N__18552\ : std_logic;
signal \N__18551\ : std_logic;
signal \N__18550\ : std_logic;
signal \N__18547\ : std_logic;
signal \N__18544\ : std_logic;
signal \N__18541\ : std_logic;
signal \N__18534\ : std_logic;
signal \N__18533\ : std_logic;
signal \N__18532\ : std_logic;
signal \N__18529\ : std_logic;
signal \N__18526\ : std_logic;
signal \N__18523\ : std_logic;
signal \N__18516\ : std_logic;
signal \N__18513\ : std_logic;
signal \N__18512\ : std_logic;
signal \N__18509\ : std_logic;
signal \N__18506\ : std_logic;
signal \N__18501\ : std_logic;
signal \N__18498\ : std_logic;
signal \N__18495\ : std_logic;
signal \N__18494\ : std_logic;
signal \N__18493\ : std_logic;
signal \N__18490\ : std_logic;
signal \N__18487\ : std_logic;
signal \N__18484\ : std_logic;
signal \N__18479\ : std_logic;
signal \N__18476\ : std_logic;
signal \N__18473\ : std_logic;
signal \N__18468\ : std_logic;
signal \N__18465\ : std_logic;
signal \N__18462\ : std_logic;
signal \N__18459\ : std_logic;
signal \N__18458\ : std_logic;
signal \N__18457\ : std_logic;
signal \N__18454\ : std_logic;
signal \N__18449\ : std_logic;
signal \N__18444\ : std_logic;
signal \N__18441\ : std_logic;
signal \N__18438\ : std_logic;
signal \N__18435\ : std_logic;
signal \N__18432\ : std_logic;
signal \N__18429\ : std_logic;
signal \N__18428\ : std_logic;
signal \N__18427\ : std_logic;
signal \N__18424\ : std_logic;
signal \N__18419\ : std_logic;
signal \N__18414\ : std_logic;
signal \N__18413\ : std_logic;
signal \N__18410\ : std_logic;
signal \N__18407\ : std_logic;
signal \N__18406\ : std_logic;
signal \N__18403\ : std_logic;
signal \N__18400\ : std_logic;
signal \N__18397\ : std_logic;
signal \N__18392\ : std_logic;
signal \N__18387\ : std_logic;
signal \N__18384\ : std_logic;
signal \N__18381\ : std_logic;
signal \N__18378\ : std_logic;
signal \N__18375\ : std_logic;
signal \N__18372\ : std_logic;
signal \N__18369\ : std_logic;
signal \N__18366\ : std_logic;
signal \N__18363\ : std_logic;
signal \N__18360\ : std_logic;
signal \N__18357\ : std_logic;
signal \N__18354\ : std_logic;
signal \N__18351\ : std_logic;
signal \N__18348\ : std_logic;
signal \N__18345\ : std_logic;
signal \N__18342\ : std_logic;
signal \N__18339\ : std_logic;
signal \N__18336\ : std_logic;
signal \N__18333\ : std_logic;
signal \N__18330\ : std_logic;
signal \N__18327\ : std_logic;
signal \N__18324\ : std_logic;
signal \N__18321\ : std_logic;
signal \N__18318\ : std_logic;
signal \N__18317\ : std_logic;
signal \N__18314\ : std_logic;
signal \N__18311\ : std_logic;
signal \N__18308\ : std_logic;
signal \N__18305\ : std_logic;
signal \N__18300\ : std_logic;
signal \N__18297\ : std_logic;
signal \N__18294\ : std_logic;
signal \N__18291\ : std_logic;
signal \N__18290\ : std_logic;
signal \N__18289\ : std_logic;
signal \N__18286\ : std_logic;
signal \N__18283\ : std_logic;
signal \N__18280\ : std_logic;
signal \N__18277\ : std_logic;
signal \N__18274\ : std_logic;
signal \N__18273\ : std_logic;
signal \N__18270\ : std_logic;
signal \N__18267\ : std_logic;
signal \N__18264\ : std_logic;
signal \N__18261\ : std_logic;
signal \N__18258\ : std_logic;
signal \N__18253\ : std_logic;
signal \N__18250\ : std_logic;
signal \N__18243\ : std_logic;
signal \N__18240\ : std_logic;
signal \N__18237\ : std_logic;
signal \N__18234\ : std_logic;
signal \N__18231\ : std_logic;
signal \N__18228\ : std_logic;
signal \N__18225\ : std_logic;
signal \N__18222\ : std_logic;
signal \N__18219\ : std_logic;
signal \N__18216\ : std_logic;
signal \N__18213\ : std_logic;
signal \N__18210\ : std_logic;
signal \N__18207\ : std_logic;
signal \N__18204\ : std_logic;
signal \N__18201\ : std_logic;
signal \N__18198\ : std_logic;
signal \N__18195\ : std_logic;
signal \N__18192\ : std_logic;
signal \N__18189\ : std_logic;
signal \N__18186\ : std_logic;
signal \N__18183\ : std_logic;
signal \N__18180\ : std_logic;
signal \N__18177\ : std_logic;
signal \N__18174\ : std_logic;
signal \N__18171\ : std_logic;
signal \N__18168\ : std_logic;
signal \N__18165\ : std_logic;
signal \N__18162\ : std_logic;
signal \N__18159\ : std_logic;
signal \N__18156\ : std_logic;
signal \N__18153\ : std_logic;
signal \N__18152\ : std_logic;
signal \N__18149\ : std_logic;
signal \N__18146\ : std_logic;
signal \N__18145\ : std_logic;
signal \N__18140\ : std_logic;
signal \N__18137\ : std_logic;
signal \N__18132\ : std_logic;
signal \N__18131\ : std_logic;
signal \N__18128\ : std_logic;
signal \N__18125\ : std_logic;
signal \N__18120\ : std_logic;
signal \N__18117\ : std_logic;
signal \N__18114\ : std_logic;
signal \N__18111\ : std_logic;
signal \N__18108\ : std_logic;
signal \N__18105\ : std_logic;
signal \N__18102\ : std_logic;
signal \N__18099\ : std_logic;
signal \N__18096\ : std_logic;
signal \N__18093\ : std_logic;
signal \N__18090\ : std_logic;
signal \N__18087\ : std_logic;
signal \N__18084\ : std_logic;
signal \N__18081\ : std_logic;
signal \N__18078\ : std_logic;
signal \N__18075\ : std_logic;
signal \N__18072\ : std_logic;
signal \N__18069\ : std_logic;
signal \N__18066\ : std_logic;
signal \N__18063\ : std_logic;
signal \N__18060\ : std_logic;
signal \N__18057\ : std_logic;
signal \N__18054\ : std_logic;
signal \N__18051\ : std_logic;
signal \N__18048\ : std_logic;
signal \N__18047\ : std_logic;
signal \N__18044\ : std_logic;
signal \N__18041\ : std_logic;
signal \N__18040\ : std_logic;
signal \N__18039\ : std_logic;
signal \N__18036\ : std_logic;
signal \N__18033\ : std_logic;
signal \N__18030\ : std_logic;
signal \N__18027\ : std_logic;
signal \N__18018\ : std_logic;
signal \N__18015\ : std_logic;
signal \N__18012\ : std_logic;
signal \N__18009\ : std_logic;
signal \N__18006\ : std_logic;
signal \N__18003\ : std_logic;
signal \N__18000\ : std_logic;
signal \N__17997\ : std_logic;
signal \N__17994\ : std_logic;
signal \N__17991\ : std_logic;
signal \N__17988\ : std_logic;
signal \N__17985\ : std_logic;
signal \N__17982\ : std_logic;
signal \N__17979\ : std_logic;
signal \N__17976\ : std_logic;
signal \N__17973\ : std_logic;
signal \N__17970\ : std_logic;
signal \N__17967\ : std_logic;
signal \N__17964\ : std_logic;
signal \N__17961\ : std_logic;
signal \N__17958\ : std_logic;
signal \N__17955\ : std_logic;
signal \N__17952\ : std_logic;
signal \N__17949\ : std_logic;
signal \N__17946\ : std_logic;
signal \N__17943\ : std_logic;
signal \N__17940\ : std_logic;
signal \N__17937\ : std_logic;
signal \N__17934\ : std_logic;
signal \N__17933\ : std_logic;
signal \N__17930\ : std_logic;
signal \N__17929\ : std_logic;
signal \N__17926\ : std_logic;
signal \N__17923\ : std_logic;
signal \N__17920\ : std_logic;
signal \N__17917\ : std_logic;
signal \N__17916\ : std_logic;
signal \N__17913\ : std_logic;
signal \N__17910\ : std_logic;
signal \N__17907\ : std_logic;
signal \N__17904\ : std_logic;
signal \N__17895\ : std_logic;
signal \N__17892\ : std_logic;
signal \N__17889\ : std_logic;
signal \N__17886\ : std_logic;
signal \N__17883\ : std_logic;
signal \N__17880\ : std_logic;
signal \N__17879\ : std_logic;
signal \N__17876\ : std_logic;
signal \N__17873\ : std_logic;
signal \N__17872\ : std_logic;
signal \N__17871\ : std_logic;
signal \N__17866\ : std_logic;
signal \N__17865\ : std_logic;
signal \N__17864\ : std_logic;
signal \N__17861\ : std_logic;
signal \N__17858\ : std_logic;
signal \N__17855\ : std_logic;
signal \N__17850\ : std_logic;
signal \N__17847\ : std_logic;
signal \N__17838\ : std_logic;
signal \N__17835\ : std_logic;
signal \N__17834\ : std_logic;
signal \N__17831\ : std_logic;
signal \N__17828\ : std_logic;
signal \N__17825\ : std_logic;
signal \N__17822\ : std_logic;
signal \N__17817\ : std_logic;
signal \N__17814\ : std_logic;
signal \N__17813\ : std_logic;
signal \N__17812\ : std_logic;
signal \N__17811\ : std_logic;
signal \N__17808\ : std_logic;
signal \N__17807\ : std_logic;
signal \N__17806\ : std_logic;
signal \N__17805\ : std_logic;
signal \N__17804\ : std_logic;
signal \N__17803\ : std_logic;
signal \N__17802\ : std_logic;
signal \N__17799\ : std_logic;
signal \N__17796\ : std_logic;
signal \N__17793\ : std_logic;
signal \N__17790\ : std_logic;
signal \N__17787\ : std_logic;
signal \N__17782\ : std_logic;
signal \N__17777\ : std_logic;
signal \N__17772\ : std_logic;
signal \N__17757\ : std_logic;
signal \N__17754\ : std_logic;
signal \N__17751\ : std_logic;
signal \N__17748\ : std_logic;
signal \N__17745\ : std_logic;
signal \N__17744\ : std_logic;
signal \N__17741\ : std_logic;
signal \N__17738\ : std_logic;
signal \N__17737\ : std_logic;
signal \N__17736\ : std_logic;
signal \N__17735\ : std_logic;
signal \N__17730\ : std_logic;
signal \N__17723\ : std_logic;
signal \N__17718\ : std_logic;
signal \N__17717\ : std_logic;
signal \N__17716\ : std_logic;
signal \N__17715\ : std_logic;
signal \N__17714\ : std_logic;
signal \N__17713\ : std_logic;
signal \N__17712\ : std_logic;
signal \N__17711\ : std_logic;
signal \N__17710\ : std_logic;
signal \N__17709\ : std_logic;
signal \N__17706\ : std_logic;
signal \N__17705\ : std_logic;
signal \N__17704\ : std_logic;
signal \N__17703\ : std_logic;
signal \N__17700\ : std_logic;
signal \N__17697\ : std_logic;
signal \N__17694\ : std_logic;
signal \N__17691\ : std_logic;
signal \N__17688\ : std_logic;
signal \N__17687\ : std_logic;
signal \N__17684\ : std_logic;
signal \N__17681\ : std_logic;
signal \N__17676\ : std_logic;
signal \N__17673\ : std_logic;
signal \N__17670\ : std_logic;
signal \N__17669\ : std_logic;
signal \N__17668\ : std_logic;
signal \N__17667\ : std_logic;
signal \N__17666\ : std_logic;
signal \N__17663\ : std_logic;
signal \N__17660\ : std_logic;
signal \N__17657\ : std_logic;
signal \N__17650\ : std_logic;
signal \N__17647\ : std_logic;
signal \N__17644\ : std_logic;
signal \N__17637\ : std_logic;
signal \N__17632\ : std_logic;
signal \N__17629\ : std_logic;
signal \N__17626\ : std_logic;
signal \N__17623\ : std_logic;
signal \N__17618\ : std_logic;
signal \N__17613\ : std_logic;
signal \N__17604\ : std_logic;
signal \N__17601\ : std_logic;
signal \N__17586\ : std_logic;
signal \N__17583\ : std_logic;
signal \N__17580\ : std_logic;
signal \N__17579\ : std_logic;
signal \N__17576\ : std_logic;
signal \N__17573\ : std_logic;
signal \N__17568\ : std_logic;
signal \N__17565\ : std_logic;
signal \N__17564\ : std_logic;
signal \N__17563\ : std_logic;
signal \N__17562\ : std_logic;
signal \N__17561\ : std_logic;
signal \N__17560\ : std_logic;
signal \N__17559\ : std_logic;
signal \N__17556\ : std_logic;
signal \N__17553\ : std_logic;
signal \N__17552\ : std_logic;
signal \N__17549\ : std_logic;
signal \N__17548\ : std_logic;
signal \N__17545\ : std_logic;
signal \N__17542\ : std_logic;
signal \N__17541\ : std_logic;
signal \N__17540\ : std_logic;
signal \N__17539\ : std_logic;
signal \N__17536\ : std_logic;
signal \N__17535\ : std_logic;
signal \N__17534\ : std_logic;
signal \N__17531\ : std_logic;
signal \N__17530\ : std_logic;
signal \N__17529\ : std_logic;
signal \N__17524\ : std_logic;
signal \N__17521\ : std_logic;
signal \N__17520\ : std_logic;
signal \N__17517\ : std_logic;
signal \N__17510\ : std_logic;
signal \N__17509\ : std_logic;
signal \N__17508\ : std_logic;
signal \N__17507\ : std_logic;
signal \N__17504\ : std_logic;
signal \N__17501\ : std_logic;
signal \N__17496\ : std_logic;
signal \N__17493\ : std_logic;
signal \N__17488\ : std_logic;
signal \N__17487\ : std_logic;
signal \N__17486\ : std_logic;
signal \N__17485\ : std_logic;
signal \N__17484\ : std_logic;
signal \N__17483\ : std_logic;
signal \N__17480\ : std_logic;
signal \N__17477\ : std_logic;
signal \N__17476\ : std_logic;
signal \N__17473\ : std_logic;
signal \N__17468\ : std_logic;
signal \N__17463\ : std_logic;
signal \N__17462\ : std_logic;
signal \N__17461\ : std_logic;
signal \N__17460\ : std_logic;
signal \N__17459\ : std_logic;
signal \N__17458\ : std_logic;
signal \N__17455\ : std_logic;
signal \N__17448\ : std_logic;
signal \N__17445\ : std_logic;
signal \N__17442\ : std_logic;
signal \N__17439\ : std_logic;
signal \N__17436\ : std_logic;
signal \N__17435\ : std_logic;
signal \N__17434\ : std_logic;
signal \N__17433\ : std_logic;
signal \N__17432\ : std_logic;
signal \N__17429\ : std_logic;
signal \N__17414\ : std_logic;
signal \N__17411\ : std_logic;
signal \N__17406\ : std_logic;
signal \N__17403\ : std_logic;
signal \N__17400\ : std_logic;
signal \N__17397\ : std_logic;
signal \N__17390\ : std_logic;
signal \N__17383\ : std_logic;
signal \N__17380\ : std_logic;
signal \N__17377\ : std_logic;
signal \N__17374\ : std_logic;
signal \N__17367\ : std_logic;
signal \N__17364\ : std_logic;
signal \N__17359\ : std_logic;
signal \N__17354\ : std_logic;
signal \N__17351\ : std_logic;
signal \N__17348\ : std_logic;
signal \N__17345\ : std_logic;
signal \N__17342\ : std_logic;
signal \N__17339\ : std_logic;
signal \N__17336\ : std_logic;
signal \N__17325\ : std_logic;
signal \N__17310\ : std_logic;
signal \N__17307\ : std_logic;
signal \N__17306\ : std_logic;
signal \N__17305\ : std_logic;
signal \N__17304\ : std_logic;
signal \N__17301\ : std_logic;
signal \N__17296\ : std_logic;
signal \N__17293\ : std_logic;
signal \N__17288\ : std_logic;
signal \N__17283\ : std_logic;
signal \N__17280\ : std_logic;
signal \N__17277\ : std_logic;
signal \N__17276\ : std_logic;
signal \N__17273\ : std_logic;
signal \N__17270\ : std_logic;
signal \N__17265\ : std_logic;
signal \N__17262\ : std_logic;
signal \N__17259\ : std_logic;
signal \N__17258\ : std_logic;
signal \N__17255\ : std_logic;
signal \N__17252\ : std_logic;
signal \N__17247\ : std_logic;
signal \N__17244\ : std_logic;
signal \N__17241\ : std_logic;
signal \N__17238\ : std_logic;
signal \N__17235\ : std_logic;
signal \N__17234\ : std_logic;
signal \N__17231\ : std_logic;
signal \N__17228\ : std_logic;
signal \N__17223\ : std_logic;
signal \N__17220\ : std_logic;
signal \N__17217\ : std_logic;
signal \N__17216\ : std_logic;
signal \N__17213\ : std_logic;
signal \N__17210\ : std_logic;
signal \N__17205\ : std_logic;
signal \N__17202\ : std_logic;
signal \N__17199\ : std_logic;
signal \N__17196\ : std_logic;
signal \N__17193\ : std_logic;
signal \N__17192\ : std_logic;
signal \N__17189\ : std_logic;
signal \N__17188\ : std_logic;
signal \N__17185\ : std_logic;
signal \N__17184\ : std_logic;
signal \N__17183\ : std_logic;
signal \N__17182\ : std_logic;
signal \N__17181\ : std_logic;
signal \N__17178\ : std_logic;
signal \N__17175\ : std_logic;
signal \N__17172\ : std_logic;
signal \N__17169\ : std_logic;
signal \N__17162\ : std_logic;
signal \N__17151\ : std_logic;
signal \N__17148\ : std_logic;
signal \N__17147\ : std_logic;
signal \N__17144\ : std_logic;
signal \N__17141\ : std_logic;
signal \N__17138\ : std_logic;
signal \N__17133\ : std_logic;
signal \N__17130\ : std_logic;
signal \N__17127\ : std_logic;
signal \N__17124\ : std_logic;
signal \N__17121\ : std_logic;
signal \N__17118\ : std_logic;
signal \N__17115\ : std_logic;
signal \N__17112\ : std_logic;
signal \N__17109\ : std_logic;
signal \N__17106\ : std_logic;
signal \N__17105\ : std_logic;
signal \N__17102\ : std_logic;
signal \N__17099\ : std_logic;
signal \N__17096\ : std_logic;
signal \N__17093\ : std_logic;
signal \N__17088\ : std_logic;
signal \N__17087\ : std_logic;
signal \N__17082\ : std_logic;
signal \N__17079\ : std_logic;
signal \N__17076\ : std_logic;
signal \N__17073\ : std_logic;
signal \N__17070\ : std_logic;
signal \N__17067\ : std_logic;
signal \N__17064\ : std_logic;
signal \N__17061\ : std_logic;
signal \N__17060\ : std_logic;
signal \N__17059\ : std_logic;
signal \N__17058\ : std_logic;
signal \N__17055\ : std_logic;
signal \N__17052\ : std_logic;
signal \N__17051\ : std_logic;
signal \N__17050\ : std_logic;
signal \N__17049\ : std_logic;
signal \N__17046\ : std_logic;
signal \N__17045\ : std_logic;
signal \N__17044\ : std_logic;
signal \N__17041\ : std_logic;
signal \N__17038\ : std_logic;
signal \N__17037\ : std_logic;
signal \N__17036\ : std_logic;
signal \N__17033\ : std_logic;
signal \N__17030\ : std_logic;
signal \N__17029\ : std_logic;
signal \N__17028\ : std_logic;
signal \N__17027\ : std_logic;
signal \N__17024\ : std_logic;
signal \N__17021\ : std_logic;
signal \N__17018\ : std_logic;
signal \N__17015\ : std_logic;
signal \N__17012\ : std_logic;
signal \N__17007\ : std_logic;
signal \N__17002\ : std_logic;
signal \N__16997\ : std_logic;
signal \N__16994\ : std_logic;
signal \N__16989\ : std_logic;
signal \N__16984\ : std_logic;
signal \N__16981\ : std_logic;
signal \N__16962\ : std_logic;
signal \N__16959\ : std_logic;
signal \N__16956\ : std_logic;
signal \N__16953\ : std_logic;
signal \N__16950\ : std_logic;
signal \N__16947\ : std_logic;
signal \N__16944\ : std_logic;
signal \N__16941\ : std_logic;
signal \N__16938\ : std_logic;
signal \N__16935\ : std_logic;
signal \N__16932\ : std_logic;
signal \N__16929\ : std_logic;
signal \N__16926\ : std_logic;
signal \N__16923\ : std_logic;
signal \N__16922\ : std_logic;
signal \N__16921\ : std_logic;
signal \N__16920\ : std_logic;
signal \N__16919\ : std_logic;
signal \N__16918\ : std_logic;
signal \N__16915\ : std_logic;
signal \N__16914\ : std_logic;
signal \N__16911\ : std_logic;
signal \N__16910\ : std_logic;
signal \N__16907\ : std_logic;
signal \N__16904\ : std_logic;
signal \N__16901\ : std_logic;
signal \N__16896\ : std_logic;
signal \N__16889\ : std_logic;
signal \N__16882\ : std_logic;
signal \N__16881\ : std_logic;
signal \N__16880\ : std_logic;
signal \N__16879\ : std_logic;
signal \N__16878\ : std_logic;
signal \N__16877\ : std_logic;
signal \N__16876\ : std_logic;
signal \N__16875\ : std_logic;
signal \N__16872\ : std_logic;
signal \N__16867\ : std_logic;
signal \N__16864\ : std_logic;
signal \N__16863\ : std_logic;
signal \N__16860\ : std_logic;
signal \N__16857\ : std_logic;
signal \N__16854\ : std_logic;
signal \N__16853\ : std_logic;
signal \N__16850\ : std_logic;
signal \N__16847\ : std_logic;
signal \N__16844\ : std_logic;
signal \N__16843\ : std_logic;
signal \N__16838\ : std_logic;
signal \N__16833\ : std_logic;
signal \N__16826\ : std_logic;
signal \N__16823\ : std_logic;
signal \N__16816\ : std_logic;
signal \N__16813\ : std_logic;
signal \N__16800\ : std_logic;
signal \N__16799\ : std_logic;
signal \N__16798\ : std_logic;
signal \N__16797\ : std_logic;
signal \N__16796\ : std_logic;
signal \N__16795\ : std_logic;
signal \N__16794\ : std_logic;
signal \N__16793\ : std_logic;
signal \N__16792\ : std_logic;
signal \N__16791\ : std_logic;
signal \N__16790\ : std_logic;
signal \N__16789\ : std_logic;
signal \N__16788\ : std_logic;
signal \N__16787\ : std_logic;
signal \N__16786\ : std_logic;
signal \N__16783\ : std_logic;
signal \N__16782\ : std_logic;
signal \N__16781\ : std_logic;
signal \N__16780\ : std_logic;
signal \N__16767\ : std_logic;
signal \N__16762\ : std_logic;
signal \N__16759\ : std_logic;
signal \N__16748\ : std_logic;
signal \N__16739\ : std_logic;
signal \N__16736\ : std_logic;
signal \N__16733\ : std_logic;
signal \N__16722\ : std_logic;
signal \N__16719\ : std_logic;
signal \N__16716\ : std_logic;
signal \N__16713\ : std_logic;
signal \N__16710\ : std_logic;
signal \N__16707\ : std_logic;
signal \N__16704\ : std_logic;
signal \N__16701\ : std_logic;
signal \N__16698\ : std_logic;
signal \N__16695\ : std_logic;
signal \N__16692\ : std_logic;
signal \N__16689\ : std_logic;
signal \N__16688\ : std_logic;
signal \N__16685\ : std_logic;
signal \N__16682\ : std_logic;
signal \N__16677\ : std_logic;
signal \N__16674\ : std_logic;
signal \N__16671\ : std_logic;
signal \N__16668\ : std_logic;
signal \N__16665\ : std_logic;
signal \N__16662\ : std_logic;
signal \N__16659\ : std_logic;
signal \N__16656\ : std_logic;
signal \N__16653\ : std_logic;
signal \N__16650\ : std_logic;
signal \N__16649\ : std_logic;
signal \N__16646\ : std_logic;
signal \N__16643\ : std_logic;
signal \N__16638\ : std_logic;
signal \N__16635\ : std_logic;
signal \N__16632\ : std_logic;
signal \N__16629\ : std_logic;
signal \N__16626\ : std_logic;
signal \N__16623\ : std_logic;
signal \N__16620\ : std_logic;
signal \N__16617\ : std_logic;
signal \N__16614\ : std_logic;
signal \N__16613\ : std_logic;
signal \N__16610\ : std_logic;
signal \N__16607\ : std_logic;
signal \N__16602\ : std_logic;
signal \N__16599\ : std_logic;
signal \N__16596\ : std_logic;
signal \N__16593\ : std_logic;
signal \N__16590\ : std_logic;
signal \N__16587\ : std_logic;
signal \N__16584\ : std_logic;
signal \N__16581\ : std_logic;
signal \N__16578\ : std_logic;
signal \N__16575\ : std_logic;
signal \N__16572\ : std_logic;
signal \N__16569\ : std_logic;
signal \N__16566\ : std_logic;
signal \N__16563\ : std_logic;
signal \N__16560\ : std_logic;
signal \N__16557\ : std_logic;
signal \N__16554\ : std_logic;
signal \N__16551\ : std_logic;
signal \N__16548\ : std_logic;
signal \N__16545\ : std_logic;
signal \N__16542\ : std_logic;
signal \N__16539\ : std_logic;
signal \N__16536\ : std_logic;
signal \N__16533\ : std_logic;
signal \N__16530\ : std_logic;
signal \N__16527\ : std_logic;
signal \N__16524\ : std_logic;
signal \N__16521\ : std_logic;
signal \N__16518\ : std_logic;
signal \N__16515\ : std_logic;
signal \N__16512\ : std_logic;
signal \N__16509\ : std_logic;
signal \N__16506\ : std_logic;
signal \N__16503\ : std_logic;
signal \N__16500\ : std_logic;
signal \N__16497\ : std_logic;
signal \N__16494\ : std_logic;
signal \N__16491\ : std_logic;
signal \N__16488\ : std_logic;
signal \N__16485\ : std_logic;
signal \N__16482\ : std_logic;
signal \N__16479\ : std_logic;
signal \N__16476\ : std_logic;
signal \N__16473\ : std_logic;
signal \N__16472\ : std_logic;
signal \N__16469\ : std_logic;
signal \N__16466\ : std_logic;
signal \N__16461\ : std_logic;
signal \N__16458\ : std_logic;
signal \N__16455\ : std_logic;
signal \N__16452\ : std_logic;
signal \N__16449\ : std_logic;
signal \N__16448\ : std_logic;
signal \N__16445\ : std_logic;
signal \N__16442\ : std_logic;
signal \N__16439\ : std_logic;
signal \N__16436\ : std_logic;
signal \N__16433\ : std_logic;
signal \N__16428\ : std_logic;
signal \N__16425\ : std_logic;
signal \N__16422\ : std_logic;
signal \N__16419\ : std_logic;
signal \N__16416\ : std_logic;
signal \N__16413\ : std_logic;
signal \N__16410\ : std_logic;
signal \N__16407\ : std_logic;
signal \N__16404\ : std_logic;
signal \N__16401\ : std_logic;
signal \N__16398\ : std_logic;
signal \N__16395\ : std_logic;
signal \N__16392\ : std_logic;
signal \N__16389\ : std_logic;
signal \N__16386\ : std_logic;
signal \N__16383\ : std_logic;
signal \N__16380\ : std_logic;
signal \N__16377\ : std_logic;
signal \N__16374\ : std_logic;
signal \N__16371\ : std_logic;
signal \N__16370\ : std_logic;
signal \N__16367\ : std_logic;
signal \N__16364\ : std_logic;
signal \N__16363\ : std_logic;
signal \N__16360\ : std_logic;
signal \N__16357\ : std_logic;
signal \N__16354\ : std_logic;
signal \N__16351\ : std_logic;
signal \N__16348\ : std_logic;
signal \N__16345\ : std_logic;
signal \N__16338\ : std_logic;
signal \N__16335\ : std_logic;
signal \N__16332\ : std_logic;
signal \N__16329\ : std_logic;
signal \N__16326\ : std_logic;
signal \N__16323\ : std_logic;
signal \N__16320\ : std_logic;
signal \N__16317\ : std_logic;
signal \N__16314\ : std_logic;
signal \N__16311\ : std_logic;
signal \N__16308\ : std_logic;
signal \N__16305\ : std_logic;
signal \N__16302\ : std_logic;
signal \N__16299\ : std_logic;
signal \N__16296\ : std_logic;
signal \N__16293\ : std_logic;
signal \N__16290\ : std_logic;
signal \N__16287\ : std_logic;
signal \N__16284\ : std_logic;
signal \N__16281\ : std_logic;
signal \N__16278\ : std_logic;
signal \N__16275\ : std_logic;
signal \N__16272\ : std_logic;
signal \N__16269\ : std_logic;
signal \N__16266\ : std_logic;
signal \N__16263\ : std_logic;
signal \N__16262\ : std_logic;
signal \N__16261\ : std_logic;
signal \N__16258\ : std_logic;
signal \N__16255\ : std_logic;
signal \N__16254\ : std_logic;
signal \N__16253\ : std_logic;
signal \N__16250\ : std_logic;
signal \N__16245\ : std_logic;
signal \N__16244\ : std_logic;
signal \N__16243\ : std_logic;
signal \N__16240\ : std_logic;
signal \N__16237\ : std_logic;
signal \N__16234\ : std_logic;
signal \N__16231\ : std_logic;
signal \N__16228\ : std_logic;
signal \N__16225\ : std_logic;
signal \N__16222\ : std_logic;
signal \N__16215\ : std_logic;
signal \N__16212\ : std_logic;
signal \N__16209\ : std_logic;
signal \N__16206\ : std_logic;
signal \N__16203\ : std_logic;
signal \N__16200\ : std_logic;
signal \N__16193\ : std_logic;
signal \N__16188\ : std_logic;
signal \N__16185\ : std_logic;
signal \N__16184\ : std_logic;
signal \N__16181\ : std_logic;
signal \N__16178\ : std_logic;
signal \N__16173\ : std_logic;
signal \N__16170\ : std_logic;
signal \N__16167\ : std_logic;
signal \N__16164\ : std_logic;
signal \N__16161\ : std_logic;
signal \N__16158\ : std_logic;
signal \N__16155\ : std_logic;
signal \N__16152\ : std_logic;
signal \N__16149\ : std_logic;
signal \N__16146\ : std_logic;
signal \N__16143\ : std_logic;
signal \N__16140\ : std_logic;
signal \N__16137\ : std_logic;
signal \N__16134\ : std_logic;
signal \N__16133\ : std_logic;
signal \N__16130\ : std_logic;
signal \N__16127\ : std_logic;
signal \N__16124\ : std_logic;
signal \N__16121\ : std_logic;
signal \N__16116\ : std_logic;
signal \N__16113\ : std_logic;
signal \N__16110\ : std_logic;
signal \N__16107\ : std_logic;
signal \N__16104\ : std_logic;
signal \N__16101\ : std_logic;
signal \N__16098\ : std_logic;
signal \N__16095\ : std_logic;
signal \N__16092\ : std_logic;
signal \N__16091\ : std_logic;
signal \N__16088\ : std_logic;
signal \N__16085\ : std_logic;
signal \N__16082\ : std_logic;
signal \N__16079\ : std_logic;
signal \N__16074\ : std_logic;
signal \N__16071\ : std_logic;
signal \N__16068\ : std_logic;
signal \N__16067\ : std_logic;
signal \N__16064\ : std_logic;
signal \N__16061\ : std_logic;
signal \N__16058\ : std_logic;
signal \N__16055\ : std_logic;
signal \N__16050\ : std_logic;
signal \N__16047\ : std_logic;
signal \N__16044\ : std_logic;
signal \N__16041\ : std_logic;
signal \N__16038\ : std_logic;
signal \N__16035\ : std_logic;
signal \N__16032\ : std_logic;
signal \N__16029\ : std_logic;
signal \N__16026\ : std_logic;
signal \N__16023\ : std_logic;
signal \N__16020\ : std_logic;
signal \N__16017\ : std_logic;
signal \N__16016\ : std_logic;
signal \N__16013\ : std_logic;
signal \N__16010\ : std_logic;
signal \N__16005\ : std_logic;
signal \N__16002\ : std_logic;
signal \N__15999\ : std_logic;
signal \N__15996\ : std_logic;
signal \N__15993\ : std_logic;
signal \N__15992\ : std_logic;
signal \N__15989\ : std_logic;
signal \N__15986\ : std_logic;
signal \N__15983\ : std_logic;
signal \N__15980\ : std_logic;
signal \N__15975\ : std_logic;
signal \N__15972\ : std_logic;
signal \N__15969\ : std_logic;
signal \N__15966\ : std_logic;
signal \N__15963\ : std_logic;
signal \N__15960\ : std_logic;
signal \N__15957\ : std_logic;
signal \N__15954\ : std_logic;
signal \N__15951\ : std_logic;
signal \N__15948\ : std_logic;
signal \N__15945\ : std_logic;
signal \N__15942\ : std_logic;
signal \N__15939\ : std_logic;
signal \N__15936\ : std_logic;
signal \N__15933\ : std_logic;
signal \N__15930\ : std_logic;
signal \N__15929\ : std_logic;
signal \N__15926\ : std_logic;
signal \N__15923\ : std_logic;
signal \N__15920\ : std_logic;
signal \N__15917\ : std_logic;
signal \N__15912\ : std_logic;
signal \N__15909\ : std_logic;
signal \N__15906\ : std_logic;
signal \N__15903\ : std_logic;
signal \N__15900\ : std_logic;
signal \N__15897\ : std_logic;
signal \N__15894\ : std_logic;
signal \N__15891\ : std_logic;
signal \N__15888\ : std_logic;
signal \N__15885\ : std_logic;
signal \N__15882\ : std_logic;
signal \N__15879\ : std_logic;
signal \N__15878\ : std_logic;
signal \N__15875\ : std_logic;
signal \N__15872\ : std_logic;
signal \N__15867\ : std_logic;
signal \N__15866\ : std_logic;
signal \N__15863\ : std_logic;
signal \N__15860\ : std_logic;
signal \N__15857\ : std_logic;
signal \N__15854\ : std_logic;
signal \N__15849\ : std_logic;
signal \N__15846\ : std_logic;
signal \N__15843\ : std_logic;
signal \N__15840\ : std_logic;
signal \N__15839\ : std_logic;
signal \N__15836\ : std_logic;
signal \N__15833\ : std_logic;
signal \N__15830\ : std_logic;
signal \N__15827\ : std_logic;
signal \N__15822\ : std_logic;
signal \N__15819\ : std_logic;
signal \N__15816\ : std_logic;
signal \N__15813\ : std_logic;
signal \N__15810\ : std_logic;
signal \N__15807\ : std_logic;
signal \N__15806\ : std_logic;
signal \N__15801\ : std_logic;
signal \N__15798\ : std_logic;
signal \N__15795\ : std_logic;
signal \N__15792\ : std_logic;
signal \N__15789\ : std_logic;
signal \N__15786\ : std_logic;
signal \N__15783\ : std_logic;
signal \N__15780\ : std_logic;
signal \N__15777\ : std_logic;
signal \N__15776\ : std_logic;
signal \N__15773\ : std_logic;
signal \N__15770\ : std_logic;
signal \N__15767\ : std_logic;
signal \N__15764\ : std_logic;
signal \N__15761\ : std_logic;
signal \N__15758\ : std_logic;
signal \N__15753\ : std_logic;
signal \N__15750\ : std_logic;
signal \N__15747\ : std_logic;
signal \N__15744\ : std_logic;
signal \N__15741\ : std_logic;
signal \N__15740\ : std_logic;
signal \N__15737\ : std_logic;
signal \N__15732\ : std_logic;
signal \N__15729\ : std_logic;
signal \N__15726\ : std_logic;
signal \N__15723\ : std_logic;
signal \N__15720\ : std_logic;
signal \N__15717\ : std_logic;
signal \N__15716\ : std_logic;
signal \N__15713\ : std_logic;
signal \N__15710\ : std_logic;
signal \N__15707\ : std_logic;
signal \N__15704\ : std_logic;
signal \N__15701\ : std_logic;
signal \N__15698\ : std_logic;
signal \N__15693\ : std_logic;
signal \N__15690\ : std_logic;
signal \N__15687\ : std_logic;
signal \N__15684\ : std_logic;
signal \N__15681\ : std_logic;
signal \N__15678\ : std_logic;
signal \N__15675\ : std_logic;
signal \N__15674\ : std_logic;
signal \N__15673\ : std_logic;
signal \N__15670\ : std_logic;
signal \N__15667\ : std_logic;
signal \N__15664\ : std_logic;
signal \N__15661\ : std_logic;
signal \N__15658\ : std_logic;
signal \N__15651\ : std_logic;
signal \N__15650\ : std_logic;
signal \N__15649\ : std_logic;
signal \N__15646\ : std_logic;
signal \N__15643\ : std_logic;
signal \N__15640\ : std_logic;
signal \N__15637\ : std_logic;
signal \N__15634\ : std_logic;
signal \N__15629\ : std_logic;
signal \N__15626\ : std_logic;
signal \N__15621\ : std_logic;
signal \N__15618\ : std_logic;
signal \N__15615\ : std_logic;
signal \N__15612\ : std_logic;
signal \N__15609\ : std_logic;
signal \N__15606\ : std_logic;
signal \N__15603\ : std_logic;
signal \N__15600\ : std_logic;
signal \N__15597\ : std_logic;
signal \N__15594\ : std_logic;
signal \N__15591\ : std_logic;
signal \N__15588\ : std_logic;
signal \N__15585\ : std_logic;
signal \N__15582\ : std_logic;
signal \N__15579\ : std_logic;
signal \N__15576\ : std_logic;
signal \N__15573\ : std_logic;
signal \N__15570\ : std_logic;
signal \N__15567\ : std_logic;
signal \N__15564\ : std_logic;
signal \N__15561\ : std_logic;
signal \N__15558\ : std_logic;
signal \N__15555\ : std_logic;
signal \N__15552\ : std_logic;
signal \N__15549\ : std_logic;
signal \N__15546\ : std_logic;
signal \N__15543\ : std_logic;
signal \N__15540\ : std_logic;
signal \N__15537\ : std_logic;
signal \N__15534\ : std_logic;
signal \N__15531\ : std_logic;
signal \N__15528\ : std_logic;
signal \N__15525\ : std_logic;
signal \N__15522\ : std_logic;
signal \N__15519\ : std_logic;
signal \N__15516\ : std_logic;
signal \N__15513\ : std_logic;
signal \N__15510\ : std_logic;
signal \N__15507\ : std_logic;
signal \N__15504\ : std_logic;
signal \N__15501\ : std_logic;
signal \N__15498\ : std_logic;
signal \N__15495\ : std_logic;
signal \N__15492\ : std_logic;
signal \N__15489\ : std_logic;
signal \N__15486\ : std_logic;
signal \N__15483\ : std_logic;
signal \N__15480\ : std_logic;
signal \N__15477\ : std_logic;
signal \N__15474\ : std_logic;
signal \N__15471\ : std_logic;
signal \N__15468\ : std_logic;
signal \N__15465\ : std_logic;
signal \N__15462\ : std_logic;
signal \N__15459\ : std_logic;
signal \N__15456\ : std_logic;
signal \N__15453\ : std_logic;
signal \N__15450\ : std_logic;
signal \N__15447\ : std_logic;
signal \N__15444\ : std_logic;
signal \N__15441\ : std_logic;
signal \N__15438\ : std_logic;
signal \N__15435\ : std_logic;
signal \N__15432\ : std_logic;
signal \N__15429\ : std_logic;
signal \N__15426\ : std_logic;
signal \N__15423\ : std_logic;
signal \N__15420\ : std_logic;
signal \N__15417\ : std_logic;
signal \N__15414\ : std_logic;
signal \N__15411\ : std_logic;
signal \N__15410\ : std_logic;
signal \N__15407\ : std_logic;
signal \N__15404\ : std_logic;
signal \N__15401\ : std_logic;
signal \N__15398\ : std_logic;
signal \N__15395\ : std_logic;
signal \N__15392\ : std_logic;
signal \N__15387\ : std_logic;
signal \N__15384\ : std_logic;
signal \N__15381\ : std_logic;
signal \N__15378\ : std_logic;
signal \N__15375\ : std_logic;
signal \N__15372\ : std_logic;
signal \N__15371\ : std_logic;
signal \N__15368\ : std_logic;
signal \N__15367\ : std_logic;
signal \N__15364\ : std_logic;
signal \N__15361\ : std_logic;
signal \N__15358\ : std_logic;
signal \N__15351\ : std_logic;
signal \N__15348\ : std_logic;
signal \N__15345\ : std_logic;
signal \N__15342\ : std_logic;
signal \N__15339\ : std_logic;
signal \N__15336\ : std_logic;
signal \N__15333\ : std_logic;
signal \N__15330\ : std_logic;
signal \N__15327\ : std_logic;
signal \N__15324\ : std_logic;
signal \N__15321\ : std_logic;
signal \N__15318\ : std_logic;
signal \N__15315\ : std_logic;
signal \N__15312\ : std_logic;
signal \N__15311\ : std_logic;
signal \N__15310\ : std_logic;
signal \N__15307\ : std_logic;
signal \N__15302\ : std_logic;
signal \N__15297\ : std_logic;
signal \N__15294\ : std_logic;
signal \N__15291\ : std_logic;
signal \N__15288\ : std_logic;
signal \N__15285\ : std_logic;
signal \N__15284\ : std_logic;
signal \N__15281\ : std_logic;
signal \N__15278\ : std_logic;
signal \N__15275\ : std_logic;
signal \N__15272\ : std_logic;
signal \N__15267\ : std_logic;
signal \N__15266\ : std_logic;
signal \N__15263\ : std_logic;
signal \N__15260\ : std_logic;
signal \N__15257\ : std_logic;
signal \N__15254\ : std_logic;
signal \N__15251\ : std_logic;
signal \N__15248\ : std_logic;
signal \N__15243\ : std_logic;
signal \N__15240\ : std_logic;
signal \N__15237\ : std_logic;
signal \N__15234\ : std_logic;
signal \N__15231\ : std_logic;
signal \N__15230\ : std_logic;
signal \N__15229\ : std_logic;
signal \N__15226\ : std_logic;
signal \N__15223\ : std_logic;
signal \N__15222\ : std_logic;
signal \N__15219\ : std_logic;
signal \N__15214\ : std_logic;
signal \N__15211\ : std_logic;
signal \N__15208\ : std_logic;
signal \N__15205\ : std_logic;
signal \N__15202\ : std_logic;
signal \N__15195\ : std_logic;
signal \N__15194\ : std_logic;
signal \N__15191\ : std_logic;
signal \N__15188\ : std_logic;
signal \N__15185\ : std_logic;
signal \N__15184\ : std_logic;
signal \N__15181\ : std_logic;
signal \N__15178\ : std_logic;
signal \N__15175\ : std_logic;
signal \N__15174\ : std_logic;
signal \N__15171\ : std_logic;
signal \N__15168\ : std_logic;
signal \N__15165\ : std_logic;
signal \N__15162\ : std_logic;
signal \N__15153\ : std_logic;
signal \N__15152\ : std_logic;
signal \N__15149\ : std_logic;
signal \N__15146\ : std_logic;
signal \N__15143\ : std_logic;
signal \N__15140\ : std_logic;
signal \N__15135\ : std_logic;
signal \N__15134\ : std_logic;
signal \N__15131\ : std_logic;
signal \N__15128\ : std_logic;
signal \N__15123\ : std_logic;
signal \N__15120\ : std_logic;
signal \N__15117\ : std_logic;
signal \N__15114\ : std_logic;
signal \N__15111\ : std_logic;
signal \N__15108\ : std_logic;
signal \N__15107\ : std_logic;
signal \N__15106\ : std_logic;
signal \N__15105\ : std_logic;
signal \N__15102\ : std_logic;
signal \N__15099\ : std_logic;
signal \N__15096\ : std_logic;
signal \N__15095\ : std_logic;
signal \N__15094\ : std_logic;
signal \N__15093\ : std_logic;
signal \N__15090\ : std_logic;
signal \N__15083\ : std_logic;
signal \N__15080\ : std_logic;
signal \N__15077\ : std_logic;
signal \N__15074\ : std_logic;
signal \N__15073\ : std_logic;
signal \N__15070\ : std_logic;
signal \N__15061\ : std_logic;
signal \N__15058\ : std_logic;
signal \N__15057\ : std_logic;
signal \N__15056\ : std_logic;
signal \N__15053\ : std_logic;
signal \N__15048\ : std_logic;
signal \N__15045\ : std_logic;
signal \N__15042\ : std_logic;
signal \N__15033\ : std_logic;
signal \N__15030\ : std_logic;
signal \N__15027\ : std_logic;
signal \N__15024\ : std_logic;
signal \N__15021\ : std_logic;
signal \N__15018\ : std_logic;
signal \N__15017\ : std_logic;
signal \N__15014\ : std_logic;
signal \N__15011\ : std_logic;
signal \N__15008\ : std_logic;
signal \N__15005\ : std_logic;
signal \N__15000\ : std_logic;
signal \N__14997\ : std_logic;
signal \N__14994\ : std_logic;
signal \N__14991\ : std_logic;
signal \N__14990\ : std_logic;
signal \N__14987\ : std_logic;
signal \N__14984\ : std_logic;
signal \N__14979\ : std_logic;
signal \N__14976\ : std_logic;
signal \N__14973\ : std_logic;
signal \N__14972\ : std_logic;
signal \N__14969\ : std_logic;
signal \N__14966\ : std_logic;
signal \N__14961\ : std_logic;
signal \N__14958\ : std_logic;
signal \N__14955\ : std_logic;
signal \N__14952\ : std_logic;
signal \N__14949\ : std_logic;
signal \N__14948\ : std_logic;
signal \N__14947\ : std_logic;
signal \N__14946\ : std_logic;
signal \N__14943\ : std_logic;
signal \N__14940\ : std_logic;
signal \N__14939\ : std_logic;
signal \N__14934\ : std_logic;
signal \N__14933\ : std_logic;
signal \N__14932\ : std_logic;
signal \N__14929\ : std_logic;
signal \N__14926\ : std_logic;
signal \N__14923\ : std_logic;
signal \N__14920\ : std_logic;
signal \N__14917\ : std_logic;
signal \N__14916\ : std_logic;
signal \N__14913\ : std_logic;
signal \N__14906\ : std_logic;
signal \N__14901\ : std_logic;
signal \N__14896\ : std_logic;
signal \N__14893\ : std_logic;
signal \N__14886\ : std_logic;
signal \N__14883\ : std_logic;
signal \N__14880\ : std_logic;
signal \N__14877\ : std_logic;
signal \N__14874\ : std_logic;
signal \N__14871\ : std_logic;
signal \N__14868\ : std_logic;
signal \N__14865\ : std_logic;
signal \N__14864\ : std_logic;
signal \N__14861\ : std_logic;
signal \N__14858\ : std_logic;
signal \N__14855\ : std_logic;
signal \N__14854\ : std_logic;
signal \N__14851\ : std_logic;
signal \N__14848\ : std_logic;
signal \N__14845\ : std_logic;
signal \N__14838\ : std_logic;
signal \N__14835\ : std_logic;
signal \N__14832\ : std_logic;
signal \N__14829\ : std_logic;
signal \N__14826\ : std_logic;
signal \N__14823\ : std_logic;
signal \N__14820\ : std_logic;
signal \N__14817\ : std_logic;
signal \N__14814\ : std_logic;
signal \N__14811\ : std_logic;
signal \N__14810\ : std_logic;
signal \N__14807\ : std_logic;
signal \N__14804\ : std_logic;
signal \N__14801\ : std_logic;
signal \N__14798\ : std_logic;
signal \N__14793\ : std_logic;
signal \N__14792\ : std_logic;
signal \N__14789\ : std_logic;
signal \N__14786\ : std_logic;
signal \N__14781\ : std_logic;
signal \N__14780\ : std_logic;
signal \N__14777\ : std_logic;
signal \N__14774\ : std_logic;
signal \N__14769\ : std_logic;
signal \N__14766\ : std_logic;
signal \N__14765\ : std_logic;
signal \N__14762\ : std_logic;
signal \N__14759\ : std_logic;
signal \N__14754\ : std_logic;
signal \N__14751\ : std_logic;
signal \N__14748\ : std_logic;
signal \N__14747\ : std_logic;
signal \N__14742\ : std_logic;
signal \N__14739\ : std_logic;
signal \N__14736\ : std_logic;
signal \N__14735\ : std_logic;
signal \N__14732\ : std_logic;
signal \N__14729\ : std_logic;
signal \N__14726\ : std_logic;
signal \N__14721\ : std_logic;
signal \N__14718\ : std_logic;
signal \N__14715\ : std_logic;
signal \N__14712\ : std_logic;
signal \N__14709\ : std_logic;
signal \N__14706\ : std_logic;
signal \N__14703\ : std_logic;
signal \N__14700\ : std_logic;
signal \N__14697\ : std_logic;
signal \N__14696\ : std_logic;
signal \N__14691\ : std_logic;
signal \N__14688\ : std_logic;
signal \N__14687\ : std_logic;
signal \N__14684\ : std_logic;
signal \N__14681\ : std_logic;
signal \N__14676\ : std_logic;
signal \N__14675\ : std_logic;
signal \N__14672\ : std_logic;
signal \N__14667\ : std_logic;
signal \N__14664\ : std_logic;
signal \N__14663\ : std_logic;
signal \N__14660\ : std_logic;
signal \N__14657\ : std_logic;
signal \N__14652\ : std_logic;
signal \N__14649\ : std_logic;
signal \N__14648\ : std_logic;
signal \N__14647\ : std_logic;
signal \N__14646\ : std_logic;
signal \N__14641\ : std_logic;
signal \N__14636\ : std_logic;
signal \N__14631\ : std_logic;
signal \N__14628\ : std_logic;
signal \N__14625\ : std_logic;
signal \N__14624\ : std_logic;
signal \N__14621\ : std_logic;
signal \N__14618\ : std_logic;
signal \N__14615\ : std_logic;
signal \N__14612\ : std_logic;
signal \N__14607\ : std_logic;
signal \N__14606\ : std_logic;
signal \N__14603\ : std_logic;
signal \N__14602\ : std_logic;
signal \N__14599\ : std_logic;
signal \N__14598\ : std_logic;
signal \N__14595\ : std_logic;
signal \N__14592\ : std_logic;
signal \N__14587\ : std_logic;
signal \N__14580\ : std_logic;
signal \N__14577\ : std_logic;
signal \N__14574\ : std_logic;
signal \N__14571\ : std_logic;
signal \N__14568\ : std_logic;
signal \N__14565\ : std_logic;
signal \N__14564\ : std_logic;
signal \N__14561\ : std_logic;
signal \N__14558\ : std_logic;
signal \N__14553\ : std_logic;
signal \N__14550\ : std_logic;
signal \N__14547\ : std_logic;
signal \N__14546\ : std_logic;
signal \N__14543\ : std_logic;
signal \N__14540\ : std_logic;
signal \N__14535\ : std_logic;
signal \N__14532\ : std_logic;
signal \N__14531\ : std_logic;
signal \N__14528\ : std_logic;
signal \N__14525\ : std_logic;
signal \N__14522\ : std_logic;
signal \N__14517\ : std_logic;
signal \N__14514\ : std_logic;
signal \N__14511\ : std_logic;
signal \N__14510\ : std_logic;
signal \N__14507\ : std_logic;
signal \N__14504\ : std_logic;
signal \N__14501\ : std_logic;
signal \N__14496\ : std_logic;
signal \N__14493\ : std_logic;
signal \N__14490\ : std_logic;
signal \N__14487\ : std_logic;
signal \N__14486\ : std_logic;
signal \N__14483\ : std_logic;
signal \N__14480\ : std_logic;
signal \N__14477\ : std_logic;
signal \N__14472\ : std_logic;
signal \N__14469\ : std_logic;
signal \N__14468\ : std_logic;
signal \N__14465\ : std_logic;
signal \N__14462\ : std_logic;
signal \N__14457\ : std_logic;
signal \N__14454\ : std_logic;
signal \N__14453\ : std_logic;
signal \N__14450\ : std_logic;
signal \N__14447\ : std_logic;
signal \N__14442\ : std_logic;
signal \N__14439\ : std_logic;
signal \N__14438\ : std_logic;
signal \N__14435\ : std_logic;
signal \N__14432\ : std_logic;
signal \N__14427\ : std_logic;
signal \N__14424\ : std_logic;
signal \N__14423\ : std_logic;
signal \N__14420\ : std_logic;
signal \N__14417\ : std_logic;
signal \N__14412\ : std_logic;
signal \N__14409\ : std_logic;
signal \N__14408\ : std_logic;
signal \N__14405\ : std_logic;
signal \N__14402\ : std_logic;
signal \N__14397\ : std_logic;
signal \N__14394\ : std_logic;
signal \N__14393\ : std_logic;
signal \N__14390\ : std_logic;
signal \N__14387\ : std_logic;
signal \N__14384\ : std_logic;
signal \N__14379\ : std_logic;
signal \N__14376\ : std_logic;
signal \N__14375\ : std_logic;
signal \N__14372\ : std_logic;
signal \N__14369\ : std_logic;
signal \N__14364\ : std_logic;
signal \N__14361\ : std_logic;
signal \N__14360\ : std_logic;
signal \N__14357\ : std_logic;
signal \N__14354\ : std_logic;
signal \N__14349\ : std_logic;
signal \N__14346\ : std_logic;
signal \N__14345\ : std_logic;
signal \N__14342\ : std_logic;
signal \N__14339\ : std_logic;
signal \N__14334\ : std_logic;
signal \N__14331\ : std_logic;
signal \N__14328\ : std_logic;
signal \N__14327\ : std_logic;
signal \N__14326\ : std_logic;
signal \N__14325\ : std_logic;
signal \N__14324\ : std_logic;
signal \N__14321\ : std_logic;
signal \N__14318\ : std_logic;
signal \N__14311\ : std_logic;
signal \N__14308\ : std_logic;
signal \N__14301\ : std_logic;
signal \N__14298\ : std_logic;
signal \N__14297\ : std_logic;
signal \N__14292\ : std_logic;
signal \N__14291\ : std_logic;
signal \N__14290\ : std_logic;
signal \N__14289\ : std_logic;
signal \N__14286\ : std_logic;
signal \N__14283\ : std_logic;
signal \N__14280\ : std_logic;
signal \N__14279\ : std_logic;
signal \N__14276\ : std_logic;
signal \N__14273\ : std_logic;
signal \N__14268\ : std_logic;
signal \N__14265\ : std_logic;
signal \N__14256\ : std_logic;
signal \N__14253\ : std_logic;
signal \N__14250\ : std_logic;
signal \N__14249\ : std_logic;
signal \N__14248\ : std_logic;
signal \N__14247\ : std_logic;
signal \N__14244\ : std_logic;
signal \N__14241\ : std_logic;
signal \N__14240\ : std_logic;
signal \N__14237\ : std_logic;
signal \N__14234\ : std_logic;
signal \N__14233\ : std_logic;
signal \N__14228\ : std_logic;
signal \N__14227\ : std_logic;
signal \N__14224\ : std_logic;
signal \N__14219\ : std_logic;
signal \N__14218\ : std_logic;
signal \N__14217\ : std_logic;
signal \N__14214\ : std_logic;
signal \N__14211\ : std_logic;
signal \N__14208\ : std_logic;
signal \N__14205\ : std_logic;
signal \N__14202\ : std_logic;
signal \N__14197\ : std_logic;
signal \N__14184\ : std_logic;
signal \N__14183\ : std_logic;
signal \N__14180\ : std_logic;
signal \N__14177\ : std_logic;
signal \N__14176\ : std_logic;
signal \N__14173\ : std_logic;
signal \N__14170\ : std_logic;
signal \N__14167\ : std_logic;
signal \N__14164\ : std_logic;
signal \N__14159\ : std_logic;
signal \N__14156\ : std_logic;
signal \N__14153\ : std_logic;
signal \N__14148\ : std_logic;
signal \N__14145\ : std_logic;
signal \N__14144\ : std_logic;
signal \N__14143\ : std_logic;
signal \N__14142\ : std_logic;
signal \N__14139\ : std_logic;
signal \N__14136\ : std_logic;
signal \N__14133\ : std_logic;
signal \N__14130\ : std_logic;
signal \N__14125\ : std_logic;
signal \N__14118\ : std_logic;
signal \N__14117\ : std_logic;
signal \N__14116\ : std_logic;
signal \N__14115\ : std_logic;
signal \N__14114\ : std_logic;
signal \N__14111\ : std_logic;
signal \N__14108\ : std_logic;
signal \N__14103\ : std_logic;
signal \N__14100\ : std_logic;
signal \N__14091\ : std_logic;
signal \N__14088\ : std_logic;
signal \N__14085\ : std_logic;
signal \N__14082\ : std_logic;
signal \N__14081\ : std_logic;
signal \N__14080\ : std_logic;
signal \N__14079\ : std_logic;
signal \N__14076\ : std_logic;
signal \N__14073\ : std_logic;
signal \N__14070\ : std_logic;
signal \N__14067\ : std_logic;
signal \N__14058\ : std_logic;
signal \N__14057\ : std_logic;
signal \N__14056\ : std_logic;
signal \N__14053\ : std_logic;
signal \N__14050\ : std_logic;
signal \N__14047\ : std_logic;
signal \N__14044\ : std_logic;
signal \N__14041\ : std_logic;
signal \N__14034\ : std_logic;
signal \N__14033\ : std_logic;
signal \N__14030\ : std_logic;
signal \N__14027\ : std_logic;
signal \N__14022\ : std_logic;
signal \N__14019\ : std_logic;
signal \N__14016\ : std_logic;
signal \N__14013\ : std_logic;
signal \N__14012\ : std_logic;
signal \N__14009\ : std_logic;
signal \N__14006\ : std_logic;
signal \N__14001\ : std_logic;
signal \N__13998\ : std_logic;
signal \N__13995\ : std_logic;
signal \N__13992\ : std_logic;
signal \N__13989\ : std_logic;
signal \N__13986\ : std_logic;
signal \N__13983\ : std_logic;
signal \N__13980\ : std_logic;
signal \N__13977\ : std_logic;
signal \N__13974\ : std_logic;
signal \N__13973\ : std_logic;
signal \N__13972\ : std_logic;
signal \N__13969\ : std_logic;
signal \N__13966\ : std_logic;
signal \N__13963\ : std_logic;
signal \N__13960\ : std_logic;
signal \N__13957\ : std_logic;
signal \N__13950\ : std_logic;
signal \N__13949\ : std_logic;
signal \N__13948\ : std_logic;
signal \N__13947\ : std_logic;
signal \N__13944\ : std_logic;
signal \N__13941\ : std_logic;
signal \N__13936\ : std_logic;
signal \N__13929\ : std_logic;
signal \N__13926\ : std_logic;
signal \N__13925\ : std_logic;
signal \N__13924\ : std_logic;
signal \N__13921\ : std_logic;
signal \N__13920\ : std_logic;
signal \N__13917\ : std_logic;
signal \N__13914\ : std_logic;
signal \N__13909\ : std_logic;
signal \N__13902\ : std_logic;
signal \N__13899\ : std_logic;
signal \N__13898\ : std_logic;
signal \N__13895\ : std_logic;
signal \N__13892\ : std_logic;
signal \N__13889\ : std_logic;
signal \N__13886\ : std_logic;
signal \N__13883\ : std_logic;
signal \N__13880\ : std_logic;
signal \N__13875\ : std_logic;
signal \N__13872\ : std_logic;
signal \N__13869\ : std_logic;
signal \N__13866\ : std_logic;
signal \N__13863\ : std_logic;
signal \N__13860\ : std_logic;
signal \N__13857\ : std_logic;
signal \N__13854\ : std_logic;
signal \N__13851\ : std_logic;
signal \N__13848\ : std_logic;
signal \N__13845\ : std_logic;
signal \N__13842\ : std_logic;
signal \N__13841\ : std_logic;
signal \N__13838\ : std_logic;
signal \N__13835\ : std_logic;
signal \N__13830\ : std_logic;
signal \N__13827\ : std_logic;
signal \N__13824\ : std_logic;
signal \N__13821\ : std_logic;
signal \N__13820\ : std_logic;
signal \N__13817\ : std_logic;
signal \N__13814\ : std_logic;
signal \N__13809\ : std_logic;
signal \N__13806\ : std_logic;
signal \N__13803\ : std_logic;
signal \N__13800\ : std_logic;
signal \N__13797\ : std_logic;
signal \N__13794\ : std_logic;
signal \N__13793\ : std_logic;
signal \N__13790\ : std_logic;
signal \N__13787\ : std_logic;
signal \N__13782\ : std_logic;
signal \N__13779\ : std_logic;
signal \N__13776\ : std_logic;
signal \N__13773\ : std_logic;
signal \N__13770\ : std_logic;
signal \N__13769\ : std_logic;
signal \N__13766\ : std_logic;
signal \N__13763\ : std_logic;
signal \N__13760\ : std_logic;
signal \N__13757\ : std_logic;
signal \N__13752\ : std_logic;
signal \N__13749\ : std_logic;
signal \N__13748\ : std_logic;
signal \N__13745\ : std_logic;
signal \N__13742\ : std_logic;
signal \N__13739\ : std_logic;
signal \N__13736\ : std_logic;
signal \N__13731\ : std_logic;
signal \N__13728\ : std_logic;
signal \N__13725\ : std_logic;
signal \N__13722\ : std_logic;
signal \N__13719\ : std_logic;
signal \N__13716\ : std_logic;
signal \N__13713\ : std_logic;
signal \N__13710\ : std_logic;
signal \N__13709\ : std_logic;
signal \N__13706\ : std_logic;
signal \N__13703\ : std_logic;
signal \N__13698\ : std_logic;
signal \N__13695\ : std_logic;
signal \N__13692\ : std_logic;
signal \N__13689\ : std_logic;
signal \N__13686\ : std_logic;
signal \N__13683\ : std_logic;
signal \N__13680\ : std_logic;
signal \N__13677\ : std_logic;
signal \N__13674\ : std_logic;
signal \N__13673\ : std_logic;
signal \N__13670\ : std_logic;
signal \N__13667\ : std_logic;
signal \N__13662\ : std_logic;
signal \N__13659\ : std_logic;
signal \N__13656\ : std_logic;
signal \N__13653\ : std_logic;
signal \N__13650\ : std_logic;
signal \N__13647\ : std_logic;
signal \N__13644\ : std_logic;
signal \N__13641\ : std_logic;
signal \N__13638\ : std_logic;
signal \N__13635\ : std_logic;
signal \N__13632\ : std_logic;
signal \N__13629\ : std_logic;
signal \N__13626\ : std_logic;
signal \N__13623\ : std_logic;
signal \N__13620\ : std_logic;
signal \N__13617\ : std_logic;
signal \N__13616\ : std_logic;
signal \N__13613\ : std_logic;
signal \N__13610\ : std_logic;
signal \N__13607\ : std_logic;
signal \N__13604\ : std_logic;
signal \N__13601\ : std_logic;
signal \N__13598\ : std_logic;
signal \N__13593\ : std_logic;
signal \N__13590\ : std_logic;
signal \N__13589\ : std_logic;
signal \N__13586\ : std_logic;
signal \N__13583\ : std_logic;
signal \N__13580\ : std_logic;
signal \N__13577\ : std_logic;
signal \N__13572\ : std_logic;
signal \N__13569\ : std_logic;
signal \N__13566\ : std_logic;
signal \N__13563\ : std_logic;
signal \N__13560\ : std_logic;
signal \N__13559\ : std_logic;
signal \N__13556\ : std_logic;
signal \N__13553\ : std_logic;
signal \N__13550\ : std_logic;
signal \N__13547\ : std_logic;
signal \N__13542\ : std_logic;
signal \N__13539\ : std_logic;
signal \N__13536\ : std_logic;
signal \N__13533\ : std_logic;
signal \N__13530\ : std_logic;
signal \N__13527\ : std_logic;
signal \N__13526\ : std_logic;
signal \N__13523\ : std_logic;
signal \N__13520\ : std_logic;
signal \N__13517\ : std_logic;
signal \N__13514\ : std_logic;
signal \N__13509\ : std_logic;
signal \N__13506\ : std_logic;
signal \N__13505\ : std_logic;
signal \N__13504\ : std_logic;
signal \N__13503\ : std_logic;
signal \N__13500\ : std_logic;
signal \N__13497\ : std_logic;
signal \N__13494\ : std_logic;
signal \N__13491\ : std_logic;
signal \N__13486\ : std_logic;
signal \N__13483\ : std_logic;
signal \N__13480\ : std_logic;
signal \N__13473\ : std_logic;
signal \N__13472\ : std_logic;
signal \N__13469\ : std_logic;
signal \N__13466\ : std_logic;
signal \N__13461\ : std_logic;
signal \N__13460\ : std_logic;
signal \N__13459\ : std_logic;
signal \N__13456\ : std_logic;
signal \N__13453\ : std_logic;
signal \N__13450\ : std_logic;
signal \N__13443\ : std_logic;
signal \N__13440\ : std_logic;
signal \N__13437\ : std_logic;
signal \N__13434\ : std_logic;
signal \N__13431\ : std_logic;
signal \N__13430\ : std_logic;
signal \N__13427\ : std_logic;
signal \N__13424\ : std_logic;
signal \N__13421\ : std_logic;
signal \N__13416\ : std_logic;
signal \N__13413\ : std_logic;
signal \N__13410\ : std_logic;
signal \N__13407\ : std_logic;
signal \N__13404\ : std_logic;
signal \N__13401\ : std_logic;
signal \N__13398\ : std_logic;
signal \N__13395\ : std_logic;
signal \N__13392\ : std_logic;
signal \N__13389\ : std_logic;
signal \N__13386\ : std_logic;
signal \N__13385\ : std_logic;
signal \N__13384\ : std_logic;
signal \N__13383\ : std_logic;
signal \N__13382\ : std_logic;
signal \N__13381\ : std_logic;
signal \N__13380\ : std_logic;
signal \N__13379\ : std_logic;
signal \N__13368\ : std_logic;
signal \N__13361\ : std_logic;
signal \N__13360\ : std_logic;
signal \N__13355\ : std_logic;
signal \N__13352\ : std_logic;
signal \N__13347\ : std_logic;
signal \N__13346\ : std_logic;
signal \N__13343\ : std_logic;
signal \N__13340\ : std_logic;
signal \N__13337\ : std_logic;
signal \N__13334\ : std_logic;
signal \N__13329\ : std_logic;
signal \N__13326\ : std_logic;
signal \N__13325\ : std_logic;
signal \N__13322\ : std_logic;
signal \N__13319\ : std_logic;
signal \N__13316\ : std_logic;
signal \N__13313\ : std_logic;
signal \N__13308\ : std_logic;
signal \N__13305\ : std_logic;
signal \N__13302\ : std_logic;
signal \N__13301\ : std_logic;
signal \N__13298\ : std_logic;
signal \N__13295\ : std_logic;
signal \N__13290\ : std_logic;
signal \N__13289\ : std_logic;
signal \N__13286\ : std_logic;
signal \N__13283\ : std_logic;
signal \N__13280\ : std_logic;
signal \N__13277\ : std_logic;
signal \N__13274\ : std_logic;
signal \N__13271\ : std_logic;
signal \N__13266\ : std_logic;
signal \N__13265\ : std_logic;
signal \N__13264\ : std_logic;
signal \N__13263\ : std_logic;
signal \N__13254\ : std_logic;
signal \N__13253\ : std_logic;
signal \N__13250\ : std_logic;
signal \N__13247\ : std_logic;
signal \N__13246\ : std_logic;
signal \N__13241\ : std_logic;
signal \N__13238\ : std_logic;
signal \N__13237\ : std_logic;
signal \N__13236\ : std_logic;
signal \N__13235\ : std_logic;
signal \N__13234\ : std_logic;
signal \N__13231\ : std_logic;
signal \N__13228\ : std_logic;
signal \N__13225\ : std_logic;
signal \N__13218\ : std_logic;
signal \N__13209\ : std_logic;
signal \N__13208\ : std_logic;
signal \N__13205\ : std_logic;
signal \N__13202\ : std_logic;
signal \N__13199\ : std_logic;
signal \N__13196\ : std_logic;
signal \N__13193\ : std_logic;
signal \N__13190\ : std_logic;
signal \N__13185\ : std_logic;
signal \N__13182\ : std_logic;
signal \N__13179\ : std_logic;
signal \N__13176\ : std_logic;
signal \N__13173\ : std_logic;
signal \N__13172\ : std_logic;
signal \N__13169\ : std_logic;
signal \N__13168\ : std_logic;
signal \N__13165\ : std_logic;
signal \N__13162\ : std_logic;
signal \N__13161\ : std_logic;
signal \N__13158\ : std_logic;
signal \N__13157\ : std_logic;
signal \N__13156\ : std_logic;
signal \N__13155\ : std_logic;
signal \N__13154\ : std_logic;
signal \N__13149\ : std_logic;
signal \N__13140\ : std_logic;
signal \N__13137\ : std_logic;
signal \N__13134\ : std_logic;
signal \N__13131\ : std_logic;
signal \N__13128\ : std_logic;
signal \N__13119\ : std_logic;
signal \N__13118\ : std_logic;
signal \N__13117\ : std_logic;
signal \N__13116\ : std_logic;
signal \N__13113\ : std_logic;
signal \N__13112\ : std_logic;
signal \N__13111\ : std_logic;
signal \N__13110\ : std_logic;
signal \N__13107\ : std_logic;
signal \N__13106\ : std_logic;
signal \N__13103\ : std_logic;
signal \N__13100\ : std_logic;
signal \N__13099\ : std_logic;
signal \N__13094\ : std_logic;
signal \N__13093\ : std_logic;
signal \N__13092\ : std_logic;
signal \N__13091\ : std_logic;
signal \N__13090\ : std_logic;
signal \N__13089\ : std_logic;
signal \N__13084\ : std_logic;
signal \N__13081\ : std_logic;
signal \N__13078\ : std_logic;
signal \N__13075\ : std_logic;
signal \N__13072\ : std_logic;
signal \N__13069\ : std_logic;
signal \N__13066\ : std_logic;
signal \N__13063\ : std_logic;
signal \N__13062\ : std_logic;
signal \N__13061\ : std_logic;
signal \N__13054\ : std_logic;
signal \N__13051\ : std_logic;
signal \N__13044\ : std_logic;
signal \N__13039\ : std_logic;
signal \N__13032\ : std_logic;
signal \N__13027\ : std_logic;
signal \N__13020\ : std_logic;
signal \N__13011\ : std_logic;
signal \N__13008\ : std_logic;
signal \N__13005\ : std_logic;
signal \N__13004\ : std_logic;
signal \N__13001\ : std_logic;
signal \N__12998\ : std_logic;
signal \N__12993\ : std_logic;
signal \N__12992\ : std_logic;
signal \N__12987\ : std_logic;
signal \N__12986\ : std_logic;
signal \N__12985\ : std_logic;
signal \N__12982\ : std_logic;
signal \N__12981\ : std_logic;
signal \N__12978\ : std_logic;
signal \N__12977\ : std_logic;
signal \N__12976\ : std_logic;
signal \N__12975\ : std_logic;
signal \N__12974\ : std_logic;
signal \N__12973\ : std_logic;
signal \N__12970\ : std_logic;
signal \N__12967\ : std_logic;
signal \N__12964\ : std_logic;
signal \N__12961\ : std_logic;
signal \N__12950\ : std_logic;
signal \N__12939\ : std_logic;
signal \N__12936\ : std_logic;
signal \N__12935\ : std_logic;
signal \N__12930\ : std_logic;
signal \N__12929\ : std_logic;
signal \N__12926\ : std_logic;
signal \N__12925\ : std_logic;
signal \N__12924\ : std_logic;
signal \N__12923\ : std_logic;
signal \N__12922\ : std_logic;
signal \N__12921\ : std_logic;
signal \N__12920\ : std_logic;
signal \N__12919\ : std_logic;
signal \N__12918\ : std_logic;
signal \N__12915\ : std_logic;
signal \N__12912\ : std_logic;
signal \N__12907\ : std_logic;
signal \N__12904\ : std_logic;
signal \N__12899\ : std_logic;
signal \N__12892\ : std_logic;
signal \N__12879\ : std_logic;
signal \N__12878\ : std_logic;
signal \N__12877\ : std_logic;
signal \N__12876\ : std_logic;
signal \N__12871\ : std_logic;
signal \N__12866\ : std_logic;
signal \N__12863\ : std_logic;
signal \N__12862\ : std_logic;
signal \N__12861\ : std_logic;
signal \N__12860\ : std_logic;
signal \N__12859\ : std_logic;
signal \N__12858\ : std_logic;
signal \N__12857\ : std_logic;
signal \N__12856\ : std_logic;
signal \N__12855\ : std_logic;
signal \N__12850\ : std_logic;
signal \N__12847\ : std_logic;
signal \N__12842\ : std_logic;
signal \N__12831\ : std_logic;
signal \N__12822\ : std_logic;
signal \N__12819\ : std_logic;
signal \N__12816\ : std_logic;
signal \N__12813\ : std_logic;
signal \N__12810\ : std_logic;
signal \N__12807\ : std_logic;
signal \N__12804\ : std_logic;
signal \N__12801\ : std_logic;
signal \N__12798\ : std_logic;
signal \N__12795\ : std_logic;
signal \N__12792\ : std_logic;
signal \N__12789\ : std_logic;
signal \N__12788\ : std_logic;
signal \N__12787\ : std_logic;
signal \N__12786\ : std_logic;
signal \N__12783\ : std_logic;
signal \N__12780\ : std_logic;
signal \N__12779\ : std_logic;
signal \N__12778\ : std_logic;
signal \N__12777\ : std_logic;
signal \N__12774\ : std_logic;
signal \N__12771\ : std_logic;
signal \N__12766\ : std_logic;
signal \N__12763\ : std_logic;
signal \N__12760\ : std_logic;
signal \N__12757\ : std_logic;
signal \N__12752\ : std_logic;
signal \N__12745\ : std_logic;
signal \N__12742\ : std_logic;
signal \N__12741\ : std_logic;
signal \N__12740\ : std_logic;
signal \N__12739\ : std_logic;
signal \N__12736\ : std_logic;
signal \N__12731\ : std_logic;
signal \N__12728\ : std_logic;
signal \N__12725\ : std_logic;
signal \N__12722\ : std_logic;
signal \N__12711\ : std_logic;
signal \N__12708\ : std_logic;
signal \N__12705\ : std_logic;
signal \N__12704\ : std_logic;
signal \N__12699\ : std_logic;
signal \N__12698\ : std_logic;
signal \N__12695\ : std_logic;
signal \N__12692\ : std_logic;
signal \N__12689\ : std_logic;
signal \N__12686\ : std_logic;
signal \N__12681\ : std_logic;
signal \N__12680\ : std_logic;
signal \N__12677\ : std_logic;
signal \N__12674\ : std_logic;
signal \N__12671\ : std_logic;
signal \N__12666\ : std_logic;
signal \N__12663\ : std_logic;
signal \N__12660\ : std_logic;
signal \N__12659\ : std_logic;
signal \N__12658\ : std_logic;
signal \N__12655\ : std_logic;
signal \N__12652\ : std_logic;
signal \N__12649\ : std_logic;
signal \N__12644\ : std_logic;
signal \N__12639\ : std_logic;
signal \N__12638\ : std_logic;
signal \N__12637\ : std_logic;
signal \N__12634\ : std_logic;
signal \N__12633\ : std_logic;
signal \N__12632\ : std_logic;
signal \N__12631\ : std_logic;
signal \N__12630\ : std_logic;
signal \N__12629\ : std_logic;
signal \N__12628\ : std_logic;
signal \N__12627\ : std_logic;
signal \N__12626\ : std_logic;
signal \N__12623\ : std_logic;
signal \N__12620\ : std_logic;
signal \N__12603\ : std_logic;
signal \N__12600\ : std_logic;
signal \N__12599\ : std_logic;
signal \N__12596\ : std_logic;
signal \N__12595\ : std_logic;
signal \N__12592\ : std_logic;
signal \N__12587\ : std_logic;
signal \N__12584\ : std_logic;
signal \N__12581\ : std_logic;
signal \N__12578\ : std_logic;
signal \N__12571\ : std_logic;
signal \N__12564\ : std_logic;
signal \N__12563\ : std_logic;
signal \N__12560\ : std_logic;
signal \N__12557\ : std_logic;
signal \N__12554\ : std_logic;
signal \N__12551\ : std_logic;
signal \N__12546\ : std_logic;
signal \N__12545\ : std_logic;
signal \N__12544\ : std_logic;
signal \N__12543\ : std_logic;
signal \N__12540\ : std_logic;
signal \N__12537\ : std_logic;
signal \N__12534\ : std_logic;
signal \N__12531\ : std_logic;
signal \N__12530\ : std_logic;
signal \N__12529\ : std_logic;
signal \N__12528\ : std_logic;
signal \N__12519\ : std_logic;
signal \N__12516\ : std_logic;
signal \N__12513\ : std_logic;
signal \N__12510\ : std_logic;
signal \N__12509\ : std_logic;
signal \N__12500\ : std_logic;
signal \N__12497\ : std_logic;
signal \N__12496\ : std_logic;
signal \N__12495\ : std_logic;
signal \N__12490\ : std_logic;
signal \N__12487\ : std_logic;
signal \N__12484\ : std_logic;
signal \N__12477\ : std_logic;
signal \N__12474\ : std_logic;
signal \N__12471\ : std_logic;
signal \N__12470\ : std_logic;
signal \N__12467\ : std_logic;
signal \N__12464\ : std_logic;
signal \N__12459\ : std_logic;
signal \N__12458\ : std_logic;
signal \N__12457\ : std_logic;
signal \N__12456\ : std_logic;
signal \N__12455\ : std_logic;
signal \N__12452\ : std_logic;
signal \N__12449\ : std_logic;
signal \N__12446\ : std_logic;
signal \N__12443\ : std_logic;
signal \N__12440\ : std_logic;
signal \N__12439\ : std_logic;
signal \N__12438\ : std_logic;
signal \N__12435\ : std_logic;
signal \N__12432\ : std_logic;
signal \N__12427\ : std_logic;
signal \N__12424\ : std_logic;
signal \N__12421\ : std_logic;
signal \N__12418\ : std_logic;
signal \N__12417\ : std_logic;
signal \N__12414\ : std_logic;
signal \N__12411\ : std_logic;
signal \N__12402\ : std_logic;
signal \N__12399\ : std_logic;
signal \N__12398\ : std_logic;
signal \N__12397\ : std_logic;
signal \N__12394\ : std_logic;
signal \N__12391\ : std_logic;
signal \N__12386\ : std_logic;
signal \N__12383\ : std_logic;
signal \N__12380\ : std_logic;
signal \N__12369\ : std_logic;
signal \N__12366\ : std_logic;
signal \N__12365\ : std_logic;
signal \N__12364\ : std_logic;
signal \N__12361\ : std_logic;
signal \N__12356\ : std_logic;
signal \N__12351\ : std_logic;
signal \N__12348\ : std_logic;
signal \N__12345\ : std_logic;
signal \N__12342\ : std_logic;
signal \N__12341\ : std_logic;
signal \N__12340\ : std_logic;
signal \N__12339\ : std_logic;
signal \N__12334\ : std_logic;
signal \N__12329\ : std_logic;
signal \N__12326\ : std_logic;
signal \N__12321\ : std_logic;
signal \N__12318\ : std_logic;
signal \N__12315\ : std_logic;
signal \N__12312\ : std_logic;
signal \N__12311\ : std_logic;
signal \N__12310\ : std_logic;
signal \N__12309\ : std_logic;
signal \N__12306\ : std_logic;
signal \N__12303\ : std_logic;
signal \N__12300\ : std_logic;
signal \N__12297\ : std_logic;
signal \N__12292\ : std_logic;
signal \N__12285\ : std_logic;
signal \N__12284\ : std_logic;
signal \N__12281\ : std_logic;
signal \N__12278\ : std_logic;
signal \N__12277\ : std_logic;
signal \N__12276\ : std_logic;
signal \N__12275\ : std_logic;
signal \N__12274\ : std_logic;
signal \N__12273\ : std_logic;
signal \N__12272\ : std_logic;
signal \N__12267\ : std_logic;
signal \N__12264\ : std_logic;
signal \N__12261\ : std_logic;
signal \N__12258\ : std_logic;
signal \N__12255\ : std_logic;
signal \N__12250\ : std_logic;
signal \N__12237\ : std_logic;
signal \N__12234\ : std_logic;
signal \N__12231\ : std_logic;
signal \N__12228\ : std_logic;
signal \N__12225\ : std_logic;
signal \N__12222\ : std_logic;
signal \N__12219\ : std_logic;
signal \N__12216\ : std_logic;
signal \N__12215\ : std_logic;
signal \N__12214\ : std_logic;
signal \N__12213\ : std_logic;
signal \N__12210\ : std_logic;
signal \N__12209\ : std_logic;
signal \N__12208\ : std_logic;
signal \N__12207\ : std_logic;
signal \N__12206\ : std_logic;
signal \N__12203\ : std_logic;
signal \N__12202\ : std_logic;
signal \N__12197\ : std_logic;
signal \N__12192\ : std_logic;
signal \N__12189\ : std_logic;
signal \N__12186\ : std_logic;
signal \N__12183\ : std_logic;
signal \N__12180\ : std_logic;
signal \N__12177\ : std_logic;
signal \N__12174\ : std_logic;
signal \N__12171\ : std_logic;
signal \N__12156\ : std_logic;
signal \N__12153\ : std_logic;
signal \N__12150\ : std_logic;
signal \N__12147\ : std_logic;
signal \N__12144\ : std_logic;
signal \N__12141\ : std_logic;
signal \N__12138\ : std_logic;
signal \N__12135\ : std_logic;
signal \N__12132\ : std_logic;
signal \N__12131\ : std_logic;
signal \N__12128\ : std_logic;
signal \N__12125\ : std_logic;
signal \N__12120\ : std_logic;
signal \N__12119\ : std_logic;
signal \N__12118\ : std_logic;
signal \N__12117\ : std_logic;
signal \N__12116\ : std_logic;
signal \N__12115\ : std_logic;
signal \N__12114\ : std_logic;
signal \N__12113\ : std_logic;
signal \N__12096\ : std_logic;
signal \N__12093\ : std_logic;
signal \N__12090\ : std_logic;
signal \N__12087\ : std_logic;
signal \N__12086\ : std_logic;
signal \N__12085\ : std_logic;
signal \N__12084\ : std_logic;
signal \N__12081\ : std_logic;
signal \N__12078\ : std_logic;
signal \N__12075\ : std_logic;
signal \N__12072\ : std_logic;
signal \N__12063\ : std_logic;
signal \N__12060\ : std_logic;
signal \N__12057\ : std_logic;
signal \N__12054\ : std_logic;
signal \N__12053\ : std_logic;
signal \N__12048\ : std_logic;
signal \N__12045\ : std_logic;
signal \N__12042\ : std_logic;
signal \N__12041\ : std_logic;
signal \N__12040\ : std_logic;
signal \N__12033\ : std_logic;
signal \N__12032\ : std_logic;
signal \N__12029\ : std_logic;
signal \N__12026\ : std_logic;
signal \N__12021\ : std_logic;
signal \N__12020\ : std_logic;
signal \N__12017\ : std_logic;
signal \N__12014\ : std_logic;
signal \N__12009\ : std_logic;
signal \N__12006\ : std_logic;
signal \N__12005\ : std_logic;
signal \N__12000\ : std_logic;
signal \N__11997\ : std_logic;
signal \N__11994\ : std_logic;
signal \N__11993\ : std_logic;
signal \N__11990\ : std_logic;
signal \N__11987\ : std_logic;
signal \N__11982\ : std_logic;
signal \N__11979\ : std_logic;
signal \N__11976\ : std_logic;
signal \N__11973\ : std_logic;
signal \N__11970\ : std_logic;
signal \N__11967\ : std_logic;
signal \N__11966\ : std_logic;
signal \N__11965\ : std_logic;
signal \N__11964\ : std_logic;
signal \N__11963\ : std_logic;
signal \N__11962\ : std_logic;
signal \N__11961\ : std_logic;
signal \N__11960\ : std_logic;
signal \N__11959\ : std_logic;
signal \N__11940\ : std_logic;
signal \N__11937\ : std_logic;
signal \N__11934\ : std_logic;
signal \N__11931\ : std_logic;
signal \N__11928\ : std_logic;
signal \N__11925\ : std_logic;
signal \N__11922\ : std_logic;
signal \N__11919\ : std_logic;
signal \N__11916\ : std_logic;
signal \N__11913\ : std_logic;
signal \N__11912\ : std_logic;
signal \N__11909\ : std_logic;
signal \N__11906\ : std_logic;
signal \N__11903\ : std_logic;
signal \N__11900\ : std_logic;
signal \N__11895\ : std_logic;
signal \N__11892\ : std_logic;
signal \N__11889\ : std_logic;
signal \N__11886\ : std_logic;
signal \N__11883\ : std_logic;
signal \N__11880\ : std_logic;
signal \N__11877\ : std_logic;
signal \N__11874\ : std_logic;
signal \N__11871\ : std_logic;
signal \N__11868\ : std_logic;
signal \N__11865\ : std_logic;
signal \N__11862\ : std_logic;
signal \N__11859\ : std_logic;
signal \N__11858\ : std_logic;
signal \N__11857\ : std_logic;
signal \N__11854\ : std_logic;
signal \N__11851\ : std_logic;
signal \N__11850\ : std_logic;
signal \N__11847\ : std_logic;
signal \N__11844\ : std_logic;
signal \N__11839\ : std_logic;
signal \N__11832\ : std_logic;
signal \N__11829\ : std_logic;
signal \N__11826\ : std_logic;
signal \N__11825\ : std_logic;
signal \N__11820\ : std_logic;
signal \N__11817\ : std_logic;
signal \N__11814\ : std_logic;
signal \N__11811\ : std_logic;
signal \N__11810\ : std_logic;
signal \N__11805\ : std_logic;
signal \N__11802\ : std_logic;
signal \N__11799\ : std_logic;
signal \N__11796\ : std_logic;
signal \N__11795\ : std_logic;
signal \N__11790\ : std_logic;
signal \N__11787\ : std_logic;
signal \N__11784\ : std_logic;
signal \N__11781\ : std_logic;
signal \N__11780\ : std_logic;
signal \N__11775\ : std_logic;
signal \N__11772\ : std_logic;
signal \N__11769\ : std_logic;
signal \N__11766\ : std_logic;
signal \N__11765\ : std_logic;
signal \N__11760\ : std_logic;
signal \N__11757\ : std_logic;
signal \N__11754\ : std_logic;
signal \N__11751\ : std_logic;
signal \N__11750\ : std_logic;
signal \N__11747\ : std_logic;
signal \N__11744\ : std_logic;
signal \N__11739\ : std_logic;
signal \N__11736\ : std_logic;
signal \N__11735\ : std_logic;
signal \N__11732\ : std_logic;
signal \N__11729\ : std_logic;
signal \N__11724\ : std_logic;
signal \N__11721\ : std_logic;
signal \N__11718\ : std_logic;
signal \N__11715\ : std_logic;
signal \N__11712\ : std_logic;
signal \N__11709\ : std_logic;
signal \N__11706\ : std_logic;
signal \N__11703\ : std_logic;
signal \N__11700\ : std_logic;
signal \N__11697\ : std_logic;
signal \N__11694\ : std_logic;
signal \N__11691\ : std_logic;
signal \N__11690\ : std_logic;
signal \N__11687\ : std_logic;
signal \N__11684\ : std_logic;
signal \N__11683\ : std_logic;
signal \N__11682\ : std_logic;
signal \N__11679\ : std_logic;
signal \N__11674\ : std_logic;
signal \N__11671\ : std_logic;
signal \N__11668\ : std_logic;
signal \N__11665\ : std_logic;
signal \N__11658\ : std_logic;
signal \N__11655\ : std_logic;
signal \N__11654\ : std_logic;
signal \N__11651\ : std_logic;
signal \N__11648\ : std_logic;
signal \N__11643\ : std_logic;
signal \N__11640\ : std_logic;
signal \N__11637\ : std_logic;
signal \N__11636\ : std_logic;
signal \N__11633\ : std_logic;
signal \N__11630\ : std_logic;
signal \N__11627\ : std_logic;
signal \N__11622\ : std_logic;
signal \N__11619\ : std_logic;
signal \N__11616\ : std_logic;
signal \N__11613\ : std_logic;
signal \N__11612\ : std_logic;
signal \N__11607\ : std_logic;
signal \N__11604\ : std_logic;
signal \N__11603\ : std_logic;
signal \N__11600\ : std_logic;
signal \N__11597\ : std_logic;
signal \N__11592\ : std_logic;
signal \N__11589\ : std_logic;
signal \N__11586\ : std_logic;
signal \N__11585\ : std_logic;
signal \N__11584\ : std_logic;
signal \N__11583\ : std_logic;
signal \N__11582\ : std_logic;
signal \N__11581\ : std_logic;
signal \N__11580\ : std_logic;
signal \N__11577\ : std_logic;
signal \N__11574\ : std_logic;
signal \N__11571\ : std_logic;
signal \N__11570\ : std_logic;
signal \N__11567\ : std_logic;
signal \N__11564\ : std_logic;
signal \N__11561\ : std_logic;
signal \N__11558\ : std_logic;
signal \N__11555\ : std_logic;
signal \N__11554\ : std_logic;
signal \N__11553\ : std_logic;
signal \N__11548\ : std_logic;
signal \N__11545\ : std_logic;
signal \N__11544\ : std_logic;
signal \N__11533\ : std_logic;
signal \N__11530\ : std_logic;
signal \N__11527\ : std_logic;
signal \N__11524\ : std_logic;
signal \N__11519\ : std_logic;
signal \N__11514\ : std_logic;
signal \N__11505\ : std_logic;
signal \N__11502\ : std_logic;
signal \N__11499\ : std_logic;
signal \N__11498\ : std_logic;
signal \N__11495\ : std_logic;
signal \N__11492\ : std_logic;
signal \N__11487\ : std_logic;
signal \N__11484\ : std_logic;
signal \N__11481\ : std_logic;
signal \N__11478\ : std_logic;
signal \N__11477\ : std_logic;
signal \N__11474\ : std_logic;
signal \N__11471\ : std_logic;
signal \N__11468\ : std_logic;
signal \N__11463\ : std_logic;
signal \N__11460\ : std_logic;
signal \N__11459\ : std_logic;
signal \N__11456\ : std_logic;
signal \N__11453\ : std_logic;
signal \N__11448\ : std_logic;
signal \N__11445\ : std_logic;
signal \N__11442\ : std_logic;
signal \N__11439\ : std_logic;
signal \N__11436\ : std_logic;
signal \N__11435\ : std_logic;
signal \N__11434\ : std_logic;
signal \N__11431\ : std_logic;
signal \N__11430\ : std_logic;
signal \N__11427\ : std_logic;
signal \N__11424\ : std_logic;
signal \N__11421\ : std_logic;
signal \N__11418\ : std_logic;
signal \N__11415\ : std_logic;
signal \N__11412\ : std_logic;
signal \N__11403\ : std_logic;
signal \N__11402\ : std_logic;
signal \N__11399\ : std_logic;
signal \N__11396\ : std_logic;
signal \N__11395\ : std_logic;
signal \N__11394\ : std_logic;
signal \N__11391\ : std_logic;
signal \N__11388\ : std_logic;
signal \N__11385\ : std_logic;
signal \N__11382\ : std_logic;
signal \N__11375\ : std_logic;
signal \N__11370\ : std_logic;
signal \N__11367\ : std_logic;
signal \N__11366\ : std_logic;
signal \N__11361\ : std_logic;
signal \N__11358\ : std_logic;
signal \N__11355\ : std_logic;
signal \N__11352\ : std_logic;
signal \N__11351\ : std_logic;
signal \N__11346\ : std_logic;
signal \N__11343\ : std_logic;
signal \N__11340\ : std_logic;
signal \N__11337\ : std_logic;
signal \N__11336\ : std_logic;
signal \N__11331\ : std_logic;
signal \N__11328\ : std_logic;
signal \N__11325\ : std_logic;
signal \N__11322\ : std_logic;
signal \N__11321\ : std_logic;
signal \N__11316\ : std_logic;
signal \N__11313\ : std_logic;
signal \N__11310\ : std_logic;
signal \N__11307\ : std_logic;
signal \N__11306\ : std_logic;
signal \N__11301\ : std_logic;
signal \N__11298\ : std_logic;
signal \N__11295\ : std_logic;
signal \N__11292\ : std_logic;
signal \N__11291\ : std_logic;
signal \N__11286\ : std_logic;
signal \N__11283\ : std_logic;
signal \N__11280\ : std_logic;
signal \N__11279\ : std_logic;
signal \N__11276\ : std_logic;
signal \N__11273\ : std_logic;
signal \N__11268\ : std_logic;
signal \N__11265\ : std_logic;
signal \N__11262\ : std_logic;
signal \N__11259\ : std_logic;
signal \N__11256\ : std_logic;
signal \N__11253\ : std_logic;
signal \N__11252\ : std_logic;
signal \N__11249\ : std_logic;
signal \N__11246\ : std_logic;
signal \N__11245\ : std_logic;
signal \N__11244\ : std_logic;
signal \N__11243\ : std_logic;
signal \N__11242\ : std_logic;
signal \N__11241\ : std_logic;
signal \N__11236\ : std_logic;
signal \N__11233\ : std_logic;
signal \N__11230\ : std_logic;
signal \N__11227\ : std_logic;
signal \N__11224\ : std_logic;
signal \N__11221\ : std_logic;
signal \N__11220\ : std_logic;
signal \N__11217\ : std_logic;
signal \N__11214\ : std_logic;
signal \N__11213\ : std_logic;
signal \N__11212\ : std_logic;
signal \N__11211\ : std_logic;
signal \N__11204\ : std_logic;
signal \N__11201\ : std_logic;
signal \N__11198\ : std_logic;
signal \N__11195\ : std_logic;
signal \N__11192\ : std_logic;
signal \N__11189\ : std_logic;
signal \N__11184\ : std_logic;
signal \N__11177\ : std_logic;
signal \N__11166\ : std_logic;
signal \N__11165\ : std_logic;
signal \N__11162\ : std_logic;
signal \N__11161\ : std_logic;
signal \N__11158\ : std_logic;
signal \N__11155\ : std_logic;
signal \N__11152\ : std_logic;
signal \N__11151\ : std_logic;
signal \N__11150\ : std_logic;
signal \N__11147\ : std_logic;
signal \N__11144\ : std_logic;
signal \N__11137\ : std_logic;
signal \N__11130\ : std_logic;
signal \N__11127\ : std_logic;
signal \N__11124\ : std_logic;
signal \N__11123\ : std_logic;
signal \N__11120\ : std_logic;
signal \N__11117\ : std_logic;
signal \N__11112\ : std_logic;
signal \N__11111\ : std_logic;
signal \N__11108\ : std_logic;
signal \N__11105\ : std_logic;
signal \N__11102\ : std_logic;
signal \N__11099\ : std_logic;
signal \N__11094\ : std_logic;
signal \N__11093\ : std_logic;
signal \N__11090\ : std_logic;
signal \N__11087\ : std_logic;
signal \N__11086\ : std_logic;
signal \N__11085\ : std_logic;
signal \N__11084\ : std_logic;
signal \N__11083\ : std_logic;
signal \N__11082\ : std_logic;
signal \N__11081\ : std_logic;
signal \N__11076\ : std_logic;
signal \N__11073\ : std_logic;
signal \N__11070\ : std_logic;
signal \N__11067\ : std_logic;
signal \N__11064\ : std_logic;
signal \N__11061\ : std_logic;
signal \N__11058\ : std_logic;
signal \N__11051\ : std_logic;
signal \N__11048\ : std_logic;
signal \N__11047\ : std_logic;
signal \N__11046\ : std_logic;
signal \N__11045\ : std_logic;
signal \N__11040\ : std_logic;
signal \N__11037\ : std_logic;
signal \N__11034\ : std_logic;
signal \N__11031\ : std_logic;
signal \N__11028\ : std_logic;
signal \N__11023\ : std_logic;
signal \N__11018\ : std_logic;
signal \N__11007\ : std_logic;
signal \N__11004\ : std_logic;
signal \N__11003\ : std_logic;
signal \N__11000\ : std_logic;
signal \N__10997\ : std_logic;
signal \N__10994\ : std_logic;
signal \N__10991\ : std_logic;
signal \N__10986\ : std_logic;
signal \N__10985\ : std_logic;
signal \N__10982\ : std_logic;
signal \N__10979\ : std_logic;
signal \N__10978\ : std_logic;
signal \N__10977\ : std_logic;
signal \N__10976\ : std_logic;
signal \N__10975\ : std_logic;
signal \N__10974\ : std_logic;
signal \N__10969\ : std_logic;
signal \N__10966\ : std_logic;
signal \N__10963\ : std_logic;
signal \N__10960\ : std_logic;
signal \N__10957\ : std_logic;
signal \N__10954\ : std_logic;
signal \N__10953\ : std_logic;
signal \N__10946\ : std_logic;
signal \N__10945\ : std_logic;
signal \N__10944\ : std_logic;
signal \N__10943\ : std_logic;
signal \N__10936\ : std_logic;
signal \N__10933\ : std_logic;
signal \N__10930\ : std_logic;
signal \N__10927\ : std_logic;
signal \N__10922\ : std_logic;
signal \N__10917\ : std_logic;
signal \N__10908\ : std_logic;
signal \N__10905\ : std_logic;
signal \N__10904\ : std_logic;
signal \N__10901\ : std_logic;
signal \N__10898\ : std_logic;
signal \N__10893\ : std_logic;
signal \N__10890\ : std_logic;
signal \N__10889\ : std_logic;
signal \N__10886\ : std_logic;
signal \N__10883\ : std_logic;
signal \N__10878\ : std_logic;
signal \N__10875\ : std_logic;
signal \N__10872\ : std_logic;
signal \N__10869\ : std_logic;
signal \N__10866\ : std_logic;
signal \N__10863\ : std_logic;
signal \N__10860\ : std_logic;
signal \N__10857\ : std_logic;
signal \N__10856\ : std_logic;
signal \N__10853\ : std_logic;
signal \N__10850\ : std_logic;
signal \N__10845\ : std_logic;
signal \N__10842\ : std_logic;
signal \N__10839\ : std_logic;
signal \N__10836\ : std_logic;
signal \N__10833\ : std_logic;
signal \N__10830\ : std_logic;
signal \N__10827\ : std_logic;
signal \N__10824\ : std_logic;
signal \N__10823\ : std_logic;
signal \N__10820\ : std_logic;
signal \N__10817\ : std_logic;
signal \N__10814\ : std_logic;
signal \N__10809\ : std_logic;
signal \N__10808\ : std_logic;
signal \N__10807\ : std_logic;
signal \N__10800\ : std_logic;
signal \N__10797\ : std_logic;
signal \N__10794\ : std_logic;
signal \N__10793\ : std_logic;
signal \N__10788\ : std_logic;
signal \N__10785\ : std_logic;
signal \N__10782\ : std_logic;
signal \N__10779\ : std_logic;
signal \N__10776\ : std_logic;
signal \N__10773\ : std_logic;
signal \N__10772\ : std_logic;
signal \N__10769\ : std_logic;
signal \N__10766\ : std_logic;
signal \N__10763\ : std_logic;
signal \N__10760\ : std_logic;
signal \N__10755\ : std_logic;
signal \N__10752\ : std_logic;
signal \N__10749\ : std_logic;
signal \N__10746\ : std_logic;
signal \N__10743\ : std_logic;
signal \N__10740\ : std_logic;
signal \N__10737\ : std_logic;
signal \N__10734\ : std_logic;
signal \N__10731\ : std_logic;
signal \N__10728\ : std_logic;
signal \N__10725\ : std_logic;
signal \N__10722\ : std_logic;
signal \N__10719\ : std_logic;
signal \N__10716\ : std_logic;
signal \N__10713\ : std_logic;
signal \N__10710\ : std_logic;
signal \N__10707\ : std_logic;
signal \N__10704\ : std_logic;
signal \N__10701\ : std_logic;
signal \N__10700\ : std_logic;
signal \N__10697\ : std_logic;
signal \N__10694\ : std_logic;
signal \N__10693\ : std_logic;
signal \N__10686\ : std_logic;
signal \N__10683\ : std_logic;
signal \N__10680\ : std_logic;
signal \N__10677\ : std_logic;
signal \N__10674\ : std_logic;
signal \N__10671\ : std_logic;
signal \N__10668\ : std_logic;
signal \N__10665\ : std_logic;
signal \N__10662\ : std_logic;
signal \N__10661\ : std_logic;
signal \N__10656\ : std_logic;
signal \N__10653\ : std_logic;
signal \N__10650\ : std_logic;
signal \N__10647\ : std_logic;
signal \N__10646\ : std_logic;
signal \N__10641\ : std_logic;
signal \N__10638\ : std_logic;
signal \N__10635\ : std_logic;
signal \N__10632\ : std_logic;
signal \N__10631\ : std_logic;
signal \N__10626\ : std_logic;
signal \N__10623\ : std_logic;
signal \N__10620\ : std_logic;
signal \N__10617\ : std_logic;
signal \N__10616\ : std_logic;
signal \N__10611\ : std_logic;
signal \N__10608\ : std_logic;
signal \N__10605\ : std_logic;
signal \N__10602\ : std_logic;
signal \N__10601\ : std_logic;
signal \N__10596\ : std_logic;
signal \N__10593\ : std_logic;
signal \N__10590\ : std_logic;
signal \N__10587\ : std_logic;
signal \N__10586\ : std_logic;
signal \N__10581\ : std_logic;
signal \N__10578\ : std_logic;
signal \N__10575\ : std_logic;
signal \N__10574\ : std_logic;
signal \N__10571\ : std_logic;
signal \N__10568\ : std_logic;
signal \N__10563\ : std_logic;
signal \N__10560\ : std_logic;
signal \N__10557\ : std_logic;
signal \N__10554\ : std_logic;
signal \N__10551\ : std_logic;
signal \N__10548\ : std_logic;
signal \N__10545\ : std_logic;
signal \N__10542\ : std_logic;
signal \N__10539\ : std_logic;
signal \N__10536\ : std_logic;
signal \N__10533\ : std_logic;
signal \N__10530\ : std_logic;
signal \N__10527\ : std_logic;
signal \N__10524\ : std_logic;
signal \N__10521\ : std_logic;
signal \N__10518\ : std_logic;
signal \N__10515\ : std_logic;
signal \N__10512\ : std_logic;
signal \N__10511\ : std_logic;
signal \N__10508\ : std_logic;
signal \N__10505\ : std_logic;
signal \N__10504\ : std_logic;
signal \N__10503\ : std_logic;
signal \N__10500\ : std_logic;
signal \N__10497\ : std_logic;
signal \N__10494\ : std_logic;
signal \N__10491\ : std_logic;
signal \N__10482\ : std_logic;
signal \N__10481\ : std_logic;
signal \N__10478\ : std_logic;
signal \N__10475\ : std_logic;
signal \N__10474\ : std_logic;
signal \N__10473\ : std_logic;
signal \N__10470\ : std_logic;
signal \N__10467\ : std_logic;
signal \N__10464\ : std_logic;
signal \N__10461\ : std_logic;
signal \N__10458\ : std_logic;
signal \N__10449\ : std_logic;
signal \N__10446\ : std_logic;
signal \N__10443\ : std_logic;
signal \N__10440\ : std_logic;
signal \N__10439\ : std_logic;
signal \N__10438\ : std_logic;
signal \N__10435\ : std_logic;
signal \N__10432\ : std_logic;
signal \N__10431\ : std_logic;
signal \N__10428\ : std_logic;
signal \N__10425\ : std_logic;
signal \N__10420\ : std_logic;
signal \N__10413\ : std_logic;
signal \N__10410\ : std_logic;
signal \N__10407\ : std_logic;
signal \N__10404\ : std_logic;
signal \N__10401\ : std_logic;
signal \N__10398\ : std_logic;
signal \N__10395\ : std_logic;
signal \N__10392\ : std_logic;
signal \N__10389\ : std_logic;
signal \N__10386\ : std_logic;
signal \N__10383\ : std_logic;
signal \N__10380\ : std_logic;
signal \N__10377\ : std_logic;
signal \N__10374\ : std_logic;
signal \N__10371\ : std_logic;
signal \N__10368\ : std_logic;
signal \N__10365\ : std_logic;
signal \N__10362\ : std_logic;
signal \N__10359\ : std_logic;
signal \N__10356\ : std_logic;
signal \N__10353\ : std_logic;
signal \N__10350\ : std_logic;
signal \N__10347\ : std_logic;
signal \N__10344\ : std_logic;
signal \N__10341\ : std_logic;
signal \N__10338\ : std_logic;
signal \N__10335\ : std_logic;
signal \N__10332\ : std_logic;
signal \N__10329\ : std_logic;
signal \N__10326\ : std_logic;
signal \N__10323\ : std_logic;
signal \N__10320\ : std_logic;
signal \N__10317\ : std_logic;
signal \N__10314\ : std_logic;
signal \N__10311\ : std_logic;
signal \N__10308\ : std_logic;
signal \N__10305\ : std_logic;
signal \N__10302\ : std_logic;
signal \N__10299\ : std_logic;
signal \N__10296\ : std_logic;
signal \N__10293\ : std_logic;
signal \N__10290\ : std_logic;
signal \N__10287\ : std_logic;
signal \N__10284\ : std_logic;
signal \N__10281\ : std_logic;
signal \N__10278\ : std_logic;
signal \N__10277\ : std_logic;
signal \N__10274\ : std_logic;
signal \N__10271\ : std_logic;
signal \N__10266\ : std_logic;
signal \N__10265\ : std_logic;
signal \N__10260\ : std_logic;
signal \N__10257\ : std_logic;
signal \N__10254\ : std_logic;
signal \N__10253\ : std_logic;
signal \N__10248\ : std_logic;
signal \N__10245\ : std_logic;
signal \N__10242\ : std_logic;
signal \N__10239\ : std_logic;
signal \N__10236\ : std_logic;
signal \N__10235\ : std_logic;
signal \N__10232\ : std_logic;
signal \N__10229\ : std_logic;
signal \N__10226\ : std_logic;
signal \N__10221\ : std_logic;
signal \N__10218\ : std_logic;
signal \N__10215\ : std_logic;
signal \N__10212\ : std_logic;
signal \N__10209\ : std_logic;
signal \N__10206\ : std_logic;
signal \N__10203\ : std_logic;
signal \N__10202\ : std_logic;
signal \N__10199\ : std_logic;
signal \N__10196\ : std_logic;
signal \N__10191\ : std_logic;
signal \N__10188\ : std_logic;
signal \N__10185\ : std_logic;
signal \N__10182\ : std_logic;
signal \N__10179\ : std_logic;
signal \N__10176\ : std_logic;
signal \N__10173\ : std_logic;
signal \N__10170\ : std_logic;
signal \N__10167\ : std_logic;
signal \N__10164\ : std_logic;
signal \N__10161\ : std_logic;
signal \N__10158\ : std_logic;
signal \N__10155\ : std_logic;
signal \N__10152\ : std_logic;
signal \N__10149\ : std_logic;
signal \N__10146\ : std_logic;
signal \N__10143\ : std_logic;
signal \N__10140\ : std_logic;
signal \N__10137\ : std_logic;
signal \N__10134\ : std_logic;
signal \N__10131\ : std_logic;
signal \N__10128\ : std_logic;
signal \N__10125\ : std_logic;
signal \N__10122\ : std_logic;
signal \N__10119\ : std_logic;
signal \N__10118\ : std_logic;
signal \N__10115\ : std_logic;
signal \N__10112\ : std_logic;
signal \N__10109\ : std_logic;
signal \N__10104\ : std_logic;
signal \N__10101\ : std_logic;
signal \N__10098\ : std_logic;
signal \N__10095\ : std_logic;
signal \N__10092\ : std_logic;
signal \N__10089\ : std_logic;
signal \N__10086\ : std_logic;
signal \N__10083\ : std_logic;
signal \N__10080\ : std_logic;
signal \N__10077\ : std_logic;
signal \N__10074\ : std_logic;
signal \N__10071\ : std_logic;
signal \N__10068\ : std_logic;
signal \N__10065\ : std_logic;
signal \N__10062\ : std_logic;
signal \N__10059\ : std_logic;
signal \N__10056\ : std_logic;
signal \N__10053\ : std_logic;
signal \N__10050\ : std_logic;
signal \N__10047\ : std_logic;
signal \N__10044\ : std_logic;
signal \N__10041\ : std_logic;
signal \N__10038\ : std_logic;
signal \N__10035\ : std_logic;
signal \N__10032\ : std_logic;
signal \N__10031\ : std_logic;
signal \N__10028\ : std_logic;
signal \N__10025\ : std_logic;
signal \N__10020\ : std_logic;
signal \N__10017\ : std_logic;
signal \N__10016\ : std_logic;
signal \N__10013\ : std_logic;
signal \N__10010\ : std_logic;
signal \N__10007\ : std_logic;
signal \N__10002\ : std_logic;
signal \N__10001\ : std_logic;
signal \N__9998\ : std_logic;
signal \N__9997\ : std_logic;
signal \N__9994\ : std_logic;
signal \N__9989\ : std_logic;
signal \N__9984\ : std_logic;
signal \N__9983\ : std_logic;
signal \N__9982\ : std_logic;
signal \N__9981\ : std_logic;
signal \N__9978\ : std_logic;
signal \N__9971\ : std_logic;
signal \N__9966\ : std_logic;
signal \N__9965\ : std_logic;
signal \N__9962\ : std_logic;
signal \N__9961\ : std_logic;
signal \N__9960\ : std_logic;
signal \N__9957\ : std_logic;
signal \N__9954\ : std_logic;
signal \N__9949\ : std_logic;
signal \N__9942\ : std_logic;
signal \N__9939\ : std_logic;
signal \N__9938\ : std_logic;
signal \N__9937\ : std_logic;
signal \N__9934\ : std_logic;
signal \N__9929\ : std_logic;
signal \N__9924\ : std_logic;
signal \N__9923\ : std_logic;
signal \N__9920\ : std_logic;
signal \N__9917\ : std_logic;
signal \N__9912\ : std_logic;
signal \N__9911\ : std_logic;
signal \N__9908\ : std_logic;
signal \N__9905\ : std_logic;
signal \N__9902\ : std_logic;
signal \N__9897\ : std_logic;
signal \N__9896\ : std_logic;
signal \N__9895\ : std_logic;
signal \N__9892\ : std_logic;
signal \N__9887\ : std_logic;
signal \N__9882\ : std_logic;
signal \N__9881\ : std_logic;
signal \N__9878\ : std_logic;
signal \N__9875\ : std_logic;
signal \N__9870\ : std_logic;
signal \N__9867\ : std_logic;
signal \N__9864\ : std_logic;
signal \N__9861\ : std_logic;
signal \N__9858\ : std_logic;
signal \N__9857\ : std_logic;
signal \N__9854\ : std_logic;
signal \N__9851\ : std_logic;
signal \N__9848\ : std_logic;
signal \N__9843\ : std_logic;
signal \N__9842\ : std_logic;
signal \N__9839\ : std_logic;
signal \N__9836\ : std_logic;
signal \N__9831\ : std_logic;
signal \N__9830\ : std_logic;
signal \N__9827\ : std_logic;
signal \N__9824\ : std_logic;
signal \N__9819\ : std_logic;
signal \N__9818\ : std_logic;
signal \N__9815\ : std_logic;
signal \N__9812\ : std_logic;
signal \N__9809\ : std_logic;
signal \N__9804\ : std_logic;
signal \N__9803\ : std_logic;
signal \N__9800\ : std_logic;
signal \N__9797\ : std_logic;
signal \N__9792\ : std_logic;
signal \N__9789\ : std_logic;
signal \N__9786\ : std_logic;
signal \N__9785\ : std_logic;
signal \N__9784\ : std_logic;
signal \N__9781\ : std_logic;
signal \N__9778\ : std_logic;
signal \N__9775\ : std_logic;
signal \N__9768\ : std_logic;
signal \N__9767\ : std_logic;
signal \N__9764\ : std_logic;
signal \N__9763\ : std_logic;
signal \N__9760\ : std_logic;
signal \N__9757\ : std_logic;
signal \N__9754\ : std_logic;
signal \N__9747\ : std_logic;
signal \N__9744\ : std_logic;
signal \N__9741\ : std_logic;
signal \N__9738\ : std_logic;
signal \N__9737\ : std_logic;
signal \N__9732\ : std_logic;
signal \N__9729\ : std_logic;
signal \N__9726\ : std_logic;
signal \N__9723\ : std_logic;
signal \N__9720\ : std_logic;
signal \N__9717\ : std_logic;
signal \N__9714\ : std_logic;
signal \N__9711\ : std_logic;
signal \N__9708\ : std_logic;
signal \N__9707\ : std_logic;
signal \N__9704\ : std_logic;
signal \N__9701\ : std_logic;
signal \N__9696\ : std_logic;
signal \N__9693\ : std_logic;
signal \N__9690\ : std_logic;
signal \N__9687\ : std_logic;
signal \N__9686\ : std_logic;
signal \N__9683\ : std_logic;
signal \N__9680\ : std_logic;
signal \N__9675\ : std_logic;
signal \N__9672\ : std_logic;
signal \N__9669\ : std_logic;
signal \N__9666\ : std_logic;
signal \N__9663\ : std_logic;
signal \N__9660\ : std_logic;
signal \N__9657\ : std_logic;
signal \N__9654\ : std_logic;
signal \N__9651\ : std_logic;
signal \N__9648\ : std_logic;
signal \N__9645\ : std_logic;
signal \N__9642\ : std_logic;
signal \N__9639\ : std_logic;
signal \N__9636\ : std_logic;
signal \N__9633\ : std_logic;
signal \N__9630\ : std_logic;
signal \N__9627\ : std_logic;
signal \N__9624\ : std_logic;
signal \N__9621\ : std_logic;
signal \N__9618\ : std_logic;
signal \N__9615\ : std_logic;
signal \N__9612\ : std_logic;
signal \N__9609\ : std_logic;
signal \N__9606\ : std_logic;
signal \N__9603\ : std_logic;
signal \N__9600\ : std_logic;
signal \N__9597\ : std_logic;
signal \N__9594\ : std_logic;
signal \N__9591\ : std_logic;
signal \N__9588\ : std_logic;
signal \N__9585\ : std_logic;
signal \N__9582\ : std_logic;
signal \N__9579\ : std_logic;
signal \N__9576\ : std_logic;
signal \N__9573\ : std_logic;
signal \N__9570\ : std_logic;
signal \N__9567\ : std_logic;
signal \N__9564\ : std_logic;
signal \N__9561\ : std_logic;
signal \N__9558\ : std_logic;
signal \N__9555\ : std_logic;
signal \N__9552\ : std_logic;
signal \N__9549\ : std_logic;
signal \N__9546\ : std_logic;
signal \N__9543\ : std_logic;
signal \N__9540\ : std_logic;
signal \N__9537\ : std_logic;
signal \N__9534\ : std_logic;
signal \N__9533\ : std_logic;
signal \N__9528\ : std_logic;
signal \N__9525\ : std_logic;
signal \N__9522\ : std_logic;
signal \N__9519\ : std_logic;
signal \N__9516\ : std_logic;
signal \N__9515\ : std_logic;
signal \N__9510\ : std_logic;
signal \N__9507\ : std_logic;
signal \N__9504\ : std_logic;
signal \N__9501\ : std_logic;
signal \N__9498\ : std_logic;
signal \N__9497\ : std_logic;
signal \N__9494\ : std_logic;
signal \N__9491\ : std_logic;
signal \N__9486\ : std_logic;
signal \N__9483\ : std_logic;
signal \N__9480\ : std_logic;
signal \N__9477\ : std_logic;
signal \N__9474\ : std_logic;
signal \N__9471\ : std_logic;
signal \N__9468\ : std_logic;
signal \N__9465\ : std_logic;
signal \N__9462\ : std_logic;
signal \N__9459\ : std_logic;
signal \N__9456\ : std_logic;
signal \N__9453\ : std_logic;
signal \N__9450\ : std_logic;
signal \N__9447\ : std_logic;
signal \N__9446\ : std_logic;
signal \N__9441\ : std_logic;
signal \N__9438\ : std_logic;
signal \N__9435\ : std_logic;
signal \N__9432\ : std_logic;
signal \N__9429\ : std_logic;
signal \N__9428\ : std_logic;
signal \N__9423\ : std_logic;
signal \N__9420\ : std_logic;
signal \N__9417\ : std_logic;
signal \N__9414\ : std_logic;
signal \N__9411\ : std_logic;
signal \N__9410\ : std_logic;
signal \N__9405\ : std_logic;
signal \N__9402\ : std_logic;
signal \N__9399\ : std_logic;
signal \N__9396\ : std_logic;
signal \N__9393\ : std_logic;
signal \N__9392\ : std_logic;
signal \N__9387\ : std_logic;
signal \N__9384\ : std_logic;
signal \N__9381\ : std_logic;
signal \N__9378\ : std_logic;
signal \N__9375\ : std_logic;
signal \N__9372\ : std_logic;
signal \N__9369\ : std_logic;
signal \N__9366\ : std_logic;
signal \N__9363\ : std_logic;
signal \N__9360\ : std_logic;
signal \N__9357\ : std_logic;
signal \N__9354\ : std_logic;
signal \N__9351\ : std_logic;
signal \N__9348\ : std_logic;
signal \N__9345\ : std_logic;
signal \N__9342\ : std_logic;
signal \N__9339\ : std_logic;
signal \N__9336\ : std_logic;
signal \N__9333\ : std_logic;
signal \N__9330\ : std_logic;
signal \N__9327\ : std_logic;
signal \N__9324\ : std_logic;
signal \N__9321\ : std_logic;
signal \N__9318\ : std_logic;
signal \N__9315\ : std_logic;
signal \N__9312\ : std_logic;
signal \N__9309\ : std_logic;
signal \N__9306\ : std_logic;
signal \N__9305\ : std_logic;
signal \N__9302\ : std_logic;
signal \N__9299\ : std_logic;
signal \N__9294\ : std_logic;
signal \N__9291\ : std_logic;
signal \N__9288\ : std_logic;
signal \N__9285\ : std_logic;
signal \N__9284\ : std_logic;
signal \N__9279\ : std_logic;
signal \N__9276\ : std_logic;
signal \N__9273\ : std_logic;
signal \N__9272\ : std_logic;
signal \N__9269\ : std_logic;
signal \N__9264\ : std_logic;
signal \N__9261\ : std_logic;
signal \N__9258\ : std_logic;
signal \N__9257\ : std_logic;
signal \N__9254\ : std_logic;
signal \N__9251\ : std_logic;
signal \N__9246\ : std_logic;
signal \N__9243\ : std_logic;
signal \N__9240\ : std_logic;
signal \N__9237\ : std_logic;
signal \N__9234\ : std_logic;
signal \N__9231\ : std_logic;
signal \N__9228\ : std_logic;
signal \N__9225\ : std_logic;
signal \N__9222\ : std_logic;
signal \N__9219\ : std_logic;
signal \N__9216\ : std_logic;
signal \N__9213\ : std_logic;
signal \N__9210\ : std_logic;
signal \N__9207\ : std_logic;
signal \N__9204\ : std_logic;
signal \N__9201\ : std_logic;
signal \N__9198\ : std_logic;
signal \N__9195\ : std_logic;
signal \N__9192\ : std_logic;
signal \N__9189\ : std_logic;
signal \N__9186\ : std_logic;
signal \N__9183\ : std_logic;
signal \N__9180\ : std_logic;
signal \N__9177\ : std_logic;
signal \N__9174\ : std_logic;
signal \N__9171\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \uart_frame_decoder.WDTZ0Z_0\ : std_logic;
signal \bfn_1_17_0_\ : std_logic;
signal \uart_frame_decoder.WDTZ0Z_1\ : std_logic;
signal \uart_frame_decoder.un1_WDT_cry_0\ : std_logic;
signal \uart_frame_decoder.WDTZ0Z_2\ : std_logic;
signal \uart_frame_decoder.un1_WDT_cry_1\ : std_logic;
signal \uart_frame_decoder.WDTZ0Z_3\ : std_logic;
signal \uart_frame_decoder.un1_WDT_cry_2\ : std_logic;
signal \uart_frame_decoder.un1_WDT_cry_3\ : std_logic;
signal \uart_frame_decoder.un1_WDT_cry_4\ : std_logic;
signal \uart_frame_decoder.un1_WDT_cry_5\ : std_logic;
signal \uart_frame_decoder.un1_WDT_cry_6\ : std_logic;
signal \uart_frame_decoder.un1_WDT_cry_7\ : std_logic;
signal \bfn_1_18_0_\ : std_logic;
signal \uart_frame_decoder.un1_WDT_cry_8\ : std_logic;
signal \uart_frame_decoder.un1_WDT_cry_9\ : std_logic;
signal \uart_frame_decoder.un1_WDT_cry_10\ : std_logic;
signal \uart_frame_decoder.un1_WDT_cry_11\ : std_logic;
signal \uart_frame_decoder.un1_WDT_cry_12\ : std_logic;
signal \uart_frame_decoder.un1_WDT_cry_13\ : std_logic;
signal \uart_frame_decoder.un1_WDT_cry_14\ : std_logic;
signal \bfn_1_19_0_\ : std_logic;
signal \uart_frame_decoder.count8_axb_1\ : std_logic;
signal \uart_frame_decoder.count8_cry_0\ : std_logic;
signal \uart_frame_decoder.count_i_2\ : std_logic;
signal \uart_frame_decoder.count8_cry_1\ : std_logic;
signal \uart_frame_decoder.count8\ : std_logic;
signal \uart_frame_decoder.count8_cry_2_c_RNICKSZ0Z21\ : std_logic;
signal \uart_frame_decoder.count8_cry_2_c_RNICKSZ0Z21_cascade_\ : std_logic;
signal \uart_frame_decoder.count_RNIV5MSZ0Z_0\ : std_logic;
signal \uart_frame_decoder.source_data_valid_2_sqmuxa_iZ0\ : std_logic;
signal \uart_frame_decoder.count8_0_i\ : std_logic;
signal \bfn_1_23_0_\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_0\ : std_logic;
signal \frame_decoder_OFF3data_2\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_1\ : std_logic;
signal \frame_decoder_OFF3data_3\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_2\ : std_logic;
signal \frame_decoder_OFF3data_4\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_3\ : std_logic;
signal \frame_decoder_OFF3data_5\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_4\ : std_logic;
signal \frame_decoder_OFF3data_6\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_5\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_6\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_7\ : std_logic;
signal \bfn_1_24_0_\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_8\ : std_logic;
signal \scaler_3.N_795_i_l_ofxZ0\ : std_logic;
signal \scaler_3.un2_source_data_0_cry_1_c_RNO_1\ : std_logic;
signal \bfn_1_25_0_\ : std_logic;
signal \scaler_3.un2_source_data_0_cry_1\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_1_c_RNIOS6I\ : std_logic;
signal \scaler_3.un2_source_data_0_cry_2\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_2_c_RNIR08I\ : std_logic;
signal \scaler_3.un2_source_data_0_cry_3\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_3_c_RNIU49I\ : std_logic;
signal \scaler_3.un2_source_data_0_cry_4\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_4_c_RNI19AI\ : std_logic;
signal \scaler_3.un2_source_data_0_cry_5\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_5_c_RNI4DBI\ : std_logic;
signal \scaler_3.un2_source_data_0_cry_6\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_6_c_RNI7HCI\ : std_logic;
signal \scaler_3.un2_source_data_0_cry_7\ : std_logic;
signal \scaler_3.un2_source_data_0_cry_8\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_7_c_RNI8JDI\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_8_c_RNIRV25\ : std_logic;
signal \bfn_1_26_0_\ : std_logic;
signal \scaler_3.un2_source_data_0_cry_9\ : std_logic;
signal \uart_frame_decoder.source_offset4data_1_sqmuxa_0\ : std_logic;
signal \bfn_1_29_0_\ : std_logic;
signal \frame_decoder_CH4data_1\ : std_logic;
signal \frame_decoder_OFF4data_1\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_0\ : std_logic;
signal \frame_decoder_CH4data_2\ : std_logic;
signal \frame_decoder_OFF4data_2\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_1\ : std_logic;
signal \frame_decoder_CH4data_3\ : std_logic;
signal \frame_decoder_OFF4data_3\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_2\ : std_logic;
signal \frame_decoder_CH4data_4\ : std_logic;
signal \frame_decoder_OFF4data_4\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_3\ : std_logic;
signal \frame_decoder_OFF4data_5\ : std_logic;
signal \frame_decoder_CH4data_5\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_4\ : std_logic;
signal \frame_decoder_CH4data_6\ : std_logic;
signal \frame_decoder_OFF4data_6\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_5\ : std_logic;
signal \scaler_4.un3_source_data_0_axb_7\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_6\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_7\ : std_logic;
signal \bfn_1_30_0_\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_8\ : std_logic;
signal \frame_decoder_OFF4data_7\ : std_logic;
signal \scaler_4.N_807_i_l_ofxZ0\ : std_logic;
signal \uart_frame_decoder.WDTZ0Z_8\ : std_logic;
signal \uart_frame_decoder.WDTZ0Z_11\ : std_logic;
signal \uart_frame_decoder.WDTZ0Z_10\ : std_logic;
signal \uart_frame_decoder.WDTZ0Z_13\ : std_logic;
signal \uart_frame_decoder.WDTZ0Z_12\ : std_logic;
signal \uart_frame_decoder.WDTZ0Z_9\ : std_logic;
signal \uart_frame_decoder.WDT_RNIAGPBZ0Z_10_cascade_\ : std_logic;
signal \uart_frame_decoder.WDT8lto13_1\ : std_logic;
signal \uart_frame_decoder.WDT8lt14_0_cascade_\ : std_logic;
signal \uart_frame_decoder.WDT8_0_i\ : std_logic;
signal \uart_frame_decoder.WDTZ0Z_6\ : std_logic;
signal \uart_frame_decoder.WDTZ0Z_5\ : std_logic;
signal \uart_frame_decoder.WDTZ0Z_7\ : std_logic;
signal \uart_frame_decoder.WDTZ0Z_4\ : std_logic;
signal \uart_frame_decoder.WDT_RNIM6B11Z0Z_4\ : std_logic;
signal \uart_frame_decoder.WDTZ0Z_15\ : std_logic;
signal \uart_frame_decoder.WDTZ0Z_14\ : std_logic;
signal \uart_frame_decoder.WDT8lt14_0\ : std_logic;
signal \uart_frame_decoder.WDT_RNIJUEI2Z0Z_15_cascade_\ : std_logic;
signal \uart_frame_decoder.state_1Z0Z_3\ : std_logic;
signal \uart_frame_decoder.state_1Z0Z_2\ : std_logic;
signal \uart_frame_decoder.state_1Z0Z_4\ : std_logic;
signal \uart_frame_decoder.countZ0Z_2\ : std_logic;
signal \uart_frame_decoder.countZ0Z_1\ : std_logic;
signal \uart_frame_decoder.count8_0\ : std_logic;
signal \uart_frame_decoder.state_1_ns_i_i_0_0_cascade_\ : std_logic;
signal \bfn_2_21_0_\ : std_logic;
signal \frame_decoder_CH2data_1\ : std_logic;
signal \frame_decoder_OFF2data_1\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_0\ : std_logic;
signal \frame_decoder_CH2data_2\ : std_logic;
signal \frame_decoder_OFF2data_2\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_1\ : std_logic;
signal \frame_decoder_CH2data_3\ : std_logic;
signal \frame_decoder_OFF2data_3\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_2\ : std_logic;
signal \frame_decoder_CH2data_4\ : std_logic;
signal \frame_decoder_OFF2data_4\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_3\ : std_logic;
signal \frame_decoder_CH2data_5\ : std_logic;
signal \frame_decoder_OFF2data_5\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_4\ : std_logic;
signal \frame_decoder_CH2data_6\ : std_logic;
signal \frame_decoder_OFF2data_6\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_5\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_6\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_7\ : std_logic;
signal \bfn_2_22_0_\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_8\ : std_logic;
signal \scaler_2.un3_source_data_0_axb_7\ : std_logic;
signal \uart_frame_decoder.source_CH1data_1_sqmuxa\ : std_logic;
signal \uart_frame_decoder.source_offset2data_1_sqmuxa_0\ : std_logic;
signal \frame_decoder_CH2data_7\ : std_logic;
signal \frame_decoder_OFF2data_7\ : std_logic;
signal \scaler_2.N_783_i_l_ofxZ0\ : std_logic;
signal \uart_frame_decoder.source_CH2data_1_sqmuxa\ : std_logic;
signal \uart_frame_decoder.source_CH2data_1_sqmuxa_0\ : std_logic;
signal \uart_frame_decoder.source_CH4data_1_sqmuxa_cascade_\ : std_logic;
signal \frame_decoder_OFF3data_7\ : std_logic;
signal \scaler_3.un3_source_data_0_axb_7\ : std_logic;
signal \uart_frame_decoder.source_offset3data_1_sqmuxa_cascade_\ : std_logic;
signal \frame_decoder_CH3data_1\ : std_logic;
signal \frame_decoder_CH3data_2\ : std_logic;
signal \frame_decoder_CH3data_3\ : std_logic;
signal \frame_decoder_CH3data_4\ : std_logic;
signal \frame_decoder_CH3data_5\ : std_logic;
signal \frame_decoder_CH3data_6\ : std_logic;
signal \frame_decoder_CH3data_7\ : std_logic;
signal \bfn_2_27_0_\ : std_logic;
signal \frame_decoder_CH1data_1\ : std_logic;
signal \frame_decoder_OFF1data_1\ : std_logic;
signal \scaler_1.un3_source_data_0_cry_0\ : std_logic;
signal \frame_decoder_CH1data_2\ : std_logic;
signal \frame_decoder_OFF1data_2\ : std_logic;
signal \scaler_1.un3_source_data_0_cry_1\ : std_logic;
signal \frame_decoder_CH1data_3\ : std_logic;
signal \frame_decoder_OFF1data_3\ : std_logic;
signal \scaler_1.un3_source_data_0_cry_2\ : std_logic;
signal \frame_decoder_OFF1data_4\ : std_logic;
signal \scaler_1.un3_source_data_0_cry_3\ : std_logic;
signal \frame_decoder_CH1data_5\ : std_logic;
signal \frame_decoder_OFF1data_5\ : std_logic;
signal \scaler_1.un3_source_data_0_cry_4\ : std_logic;
signal \frame_decoder_OFF1data_6\ : std_logic;
signal \frame_decoder_CH1data_6\ : std_logic;
signal \scaler_1.un3_source_data_0_cry_5\ : std_logic;
signal \scaler_1.un3_source_data_0_cry_6\ : std_logic;
signal \scaler_1.un3_source_data_0_cry_7\ : std_logic;
signal \bfn_2_28_0_\ : std_logic;
signal \scaler_1.un3_source_data_0_cry_8\ : std_logic;
signal \scaler_1.N_771_i_l_ofxZ0\ : std_logic;
signal \frame_decoder_CH4data_0\ : std_logic;
signal \frame_decoder_OFF4data_0\ : std_logic;
signal \scaler_4.un2_source_data_0_cry_1_c_RNO_2\ : std_logic;
signal \bfn_2_29_0_\ : std_logic;
signal \scaler_4.un2_source_data_0\ : std_logic;
signal \scaler_4.un2_source_data_0_cry_1\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_1_c_RNIRSJI\ : std_logic;
signal \scaler_4.un2_source_data_0_cry_2\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_2_c_RNIU0LI\ : std_logic;
signal \scaler_4.un2_source_data_0_cry_3\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_3_c_RNI15MI\ : std_logic;
signal \scaler_4.un2_source_data_0_cry_4\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_4_c_RNI49NI\ : std_logic;
signal \scaler_4.un2_source_data_0_cry_5\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_5_c_RNI7DOI\ : std_logic;
signal \scaler_4.un2_source_data_0_cry_6\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_6_c_RNIAHPI\ : std_logic;
signal \scaler_4.un2_source_data_0_cry_7\ : std_logic;
signal \scaler_4.un2_source_data_0_cry_8\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_7_c_RNIBJQI\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_8_c_RNIS918\ : std_logic;
signal \bfn_2_30_0_\ : std_logic;
signal \scaler_4.un2_source_data_0_cry_9\ : std_logic;
signal \uart.CO1\ : std_logic;
signal \uart.N_133_0\ : std_logic;
signal \uart.N_177_cascade_\ : std_logic;
signal \uart.state_srsts_i_0_3\ : std_logic;
signal \uart.N_168_1_cascade_\ : std_logic;
signal \uart.N_154_0\ : std_logic;
signal \uart.data_Auxce_0_0_0\ : std_logic;
signal \uart.data_Auxce_0_1\ : std_logic;
signal \uart.data_Auxce_0_3\ : std_logic;
signal \uart.data_Auxce_0_5\ : std_logic;
signal \uart.data_Auxce_0_6\ : std_logic;
signal \uart.N_177\ : std_logic;
signal \uart.state_srsts_0_0_0_cascade_\ : std_logic;
signal \uart_frame_decoder.state_1_RNI592GZ0Z_10\ : std_logic;
signal \uart_frame_decoder.state_1_RNO_3Z0Z_0\ : std_logic;
signal \uart_frame_decoder.N_168_i_1\ : std_logic;
signal \uart_frame_decoder.state_1_RNO_2Z0Z_0\ : std_logic;
signal \uart_frame_decoder.state_1Z0Z_7\ : std_logic;
signal \uart_frame_decoder.state_1Z0Z_0\ : std_logic;
signal \uart_frame_decoder.N_79_4\ : std_logic;
signal \uart_frame_decoder.state_1_ns_0_i_a2_0_0_1\ : std_logic;
signal \uart.data_AuxZ1Z_0\ : std_logic;
signal uart_data_0 : std_logic;
signal \uart_frame_decoder.state_1Z0Z_1\ : std_logic;
signal \uart_frame_decoder.state_1_ns_0_i_a2_0_0_1Z0Z_2_cascade_\ : std_logic;
signal \uart_frame_decoder.state_1_ns_0_i_a2_0_2\ : std_logic;
signal \uart.data_AuxZ0Z_5\ : std_logic;
signal uart_data_5 : std_logic;
signal \uart.data_AuxZ1Z_2\ : std_logic;
signal uart_data_2 : std_logic;
signal \uart.data_AuxZ0Z_7\ : std_logic;
signal \uart.data_AuxZ1Z_1\ : std_logic;
signal \bfn_3_21_0_\ : std_logic;
signal \scaler_2.un2_source_data_0_cry_1\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_1_c_RNILSPH\ : std_logic;
signal \scaler_2.un2_source_data_0_cry_2\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_2_c_RNIO0RH\ : std_logic;
signal \scaler_2.un2_source_data_0_cry_3\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_3_c_RNIR4SH\ : std_logic;
signal \scaler_2.un2_source_data_0_cry_4\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_4_c_RNIU8TH\ : std_logic;
signal \scaler_2.un2_source_data_0_cry_5\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_5_c_RNI1DUH\ : std_logic;
signal \scaler_2.un2_source_data_0_cry_6\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_6_c_RNI4HVH\ : std_logic;
signal \scaler_2.un2_source_data_0_cry_7\ : std_logic;
signal \scaler_2.un2_source_data_0_cry_8\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_7_c_RNI5J0I\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_8_c_RNIQL42\ : std_logic;
signal \bfn_3_22_0_\ : std_logic;
signal \scaler_2.un2_source_data_0_cry_9\ : std_logic;
signal \scaler_3.un2_source_data_0\ : std_logic;
signal \uart_frame_decoder.source_offset2data_1_sqmuxa\ : std_logic;
signal \uart_frame_decoder.state_1Z0Z_8\ : std_logic;
signal \uart_frame_decoder.source_offset3data_1_sqmuxa\ : std_logic;
signal \uart_frame_decoder.state_1Z0Z_9\ : std_logic;
signal \uart_frame_decoder.state_1Z0Z_5\ : std_logic;
signal \uart_frame_decoder.source_CH4data_1_sqmuxa\ : std_logic;
signal uart_data_7 : std_logic;
signal \frame_decoder_CH4data_7\ : std_logic;
signal \uart_frame_decoder.source_CH4data_1_sqmuxa_0\ : std_logic;
signal \uart_frame_decoder.source_CH3data_1_sqmuxa\ : std_logic;
signal \uart_frame_decoder.source_CH3data_1_sqmuxa_0\ : std_logic;
signal \frame_decoder_OFF1data_0\ : std_logic;
signal \frame_decoder_CH1data_0\ : std_logic;
signal \frame_decoder_OFF1data_7\ : std_logic;
signal \frame_decoder_CH1data_7\ : std_logic;
signal \scaler_1.un3_source_data_0_axb_7\ : std_logic;
signal \bfn_3_26_0_\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_6\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_7\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_8\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_9\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_10\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_11\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_12\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_13\ : std_logic;
signal scaler_4_data_14 : std_logic;
signal \bfn_3_27_0_\ : std_logic;
signal \scaler_1.un2_source_data_0_cry_1_c_RNOZ0\ : std_logic;
signal \bfn_3_28_0_\ : std_logic;
signal \scaler_1.un2_source_data_0\ : std_logic;
signal \scaler_1.un2_source_data_0_cry_1\ : std_logic;
signal \scaler_1.un3_source_data_0_cry_1_c_RNIISC11\ : std_logic;
signal \scaler_1.un2_source_data_0_cry_2\ : std_logic;
signal \scaler_1.un3_source_data_0_cry_2_c_RNIL0E11\ : std_logic;
signal \scaler_1.un2_source_data_0_cry_3\ : std_logic;
signal \scaler_1.un3_source_data_0_cry_3_c_RNIO4F11\ : std_logic;
signal \scaler_1.un2_source_data_0_cry_4\ : std_logic;
signal \scaler_1.un3_source_data_0_cry_4_c_RNIR8G11\ : std_logic;
signal \scaler_1.un2_source_data_0_cry_5\ : std_logic;
signal \scaler_1.un3_source_data_0_cry_5_c_RNIUCH11\ : std_logic;
signal \scaler_1.un2_source_data_0_cry_6\ : std_logic;
signal \scaler_1.un3_source_data_0_cry_6_c_RNI1HI11\ : std_logic;
signal \scaler_1.un2_source_data_0_cry_7\ : std_logic;
signal \scaler_1.un2_source_data_0_cry_8\ : std_logic;
signal \scaler_1.un3_source_data_0_cry_7_c_RNI2JJ11\ : std_logic;
signal \scaler_1.un3_source_data_0_cry_8_c_RNIPB6F\ : std_logic;
signal \bfn_3_29_0_\ : std_logic;
signal \scaler_1.un2_source_data_0_cry_9\ : std_logic;
signal frame_decoder_dv_c_0_g : std_logic;
signal \frame_decoder_OFF3data_1\ : std_logic;
signal \uart_frame_decoder.source_offset3data_1_sqmuxa_0\ : std_logic;
signal \uart_sync.aux_2__0_Z0Z_0\ : std_logic;
signal \uart_sync.aux_3__0_Z0Z_0\ : std_logic;
signal \uart.N_151\ : std_logic;
signal \uart.stateZ0Z_2\ : std_logic;
signal \uart.N_159\ : std_logic;
signal \uart.timer_Count_0_sqmuxa_1_cascade_\ : std_logic;
signal \uart.N_180\ : std_logic;
signal \uart.N_180_cascade_\ : std_logic;
signal \uart.un1_state_5_0\ : std_logic;
signal \uart.N_143_0\ : std_logic;
signal \reset_module_System.count_1_1_cascade_\ : std_logic;
signal \uart.N_153_0_cascade_\ : std_logic;
signal \uart.state_srsts_i_a3_0_0_3_cascade_\ : std_logic;
signal \uart.N_170\ : std_logic;
signal \uart.un1_state_2_0_a3_2\ : std_logic;
signal \uart.N_146_0\ : std_logic;
signal \uart.un1_state_2_0\ : std_logic;
signal \reset_module_System.reset6_11_cascade_\ : std_logic;
signal \reset_module_System.reset6_19\ : std_logic;
signal \reset_module_System.reset6_19_cascade_\ : std_logic;
signal \uart.data_Auxce_0_0_4\ : std_logic;
signal \reset_module_System.reset6_14\ : std_logic;
signal \uart.state_RNIAFHLZ0Z_3\ : std_logic;
signal \uart.N_153_0\ : std_logic;
signal \uart.stateZ0Z_3\ : std_logic;
signal \uart.N_168_1\ : std_logic;
signal \uart.N_167\ : std_logic;
signal \uart.stateZ0Z_4\ : std_logic;
signal \uart.bit_CountZ0Z_2\ : std_logic;
signal \uart.bit_CountZ0Z_1\ : std_logic;
signal \uart.bit_CountZ0Z_0\ : std_logic;
signal \uart.data_Auxce_0_0_2\ : std_logic;
signal \reset_module_System.reset6_13\ : std_logic;
signal \reset_module_System.reset6_3\ : std_logic;
signal \reset_module_System.reset6_17\ : std_logic;
signal uart_data_1 : std_logic;
signal \uart_frame_decoder.state_1_ns_0_i_a2_1_1Z0Z_2_cascade_\ : std_logic;
signal \uart_frame_decoder.state_1_ns_0_i_a2_1Z0Z_2\ : std_logic;
signal \uart.stateZ0Z_0\ : std_logic;
signal \uart.stateZ0Z_1\ : std_logic;
signal uart_input_sync : std_logic;
signal \uart.data_AuxZ0Z_3\ : std_logic;
signal uart_data_3 : std_logic;
signal \uart.data_AuxZ0Z_6\ : std_logic;
signal uart_data_6 : std_logic;
signal \uart_frame_decoder.state_1Z0Z_6\ : std_logic;
signal \uart_frame_decoder.source_offset1data_1_sqmuxa\ : std_logic;
signal \uart_frame_decoder.source_offset1data_1_sqmuxa_cascade_\ : std_logic;
signal \uart_frame_decoder.source_offset1data_1_sqmuxa_0\ : std_logic;
signal \uart.data_rdyc_1\ : std_logic;
signal \uart.data_AuxZ0Z_4\ : std_logic;
signal \uart.state_RNIQABT2Z0Z_4\ : std_logic;
signal \uart_frame_decoder.state_1_ns_0_i_o2_0_10\ : std_logic;
signal \uart_frame_decoder.source_offset4data_1_sqmuxa\ : std_logic;
signal \uart_frame_decoder.WDT_RNIJUEI2Z0Z_15\ : std_logic;
signal scaler_4_data_11 : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_10_THRU_CO\ : std_logic;
signal \uart_frame_decoder.state_1Z0Z_10\ : std_logic;
signal uart_data_rdy : std_logic;
signal \uart_frame_decoder.count8_THRU_CO\ : std_logic;
signal scaler_4_data_6 : std_logic;
signal \frame_decoder_OFF3data_0\ : std_logic;
signal \frame_decoder_CH3data_0\ : std_logic;
signal \bfn_4_24_0_\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_6\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_7\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_8\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_9\ : std_logic;
signal scaler_2_data_11 : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_10_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_10\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_11\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_12\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_13\ : std_logic;
signal scaler_2_data_14 : std_logic;
signal \bfn_4_25_0_\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_9_THRU_CO\ : std_logic;
signal scaler_4_data_10 : std_logic;
signal scaler_2_data_10 : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_9_THRU_CO\ : std_logic;
signal scaler_4_data_13 : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_12_THRU_CO\ : std_logic;
signal scaler_3_data_6 : std_logic;
signal \bfn_4_27_0_\ : std_logic;
signal scaler_3_data_7 : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_6_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_6\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_7\ : std_logic;
signal scaler_3_data_9 : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_8_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_8\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_9\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_10\ : std_logic;
signal scaler_3_data_12 : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_11_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_11\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_12\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_13\ : std_logic;
signal scaler_3_data_14 : std_logic;
signal \bfn_4_28_0_\ : std_logic;
signal scaler_1_data_6 : std_logic;
signal \bfn_4_29_0_\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_6\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_7\ : std_logic;
signal scaler_1_data_9 : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_8_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_8\ : std_logic;
signal scaler_1_data_10 : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_9_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_9\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_10\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_11\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_12\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_13\ : std_logic;
signal scaler_1_data_14 : std_logic;
signal \bfn_4_30_0_\ : std_logic;
signal \uart_sync.aux_1__0_Z0Z_0\ : std_logic;
signal \uart.timer_CountZ0Z_1\ : std_logic;
signal \bfn_5_15_0_\ : std_logic;
signal \uart.timer_CountZ0Z_2\ : std_logic;
signal \uart.un4_timer_Count_1_cry_1\ : std_logic;
signal \uart.timer_CountZ0Z_3\ : std_logic;
signal \uart.un4_timer_Count_1_cry_2\ : std_logic;
signal \uart.un4_timer_Count_1_cry_3\ : std_logic;
signal \uart.timer_CountZ0Z_5\ : std_logic;
signal \uart.un4_timer_Count_1_cry_4\ : std_logic;
signal \uart.timer_CountZ0Z_6\ : std_logic;
signal \uart.un4_timer_Count_1_cry_5\ : std_logic;
signal \uart.un4_timer_Count_1_cry_6\ : std_logic;
signal \uart.timer_CountZ0Z_7\ : std_logic;
signal \uart.timer_Count_1_sqmuxa_i\ : std_logic;
signal \uart.timer_CountZ0Z_0\ : std_logic;
signal \uart.timer_CountZ0Z_4\ : std_logic;
signal \uart.un1_state_2_0_a3_0\ : std_logic;
signal \reset_module_System.countZ0Z_0\ : std_logic;
signal \reset_module_System.countZ0Z_1\ : std_logic;
signal \bfn_5_17_0_\ : std_logic;
signal \reset_module_System.countZ0Z_2\ : std_logic;
signal \reset_module_System.count_1_2\ : std_logic;
signal \reset_module_System.count_1_cry_1\ : std_logic;
signal \reset_module_System.countZ0Z_3\ : std_logic;
signal \reset_module_System.count_1_cry_2\ : std_logic;
signal \reset_module_System.countZ0Z_4\ : std_logic;
signal \reset_module_System.count_1_cry_3\ : std_logic;
signal \reset_module_System.countZ0Z_5\ : std_logic;
signal \reset_module_System.count_1_cry_4\ : std_logic;
signal \reset_module_System.countZ0Z_6\ : std_logic;
signal \reset_module_System.count_1_cry_5\ : std_logic;
signal \reset_module_System.countZ0Z_7\ : std_logic;
signal \reset_module_System.count_1_cry_6\ : std_logic;
signal \reset_module_System.countZ0Z_8\ : std_logic;
signal \reset_module_System.count_1_cry_7\ : std_logic;
signal \reset_module_System.count_1_cry_8\ : std_logic;
signal \reset_module_System.countZ0Z_9\ : std_logic;
signal \bfn_5_18_0_\ : std_logic;
signal \reset_module_System.countZ0Z_10\ : std_logic;
signal \reset_module_System.count_1_cry_9\ : std_logic;
signal \reset_module_System.countZ0Z_11\ : std_logic;
signal \reset_module_System.count_1_cry_10\ : std_logic;
signal \reset_module_System.countZ0Z_12\ : std_logic;
signal \reset_module_System.count_1_cry_11\ : std_logic;
signal \reset_module_System.count_1_cry_12\ : std_logic;
signal \reset_module_System.countZ0Z_14\ : std_logic;
signal \reset_module_System.count_1_cry_13\ : std_logic;
signal \reset_module_System.count_1_cry_14\ : std_logic;
signal \reset_module_System.countZ0Z_16\ : std_logic;
signal \reset_module_System.count_1_cry_15\ : std_logic;
signal \reset_module_System.count_1_cry_16\ : std_logic;
signal \reset_module_System.countZ0Z_17\ : std_logic;
signal \bfn_5_19_0_\ : std_logic;
signal \reset_module_System.countZ0Z_18\ : std_logic;
signal \reset_module_System.count_1_cry_17\ : std_logic;
signal \reset_module_System.count_1_cry_18\ : std_logic;
signal \reset_module_System.countZ0Z_20\ : std_logic;
signal \reset_module_System.count_1_cry_19\ : std_logic;
signal \reset_module_System.count_1_cry_20\ : std_logic;
signal \reset_module_System.countZ0Z_19\ : std_logic;
signal \reset_module_System.countZ0Z_15\ : std_logic;
signal \reset_module_System.countZ0Z_21\ : std_logic;
signal \reset_module_System.countZ0Z_13\ : std_logic;
signal \reset_module_System.reset6_15\ : std_logic;
signal scaler_3_data_4 : std_logic;
signal \scaler_2.un2_source_data_0\ : std_logic;
signal \scaler_2.un2_source_data_0_cry_1_c_RNO_0\ : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_4\ : std_logic;
signal \ppm_encoder_1.aileronZ0Z_4\ : std_logic;
signal scaler_2_data_6 : std_logic;
signal \ppm_encoder_1.aileronZ0Z_6\ : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_6\ : std_logic;
signal \ppm_encoder_1.pulses2count_9_0_o2_0_6_cascade_\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_rn_0_6\ : std_logic;
signal \ppm_encoder_1.un2_throttle_0_6_cascade_\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_axb_6_cascade_\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_sn_6\ : std_logic;
signal \ppm_encoder_1.N_415\ : std_logic;
signal \ppm_encoder_1.N_414_cascade_\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_1_10_cascade_\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_axb_10_cascade_\ : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_9\ : std_logic;
signal \ppm_encoder_1.N_412\ : std_logic;
signal \ppm_encoder_1.N_411_cascade_\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_1_9_cascade_\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_axb_9\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_8_THRU_CO\ : std_logic;
signal scaler_2_data_9 : std_logic;
signal \ppm_encoder_1.aileronZ0Z_9\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_8_THRU_CO\ : std_logic;
signal scaler_4_data_9 : std_logic;
signal scaler_3_data_10 : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_9_THRU_CO\ : std_logic;
signal \frame_decoder_OFF2data_0\ : std_logic;
signal \frame_decoder_CH2data_0\ : std_logic;
signal scaler_2_data_4 : std_logic;
signal scaler_4_data_12 : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_11_THRU_CO\ : std_logic;
signal uart_data_4 : std_logic;
signal \frame_decoder_CH1data_4\ : std_logic;
signal \uart_frame_decoder.source_CH1data_1_sqmuxa_0\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_11_THRU_CO\ : std_logic;
signal scaler_1_data_12 : std_logic;
signal scaler_1_data_13 : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_12_THRU_CO\ : std_logic;
signal frame_decoder_dv_c : std_logic;
signal frame_decoder_dv_c_0 : std_logic;
signal uart_input_c : std_logic;
signal \uart_sync.aux_0__0_Z0Z_0\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_6\ : std_logic;
signal \ppm_encoder_1.pulses2count_9_0_o2_0_6\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_axb_11_cascade_\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_2_11\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_i_i_1_1_4_cascade_\ : std_logic;
signal \ppm_encoder_1.N_462\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_0_cascade_\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_i_i_1_4\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_axb_4_cascade_\ : std_logic;
signal \bfn_7_23_0_\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_0\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_1\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_2\ : std_logic;
signal \ppm_encoder_1.init_pulses_RNI398E4Z0Z_4\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_4\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_3\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_4\ : std_logic;
signal \ppm_encoder_1.init_pulses_RNI6UPC6Z0Z_6\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_5\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_6\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_7\ : std_logic;
signal \bfn_7_24_0_\ : std_logic;
signal \ppm_encoder_1.init_pulses_RNI31EQ5Z0Z_9\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_8\ : std_logic;
signal \ppm_encoder_1.init_pulses_RNIJ2JB5Z0Z_10\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_9\ : std_logic;
signal \ppm_encoder_1.init_pulses_RNIV8JB5Z0Z_11\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_10\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_11\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_12\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_13\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_14\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_15\ : std_logic;
signal \bfn_7_25_0_\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_axb_17\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_16\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_17\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_axb_14_cascade_\ : std_logic;
signal \ppm_encoder_1.init_pulses_RNINK8A6Z0Z_14\ : std_logic;
signal \ppm_encoder_1.init_pulses_RNIJJM71Z0Z_15\ : std_logic;
signal \ppm_encoder_1.N_403\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_14\ : std_logic;
signal \ppm_encoder_1.N_114_cascade_\ : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_10\ : std_logic;
signal \ppm_encoder_1.aileronZ0Z_10\ : std_logic;
signal \ppm_encoder_1.N_348_cascade_\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_14\ : std_logic;
signal \ppm_encoder_1.init_pulses_18_i_0_14_cascade_\ : std_logic;
signal \ppm_encoder_1.init_pulses_18_i_a2_0_14\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_16\ : std_logic;
signal \ppm_encoder_1.N_241_cascade_\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_13\ : std_logic;
signal \ppm_encoder_1.pulses2count_9_0_o2_0_13_cascade_\ : std_logic;
signal scaler_2_data_13 : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_12_THRU_CO\ : std_logic;
signal \ppm_encoder_1.aileronZ0Z_13\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_0_13_cascade_\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_axb_13_cascade_\ : std_logic;
signal \ppm_encoder_1.init_pulses_RNIC11J5Z0Z_13\ : std_logic;
signal scaler_3_data_13 : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_12_THRU_CO\ : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_13\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_1_11\ : std_logic;
signal scaler_3_data_11 : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_10_THRU_CO\ : std_logic;
signal scaler_1_data_11 : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_10_THRU_CO\ : std_logic;
signal scaler_2_data_12 : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_11_THRU_CO\ : std_logic;
signal \ppm_encoder_1.N_418\ : std_logic;
signal \ppm_encoder_1.N_417_cascade_\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_1_8_cascade_\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_7_THRU_CO\ : std_logic;
signal scaler_2_data_8 : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_7_THRU_CO\ : std_logic;
signal scaler_1_data_8 : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_7_THRU_CO\ : std_logic;
signal scaler_3_data_8 : std_logic;
signal scaler_3_data_5 : std_logic;
signal scaler_4_data_4 : std_logic;
signal scaler_1_data_4 : std_logic;
signal scaler_1_data_5 : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_5\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_axb_5_1_sn_cascade_\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_axb_5_1_cascade_\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_axb_5_cascade_\ : std_logic;
signal \ppm_encoder_1.init_pulses_RNIT8FS5Z0Z_5\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_axb_5_1_rn_0\ : std_logic;
signal scaler_2_data_5 : std_logic;
signal \ppm_encoder_1.aileronZ0Z_5\ : std_logic;
signal scaler_4_data_5 : std_logic;
signal \ppm_encoder_1.scaler_1_dv_0\ : std_logic;
signal \ppm_encoder_1.N_252_i_i\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_axb_8\ : std_logic;
signal \ppm_encoder_1.init_pulses_RNITQDQ5Z0Z_8\ : std_logic;
signal \ppm_encoder_1.N_235_cascade_\ : std_logic;
signal \ppm_encoder_1.init_pulses_RNIUBDK6Z0Z_7\ : std_logic;
signal \ppm_encoder_1.N_114\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_1_12\ : std_logic;
signal \ppm_encoder_1.N_407_cascade_\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_axb_2_1_cascade_\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_axb_2_cascade_\ : std_logic;
signal \ppm_encoder_1.init_pulses_RNIE48O3Z0Z_2\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_0_14\ : std_logic;
signal \ppm_encoder_1.N_251_i_i\ : std_logic;
signal \ppm_encoder_1.aileronZ0Z_14\ : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_14\ : std_logic;
signal \ppm_encoder_1.pulses2count_9_i_o2_0_14\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_2_12\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_axb_12_cascade_\ : std_logic;
signal \ppm_encoder_1.init_pulses_RNI5FJB5Z0Z_12\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_6_cascade_\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_13\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_13\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_17\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_18\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_1\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_15\ : std_logic;
signal \ppm_encoder_1.N_245_i_i\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_9\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_10\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_11\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_12\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_2\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_3\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_5\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_6\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_7\ : std_logic;
signal \ppm_encoder_1.N_241\ : std_logic;
signal \ppm_encoder_1.N_348\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_8\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_7_THRU_CO\ : std_logic;
signal scaler_4_data_8 : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_6_THRU_CO\ : std_logic;
signal scaler_1_data_7 : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_6_THRU_CO\ : std_logic;
signal scaler_4_data_7 : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_sn_7_cascade_\ : std_logic;
signal \ppm_encoder_1.un2_throttle_0_0_7_cascade_\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_axb_7\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0\ : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_7\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_rn_0_7\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_6_THRU_CO\ : std_logic;
signal scaler_2_data_7 : std_logic;
signal \ppm_encoder_1.aileronZ0Z_7\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_axb_1_cascade_\ : std_logic;
signal \ppm_encoder_1.init_pulses_RNIOC8K3Z0Z_1\ : std_logic;
signal \ppm_encoder_1.N_426\ : std_logic;
signal \ppm_encoder_1.N_246\ : std_logic;
signal \ppm_encoder_1.N_426_cascade_\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_axb_3_cascade_\ : std_logic;
signal \ppm_encoder_1.init_pulses_RNISG8K3Z0Z_3\ : std_logic;
signal scaler_1_dv : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_1\ : std_logic;
signal \ppm_encoder_1.N_248_i_i\ : std_logic;
signal \ppm_encoder_1.N_250_i_i\ : std_logic;
signal \ppm_encoder_1.N_254_i_i\ : std_logic;
signal \ppm_encoder_1.PPM_STATE_fast_RNICIABZ0Z_0_cascade_\ : std_logic;
signal \ppm_encoder_1.N_246_i_i\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_1\ : std_logic;
signal \ppm_encoder_1.N_256_i_i\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_3_repZ0Z1\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_axb_16\ : std_logic;
signal \ppm_encoder_1.N_305\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIK17JZ0Z_3\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_2_cascade_\ : std_logic;
signal \ppm_encoder_1.N_260_i_i\ : std_logic;
signal \ppm_encoder_1.PPM_STATE_fast_RNI4RFRZ0Z_0_cascade_\ : std_logic;
signal \ppm_encoder_1.init_pulses_RNI83R42Z0Z_0\ : std_logic;
signal \bfn_9_26_0_\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_1\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_1\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_0\ : std_logic;
signal \ppm_encoder_1.init_pulses_RNIGLA33Z0Z_2\ : std_logic;
signal \ppm_encoder_1.N_249_i_i\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_2\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_1\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_3\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_3\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_2\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_4\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_4\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_3\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_5\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_5\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_4\ : std_logic;
signal \ppm_encoder_1.init_pulses_RNI69BV2Z0Z_6\ : std_logic;
signal \ppm_encoder_1.N_253_i_i\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_6\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_5\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_7\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_6\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_7\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_8\ : std_logic;
signal \bfn_9_27_0_\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_9\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_9\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_8\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_10\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_10\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_9\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_11\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_11\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_10\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_12\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_12\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_11\ : std_logic;
signal \ppm_encoder_1.N_259_i_i\ : std_logic;
signal \ppm_encoder_1.init_pulses_RNIKON03Z0Z_13\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_13\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_12\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_13_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_13\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_15\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_14\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_15\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_16\ : std_logic;
signal \bfn_9_28_0_\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_17\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_16\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_17\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_18\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_16\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_14\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_17\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_ns_2\ : std_logic;
signal \ppm_encoder_1.N_204_cascade_\ : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_8\ : std_logic;
signal \ppm_encoder_1.aileronZ0Z_8\ : std_logic;
signal \ppm_encoder_1.N_379_cascade_\ : std_logic;
signal \ppm_encoder_1.rudderZ0Z_8\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_7\ : std_logic;
signal \ppm_encoder_1.pulses2count_9_i_o2_0_7\ : std_logic;
signal \ppm_encoder_1.rudderZ0Z_12\ : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_11\ : std_logic;
signal \ppm_encoder_1.pulses2count_9_i_0_8\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_8\ : std_logic;
signal \ppm_encoder_1.rudderZ0Z_11\ : std_logic;
signal \ppm_encoder_1.N_391\ : std_logic;
signal \ppm_encoder_1.aileronZ0Z_12\ : std_logic;
signal \ppm_encoder_1.N_396\ : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_12\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_9\ : std_logic;
signal \ppm_encoder_1.N_325\ : std_logic;
signal \ppm_encoder_1.N_327_cascade_\ : std_logic;
signal \ppm_encoder_1.rudderZ0Z_9\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_5\ : std_logic;
signal \ppm_encoder_1.pulses2count_9_i_o2_0_5\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_8\ : std_logic;
signal \ppm_encoder_1.N_204\ : std_logic;
signal \ppm_encoder_1.N_255_i_i\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_12\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_12\ : std_logic;
signal \ppm_encoder_1.N_258_i_i\ : std_logic;
signal \ppm_encoder_1.N_257_i_i\ : std_logic;
signal \ppm_encoder_1.rudderZ0Z_6\ : std_logic;
signal \ppm_encoder_1.pulses2count_9_0_0_6\ : std_logic;
signal \ppm_encoder_1.N_301\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_6\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_6\ : std_logic;
signal \ppm_encoder_1.N_302\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_7\ : std_logic;
signal \ppm_encoder_1.pulses2count_9_0_2_12\ : std_logic;
signal \ppm_encoder_1.N_393\ : std_logic;
signal \ppm_encoder_1.pulses2count_9_0_0_12\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_3\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_3_repZ0Z2\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z1\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_7\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_7\ : std_logic;
signal \ppm_encoder_1.PPM_STATE_fastZ0Z_0\ : std_logic;
signal \ppm_encoder_1.aileronZ0Z_11\ : std_logic;
signal \ppm_encoder_1.init_pulses_RNILB4MZ0Z_0\ : std_logic;
signal \ppm_encoder_1.N_247_i_i\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z2\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z2\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z2\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_11\ : std_logic;
signal \ppm_encoder_1.N_441_cascade_\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_11\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_18\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_10\ : std_logic;
signal \ppm_encoder_1.rudderZ0Z_10\ : std_logic;
signal \ppm_encoder_1.N_383\ : std_logic;
signal \ppm_encoder_1.N_385_cascade_\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_4\ : std_logic;
signal \ppm_encoder_1.N_369\ : std_logic;
signal \ppm_encoder_1.N_371_cascade_\ : std_logic;
signal \ppm_encoder_1.rudderZ0Z_4\ : std_logic;
signal \ppm_encoder_1.rudderZ0Z_13\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_15\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_2\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_3\ : std_logic;
signal \ppm_encoder_1.N_360\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_2\ : std_logic;
signal \ppm_encoder_1.pulses2count_9_0_0_3\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_2\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_3\ : std_logic;
signal \ppm_encoder_1.N_365\ : std_logic;
signal \ppm_encoder_1.N_443\ : std_logic;
signal \ppm_encoder_1.pulses2count_9_0_2_1\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_1\ : std_logic;
signal \bfn_11_24_0_\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_0\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_2\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_1\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_3\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_2\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_3\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_4\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_5\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_6\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_7\ : std_logic;
signal \bfn_11_25_0_\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_8\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_9\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_10\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_11\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_12\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_13\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_14\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_15\ : std_logic;
signal \bfn_11_26_0_\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_16\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_17\ : std_logic;
signal \ppm_encoder_1.N_512_g\ : std_logic;
signal \ppm_encoder_1.N_247\ : std_logic;
signal \ppm_encoder_1.pulses2count_9_0_2_11\ : std_logic;
signal \ppm_encoder_1.N_388\ : std_logic;
signal \ppm_encoder_1.pulses2count_9_0_0_11\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_13\ : std_logic;
signal \ppm_encoder_1.pulses2count_9_0_0_13\ : std_logic;
signal \ppm_encoder_1.N_303\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_16\ : std_logic;
signal \ppm_encoder_1.PPM_STATE_fast_RNICIABZ0Z_0\ : std_logic;
signal \ppm_encoder_1.N_238_i_0\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_17\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_18\ : std_logic;
signal \ppm_encoder_1.rudderZ0Z_5\ : std_logic;
signal \ppm_encoder_1.rudderZ0Z_7\ : std_logic;
signal \ppm_encoder_1.pulses2count_9_i_0_7\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_0\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_1\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_1\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_0\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNELZ0Z_1\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNELZ0Z_0\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_15\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNELZ0Z_3\ : std_logic;
signal \ppm_encoder_1.N_235\ : std_logic;
signal \ppm_encoder_1.rudderZ0Z_14\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_14\ : std_logic;
signal \ppm_encoder_1.pulses2count_9_i_0_14_cascade_\ : std_logic;
signal \ppm_encoder_1.N_304\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_4\ : std_logic;
signal \ppm_encoder_1.pulses2count_9_i_1_4\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_4\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_4\ : std_logic;
signal \ppm_encoder_1.N_300\ : std_logic;
signal \ppm_encoder_1.pulses2count_9_i_0_5\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_5\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_5\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_10\ : std_logic;
signal \ppm_encoder_1.pulses2count_9_i_1_10\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_10\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_11\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_11\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_10\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_14\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_15\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_7\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_5\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_14\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_6\ : std_logic;
signal \ppm_encoder_1.un1_PPM_STATE_0_sqmuxa_0_i_0_a2_1\ : std_logic;
signal \ppm_encoder_1.un1_PPM_STATE_0_sqmuxa_0_i_0_a2_16_4_cascade_\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_12\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_13\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_12\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_18\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_18\ : std_logic;
signal \ppm_encoder_1.un1_PPM_STATE_0_sqmuxa_0_i_0_a2_2_3\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_15\ : std_logic;
signal \ppm_encoder_1.un1_PPM_STATE_0_sqmuxa_0_i_0_a2_2_4\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_13\ : std_logic;
signal \ppm_encoder_1.un1_PPM_STATE_0_sqmuxa_0_i_0_a2_2\ : std_logic;
signal \ppm_encoder_1.un1_PPM_STATE_1_sqmuxa_i_i_a2_0_1\ : std_logic;
signal \ppm_encoder_1.un1_PPM_STATE_0_sqmuxa_0_i_0_a2_16_4\ : std_logic;
signal \ppm_encoder_1.un1_PPM_STATE_0_sqmuxa_0_i_0_a2_2_cascade_\ : std_logic;
signal \ppm_encoder_1.un1_PPM_STATE_0_sqmuxa_0_i_0_a2_16_5\ : std_logic;
signal \ppm_encoder_1.counter24_0_I_57_c_RNIJMMDZ0\ : std_logic;
signal \ppm_encoder_1.N_431_cascade_\ : std_logic;
signal \ppm_encoder_1.PPM_STATEZ0Z_1\ : std_logic;
signal ppm_output_c : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_16\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_17\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_17\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_16\ : std_logic;
signal \ppm_encoder_1.pulses2count_9_i_1_8\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_8\ : std_logic;
signal \ppm_encoder_1.pulses2count_9_i_0_1_9\ : std_logic;
signal \ppm_encoder_1.N_441\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_9\ : std_logic;
signal \ppm_encoder_1.N_244\ : std_logic;
signal \ppm_encoder_1.pulses2count_9_0_1_0\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNELZ0Z_2\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_0\ : std_logic;
signal clk_system_c_g : std_logic;
signal \ppm_encoder_1.N_238_i_0_g\ : std_logic;
signal reset_system_g : std_logic;
signal \ppm_encoder_1.counter24_0_I_1_c_RNOZ0\ : std_logic;
signal \bfn_13_24_0_\ : std_logic;
signal \ppm_encoder_1.counter24_0_I_9_c_RNOZ0\ : std_logic;
signal \ppm_encoder_1.counter24_0_data_tmp_0\ : std_logic;
signal \ppm_encoder_1.counter24_0_I_15_c_RNOZ0\ : std_logic;
signal \ppm_encoder_1.counter24_0_data_tmp_1\ : std_logic;
signal \ppm_encoder_1.counter24_0_I_21_c_RNOZ0\ : std_logic;
signal \ppm_encoder_1.counter24_0_data_tmp_2\ : std_logic;
signal \ppm_encoder_1.counter24_0_data_tmp_3\ : std_logic;
signal \ppm_encoder_1.counter24_0_I_33_c_RNOZ0\ : std_logic;
signal \ppm_encoder_1.counter24_0_data_tmp_4\ : std_logic;
signal \ppm_encoder_1.counter24_0_I_39_c_RNOZ0\ : std_logic;
signal \ppm_encoder_1.counter24_0_data_tmp_5\ : std_logic;
signal \ppm_encoder_1.counter24_0_I_45_c_RNOZ0\ : std_logic;
signal \ppm_encoder_1.counter24_0_data_tmp_6\ : std_logic;
signal \ppm_encoder_1.counter24_0_data_tmp_7\ : std_logic;
signal \ppm_encoder_1.counter24_0_I_51_c_RNOZ0\ : std_logic;
signal \bfn_13_25_0_\ : std_logic;
signal \ppm_encoder_1.counter24_0_I_57_c_RNOZ0\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \ppm_encoder_1.counter24_0_data_tmp_8\ : std_logic;
signal \ppm_encoder_1.counter24_0_N_2\ : std_logic;
signal \ppm_encoder_1.N_330\ : std_logic;
signal \ppm_encoder_1.counter24_0_N_2_THRU_CO\ : std_logic;
signal reset_system : std_logic;
signal \ppm_encoder_1.PPM_STATEZ0Z_0\ : std_logic;
signal \ppm_encoder_1.counter24_0_I_57_c_RNIGCOZ0Z83\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_9\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_8\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_9\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_8\ : std_logic;
signal \ppm_encoder_1.counter24_0_I_27_c_RNOZ0\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal clk_system_wire : std_logic;
signal ppm_output_wire : std_logic;
signal frame_decoder_dv_wire : std_logic;
signal uart_input_wire : std_logic;
signal uart_input_debug_wire : std_logic;

begin
    clk_system_wire <= clk_system;
    ppm_output <= ppm_output_wire;
    frame_decoder_dv <= frame_decoder_dv_wire;
    uart_input_wire <= uart_input;
    uart_input_debug <= uart_input_debug_wire;

    \clk_system_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__24856\,
            GLOBALBUFFEROUTPUT => clk_system_c_g
        );

    \clk_system_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24858\,
            DIN => \N__24857\,
            DOUT => \N__24856\,
            PACKAGEPIN => clk_system_wire
        );

    \clk_system_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__24858\,
            PADOUT => \N__24857\,
            PADIN => \N__24856\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ppm_output_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24847\,
            DIN => \N__24846\,
            DOUT => \N__24845\,
            PACKAGEPIN => ppm_output_wire
        );

    \ppm_output_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__24847\,
            PADOUT => \N__24846\,
            PADIN => \N__24845\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__22803\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \frame_decoder_dv_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24838\,
            DIN => \N__24837\,
            DOUT => \N__24836\,
            PACKAGEPIN => frame_decoder_dv_wire
        );

    \frame_decoder_dv_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__24838\,
            PADOUT => \N__24837\,
            PADIN => \N__24836\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__14955\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \uart_input_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24829\,
            DIN => \N__24828\,
            DOUT => \N__24827\,
            PACKAGEPIN => uart_input_wire
        );

    \uart_input_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__24829\,
            PADOUT => \N__24828\,
            PADIN => \N__24827\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => uart_input_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \uart_input_debug_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24820\,
            DIN => \N__24819\,
            DOUT => \N__24818\,
            PACKAGEPIN => uart_input_debug_wire
        );

    \uart_input_debug_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__24820\,
            PADOUT => \N__24819\,
            PADIN => \N__24818\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__15410\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__5994\ : InMux
    port map (
            O => \N__24801\,
            I => \N__24798\
        );

    \I__5993\ : LocalMux
    port map (
            O => \N__24798\,
            I => \ppm_encoder_1.counter24_0_I_39_c_RNOZ0\
        );

    \I__5992\ : InMux
    port map (
            O => \N__24795\,
            I => \N__24792\
        );

    \I__5991\ : LocalMux
    port map (
            O => \N__24792\,
            I => \ppm_encoder_1.counter24_0_I_45_c_RNOZ0\
        );

    \I__5990\ : CascadeMux
    port map (
            O => \N__24789\,
            I => \N__24786\
        );

    \I__5989\ : InMux
    port map (
            O => \N__24786\,
            I => \N__24783\
        );

    \I__5988\ : LocalMux
    port map (
            O => \N__24783\,
            I => \N__24780\
        );

    \I__5987\ : Odrv4
    port map (
            O => \N__24780\,
            I => \ppm_encoder_1.counter24_0_I_51_c_RNOZ0\
        );

    \I__5986\ : InMux
    port map (
            O => \N__24777\,
            I => \N__24774\
        );

    \I__5985\ : LocalMux
    port map (
            O => \N__24774\,
            I => \ppm_encoder_1.counter24_0_I_57_c_RNOZ0\
        );

    \I__5984\ : CascadeMux
    port map (
            O => \N__24771\,
            I => \N__24764\
        );

    \I__5983\ : CascadeMux
    port map (
            O => \N__24770\,
            I => \N__24761\
        );

    \I__5982\ : CascadeMux
    port map (
            O => \N__24769\,
            I => \N__24758\
        );

    \I__5981\ : CascadeMux
    port map (
            O => \N__24768\,
            I => \N__24754\
        );

    \I__5980\ : CascadeMux
    port map (
            O => \N__24767\,
            I => \N__24751\
        );

    \I__5979\ : InMux
    port map (
            O => \N__24764\,
            I => \N__24738\
        );

    \I__5978\ : InMux
    port map (
            O => \N__24761\,
            I => \N__24735\
        );

    \I__5977\ : InMux
    port map (
            O => \N__24758\,
            I => \N__24732\
        );

    \I__5976\ : CascadeMux
    port map (
            O => \N__24757\,
            I => \N__24729\
        );

    \I__5975\ : InMux
    port map (
            O => \N__24754\,
            I => \N__24726\
        );

    \I__5974\ : InMux
    port map (
            O => \N__24751\,
            I => \N__24723\
        );

    \I__5973\ : CascadeMux
    port map (
            O => \N__24750\,
            I => \N__24720\
        );

    \I__5972\ : CascadeMux
    port map (
            O => \N__24749\,
            I => \N__24717\
        );

    \I__5971\ : CascadeMux
    port map (
            O => \N__24748\,
            I => \N__24713\
        );

    \I__5970\ : CascadeMux
    port map (
            O => \N__24747\,
            I => \N__24709\
        );

    \I__5969\ : CascadeMux
    port map (
            O => \N__24746\,
            I => \N__24706\
        );

    \I__5968\ : CascadeMux
    port map (
            O => \N__24745\,
            I => \N__24703\
        );

    \I__5967\ : CascadeMux
    port map (
            O => \N__24744\,
            I => \N__24700\
        );

    \I__5966\ : CascadeMux
    port map (
            O => \N__24743\,
            I => \N__24697\
        );

    \I__5965\ : CascadeMux
    port map (
            O => \N__24742\,
            I => \N__24694\
        );

    \I__5964\ : CascadeMux
    port map (
            O => \N__24741\,
            I => \N__24691\
        );

    \I__5963\ : LocalMux
    port map (
            O => \N__24738\,
            I => \N__24687\
        );

    \I__5962\ : LocalMux
    port map (
            O => \N__24735\,
            I => \N__24682\
        );

    \I__5961\ : LocalMux
    port map (
            O => \N__24732\,
            I => \N__24682\
        );

    \I__5960\ : InMux
    port map (
            O => \N__24729\,
            I => \N__24679\
        );

    \I__5959\ : LocalMux
    port map (
            O => \N__24726\,
            I => \N__24674\
        );

    \I__5958\ : LocalMux
    port map (
            O => \N__24723\,
            I => \N__24674\
        );

    \I__5957\ : InMux
    port map (
            O => \N__24720\,
            I => \N__24671\
        );

    \I__5956\ : InMux
    port map (
            O => \N__24717\,
            I => \N__24668\
        );

    \I__5955\ : InMux
    port map (
            O => \N__24716\,
            I => \N__24665\
        );

    \I__5954\ : InMux
    port map (
            O => \N__24713\,
            I => \N__24660\
        );

    \I__5953\ : InMux
    port map (
            O => \N__24712\,
            I => \N__24660\
        );

    \I__5952\ : InMux
    port map (
            O => \N__24709\,
            I => \N__24651\
        );

    \I__5951\ : InMux
    port map (
            O => \N__24706\,
            I => \N__24651\
        );

    \I__5950\ : InMux
    port map (
            O => \N__24703\,
            I => \N__24651\
        );

    \I__5949\ : InMux
    port map (
            O => \N__24700\,
            I => \N__24651\
        );

    \I__5948\ : InMux
    port map (
            O => \N__24697\,
            I => \N__24644\
        );

    \I__5947\ : InMux
    port map (
            O => \N__24694\,
            I => \N__24644\
        );

    \I__5946\ : InMux
    port map (
            O => \N__24691\,
            I => \N__24644\
        );

    \I__5945\ : CascadeMux
    port map (
            O => \N__24690\,
            I => \N__24641\
        );

    \I__5944\ : Span4Mux_h
    port map (
            O => \N__24687\,
            I => \N__24634\
        );

    \I__5943\ : Span4Mux_v
    port map (
            O => \N__24682\,
            I => \N__24634\
        );

    \I__5942\ : LocalMux
    port map (
            O => \N__24679\,
            I => \N__24634\
        );

    \I__5941\ : Span4Mux_v
    port map (
            O => \N__24674\,
            I => \N__24629\
        );

    \I__5940\ : LocalMux
    port map (
            O => \N__24671\,
            I => \N__24629\
        );

    \I__5939\ : LocalMux
    port map (
            O => \N__24668\,
            I => \N__24624\
        );

    \I__5938\ : LocalMux
    port map (
            O => \N__24665\,
            I => \N__24624\
        );

    \I__5937\ : LocalMux
    port map (
            O => \N__24660\,
            I => \N__24617\
        );

    \I__5936\ : LocalMux
    port map (
            O => \N__24651\,
            I => \N__24617\
        );

    \I__5935\ : LocalMux
    port map (
            O => \N__24644\,
            I => \N__24617\
        );

    \I__5934\ : InMux
    port map (
            O => \N__24641\,
            I => \N__24614\
        );

    \I__5933\ : Span4Mux_v
    port map (
            O => \N__24634\,
            I => \N__24611\
        );

    \I__5932\ : Sp12to4
    port map (
            O => \N__24629\,
            I => \N__24608\
        );

    \I__5931\ : Span4Mux_v
    port map (
            O => \N__24624\,
            I => \N__24605\
        );

    \I__5930\ : Sp12to4
    port map (
            O => \N__24617\,
            I => \N__24602\
        );

    \I__5929\ : LocalMux
    port map (
            O => \N__24614\,
            I => \N__24599\
        );

    \I__5928\ : Span4Mux_h
    port map (
            O => \N__24611\,
            I => \N__24596\
        );

    \I__5927\ : Span12Mux_s11_v
    port map (
            O => \N__24608\,
            I => \N__24587\
        );

    \I__5926\ : Sp12to4
    port map (
            O => \N__24605\,
            I => \N__24587\
        );

    \I__5925\ : Span12Mux_s11_v
    port map (
            O => \N__24602\,
            I => \N__24587\
        );

    \I__5924\ : Span12Mux_s2_h
    port map (
            O => \N__24599\,
            I => \N__24587\
        );

    \I__5923\ : Odrv4
    port map (
            O => \N__24596\,
            I => \CONSTANT_ONE_NET\
        );

    \I__5922\ : Odrv12
    port map (
            O => \N__24587\,
            I => \CONSTANT_ONE_NET\
        );

    \I__5921\ : InMux
    port map (
            O => \N__24582\,
            I => \ppm_encoder_1.counter24_0_N_2\
        );

    \I__5920\ : InMux
    port map (
            O => \N__24579\,
            I => \N__24570\
        );

    \I__5919\ : InMux
    port map (
            O => \N__24578\,
            I => \N__24570\
        );

    \I__5918\ : InMux
    port map (
            O => \N__24577\,
            I => \N__24570\
        );

    \I__5917\ : LocalMux
    port map (
            O => \N__24570\,
            I => \N__24566\
        );

    \I__5916\ : InMux
    port map (
            O => \N__24569\,
            I => \N__24563\
        );

    \I__5915\ : Odrv4
    port map (
            O => \N__24566\,
            I => \ppm_encoder_1.N_330\
        );

    \I__5914\ : LocalMux
    port map (
            O => \N__24563\,
            I => \ppm_encoder_1.N_330\
        );

    \I__5913\ : InMux
    port map (
            O => \N__24558\,
            I => \N__24555\
        );

    \I__5912\ : LocalMux
    port map (
            O => \N__24555\,
            I => \N__24551\
        );

    \I__5911\ : InMux
    port map (
            O => \N__24554\,
            I => \N__24547\
        );

    \I__5910\ : Span12Mux_s5_v
    port map (
            O => \N__24551\,
            I => \N__24544\
        );

    \I__5909\ : InMux
    port map (
            O => \N__24550\,
            I => \N__24541\
        );

    \I__5908\ : LocalMux
    port map (
            O => \N__24547\,
            I => \ppm_encoder_1.counter24_0_N_2_THRU_CO\
        );

    \I__5907\ : Odrv12
    port map (
            O => \N__24544\,
            I => \ppm_encoder_1.counter24_0_N_2_THRU_CO\
        );

    \I__5906\ : LocalMux
    port map (
            O => \N__24541\,
            I => \ppm_encoder_1.counter24_0_N_2_THRU_CO\
        );

    \I__5905\ : CascadeMux
    port map (
            O => \N__24534\,
            I => \N__24530\
        );

    \I__5904\ : CascadeMux
    port map (
            O => \N__24533\,
            I => \N__24525\
        );

    \I__5903\ : InMux
    port map (
            O => \N__24530\,
            I => \N__24517\
        );

    \I__5902\ : InMux
    port map (
            O => \N__24529\,
            I => \N__24517\
        );

    \I__5901\ : InMux
    port map (
            O => \N__24528\,
            I => \N__24517\
        );

    \I__5900\ : InMux
    port map (
            O => \N__24525\,
            I => \N__24514\
        );

    \I__5899\ : IoInMux
    port map (
            O => \N__24524\,
            I => \N__24511\
        );

    \I__5898\ : LocalMux
    port map (
            O => \N__24517\,
            I => \N__24508\
        );

    \I__5897\ : LocalMux
    port map (
            O => \N__24514\,
            I => \N__24504\
        );

    \I__5896\ : LocalMux
    port map (
            O => \N__24511\,
            I => \N__24501\
        );

    \I__5895\ : Span4Mux_h
    port map (
            O => \N__24508\,
            I => \N__24497\
        );

    \I__5894\ : InMux
    port map (
            O => \N__24507\,
            I => \N__24494\
        );

    \I__5893\ : Span4Mux_v
    port map (
            O => \N__24504\,
            I => \N__24491\
        );

    \I__5892\ : IoSpan4Mux
    port map (
            O => \N__24501\,
            I => \N__24488\
        );

    \I__5891\ : InMux
    port map (
            O => \N__24500\,
            I => \N__24483\
        );

    \I__5890\ : Span4Mux_h
    port map (
            O => \N__24497\,
            I => \N__24480\
        );

    \I__5889\ : LocalMux
    port map (
            O => \N__24494\,
            I => \N__24477\
        );

    \I__5888\ : Span4Mux_h
    port map (
            O => \N__24491\,
            I => \N__24474\
        );

    \I__5887\ : Span4Mux_s3_v
    port map (
            O => \N__24488\,
            I => \N__24471\
        );

    \I__5886\ : InMux
    port map (
            O => \N__24487\,
            I => \N__24468\
        );

    \I__5885\ : InMux
    port map (
            O => \N__24486\,
            I => \N__24464\
        );

    \I__5884\ : LocalMux
    port map (
            O => \N__24483\,
            I => \N__24457\
        );

    \I__5883\ : Span4Mux_v
    port map (
            O => \N__24480\,
            I => \N__24457\
        );

    \I__5882\ : Span4Mux_h
    port map (
            O => \N__24477\,
            I => \N__24452\
        );

    \I__5881\ : Span4Mux_h
    port map (
            O => \N__24474\,
            I => \N__24452\
        );

    \I__5880\ : Span4Mux_v
    port map (
            O => \N__24471\,
            I => \N__24449\
        );

    \I__5879\ : LocalMux
    port map (
            O => \N__24468\,
            I => \N__24446\
        );

    \I__5878\ : InMux
    port map (
            O => \N__24467\,
            I => \N__24443\
        );

    \I__5877\ : LocalMux
    port map (
            O => \N__24464\,
            I => \N__24440\
        );

    \I__5876\ : InMux
    port map (
            O => \N__24463\,
            I => \N__24435\
        );

    \I__5875\ : InMux
    port map (
            O => \N__24462\,
            I => \N__24435\
        );

    \I__5874\ : Span4Mux_v
    port map (
            O => \N__24457\,
            I => \N__24432\
        );

    \I__5873\ : Span4Mux_v
    port map (
            O => \N__24452\,
            I => \N__24429\
        );

    \I__5872\ : Span4Mux_v
    port map (
            O => \N__24449\,
            I => \N__24426\
        );

    \I__5871\ : Odrv12
    port map (
            O => \N__24446\,
            I => reset_system
        );

    \I__5870\ : LocalMux
    port map (
            O => \N__24443\,
            I => reset_system
        );

    \I__5869\ : Odrv4
    port map (
            O => \N__24440\,
            I => reset_system
        );

    \I__5868\ : LocalMux
    port map (
            O => \N__24435\,
            I => reset_system
        );

    \I__5867\ : Odrv4
    port map (
            O => \N__24432\,
            I => reset_system
        );

    \I__5866\ : Odrv4
    port map (
            O => \N__24429\,
            I => reset_system
        );

    \I__5865\ : Odrv4
    port map (
            O => \N__24426\,
            I => reset_system
        );

    \I__5864\ : InMux
    port map (
            O => \N__24411\,
            I => \N__24408\
        );

    \I__5863\ : LocalMux
    port map (
            O => \N__24408\,
            I => \N__24402\
        );

    \I__5862\ : InMux
    port map (
            O => \N__24407\,
            I => \N__24398\
        );

    \I__5861\ : InMux
    port map (
            O => \N__24406\,
            I => \N__24395\
        );

    \I__5860\ : CascadeMux
    port map (
            O => \N__24405\,
            I => \N__24390\
        );

    \I__5859\ : Span4Mux_h
    port map (
            O => \N__24402\,
            I => \N__24387\
        );

    \I__5858\ : InMux
    port map (
            O => \N__24401\,
            I => \N__24384\
        );

    \I__5857\ : LocalMux
    port map (
            O => \N__24398\,
            I => \N__24379\
        );

    \I__5856\ : LocalMux
    port map (
            O => \N__24395\,
            I => \N__24379\
        );

    \I__5855\ : InMux
    port map (
            O => \N__24394\,
            I => \N__24374\
        );

    \I__5854\ : InMux
    port map (
            O => \N__24393\,
            I => \N__24374\
        );

    \I__5853\ : InMux
    port map (
            O => \N__24390\,
            I => \N__24371\
        );

    \I__5852\ : Odrv4
    port map (
            O => \N__24387\,
            I => \ppm_encoder_1.PPM_STATEZ0Z_0\
        );

    \I__5851\ : LocalMux
    port map (
            O => \N__24384\,
            I => \ppm_encoder_1.PPM_STATEZ0Z_0\
        );

    \I__5850\ : Odrv4
    port map (
            O => \N__24379\,
            I => \ppm_encoder_1.PPM_STATEZ0Z_0\
        );

    \I__5849\ : LocalMux
    port map (
            O => \N__24374\,
            I => \ppm_encoder_1.PPM_STATEZ0Z_0\
        );

    \I__5848\ : LocalMux
    port map (
            O => \N__24371\,
            I => \ppm_encoder_1.PPM_STATEZ0Z_0\
        );

    \I__5847\ : IoInMux
    port map (
            O => \N__24360\,
            I => \N__24357\
        );

    \I__5846\ : LocalMux
    port map (
            O => \N__24357\,
            I => \N__24354\
        );

    \I__5845\ : Span12Mux_s5_v
    port map (
            O => \N__24354\,
            I => \N__24351\
        );

    \I__5844\ : Odrv12
    port map (
            O => \N__24351\,
            I => \ppm_encoder_1.counter24_0_I_57_c_RNIGCOZ0Z83\
        );

    \I__5843\ : InMux
    port map (
            O => \N__24348\,
            I => \N__24342\
        );

    \I__5842\ : InMux
    port map (
            O => \N__24347\,
            I => \N__24339\
        );

    \I__5841\ : InMux
    port map (
            O => \N__24346\,
            I => \N__24336\
        );

    \I__5840\ : InMux
    port map (
            O => \N__24345\,
            I => \N__24333\
        );

    \I__5839\ : LocalMux
    port map (
            O => \N__24342\,
            I => \N__24330\
        );

    \I__5838\ : LocalMux
    port map (
            O => \N__24339\,
            I => \ppm_encoder_1.counterZ0Z_9\
        );

    \I__5837\ : LocalMux
    port map (
            O => \N__24336\,
            I => \ppm_encoder_1.counterZ0Z_9\
        );

    \I__5836\ : LocalMux
    port map (
            O => \N__24333\,
            I => \ppm_encoder_1.counterZ0Z_9\
        );

    \I__5835\ : Odrv12
    port map (
            O => \N__24330\,
            I => \ppm_encoder_1.counterZ0Z_9\
        );

    \I__5834\ : InMux
    port map (
            O => \N__24321\,
            I => \N__24318\
        );

    \I__5833\ : LocalMux
    port map (
            O => \N__24318\,
            I => \N__24315\
        );

    \I__5832\ : Odrv12
    port map (
            O => \N__24315\,
            I => \ppm_encoder_1.pulses2countZ0Z_8\
        );

    \I__5831\ : CascadeMux
    port map (
            O => \N__24312\,
            I => \N__24309\
        );

    \I__5830\ : InMux
    port map (
            O => \N__24309\,
            I => \N__24306\
        );

    \I__5829\ : LocalMux
    port map (
            O => \N__24306\,
            I => \N__24303\
        );

    \I__5828\ : Odrv4
    port map (
            O => \N__24303\,
            I => \ppm_encoder_1.pulses2countZ0Z_9\
        );

    \I__5827\ : InMux
    port map (
            O => \N__24300\,
            I => \N__24295\
        );

    \I__5826\ : InMux
    port map (
            O => \N__24299\,
            I => \N__24292\
        );

    \I__5825\ : InMux
    port map (
            O => \N__24298\,
            I => \N__24289\
        );

    \I__5824\ : LocalMux
    port map (
            O => \N__24295\,
            I => \N__24286\
        );

    \I__5823\ : LocalMux
    port map (
            O => \N__24292\,
            I => \ppm_encoder_1.counterZ0Z_8\
        );

    \I__5822\ : LocalMux
    port map (
            O => \N__24289\,
            I => \ppm_encoder_1.counterZ0Z_8\
        );

    \I__5821\ : Odrv4
    port map (
            O => \N__24286\,
            I => \ppm_encoder_1.counterZ0Z_8\
        );

    \I__5820\ : InMux
    port map (
            O => \N__24279\,
            I => \N__24276\
        );

    \I__5819\ : LocalMux
    port map (
            O => \N__24276\,
            I => \ppm_encoder_1.counter24_0_I_27_c_RNOZ0\
        );

    \I__5818\ : InMux
    port map (
            O => \N__24273\,
            I => \N__24270\
        );

    \I__5817\ : LocalMux
    port map (
            O => \N__24270\,
            I => \N__24267\
        );

    \I__5816\ : Span4Mux_v
    port map (
            O => \N__24267\,
            I => \N__24264\
        );

    \I__5815\ : Odrv4
    port map (
            O => \N__24264\,
            I => \ppm_encoder_1.pulses2count_9_i_0_1_9\
        );

    \I__5814\ : InMux
    port map (
            O => \N__24261\,
            I => \N__24250\
        );

    \I__5813\ : InMux
    port map (
            O => \N__24260\,
            I => \N__24247\
        );

    \I__5812\ : InMux
    port map (
            O => \N__24259\,
            I => \N__24240\
        );

    \I__5811\ : InMux
    port map (
            O => \N__24258\,
            I => \N__24240\
        );

    \I__5810\ : InMux
    port map (
            O => \N__24257\,
            I => \N__24240\
        );

    \I__5809\ : InMux
    port map (
            O => \N__24256\,
            I => \N__24237\
        );

    \I__5808\ : InMux
    port map (
            O => \N__24255\,
            I => \N__24232\
        );

    \I__5807\ : InMux
    port map (
            O => \N__24254\,
            I => \N__24229\
        );

    \I__5806\ : CascadeMux
    port map (
            O => \N__24253\,
            I => \N__24226\
        );

    \I__5805\ : LocalMux
    port map (
            O => \N__24250\,
            I => \N__24222\
        );

    \I__5804\ : LocalMux
    port map (
            O => \N__24247\,
            I => \N__24219\
        );

    \I__5803\ : LocalMux
    port map (
            O => \N__24240\,
            I => \N__24216\
        );

    \I__5802\ : LocalMux
    port map (
            O => \N__24237\,
            I => \N__24213\
        );

    \I__5801\ : InMux
    port map (
            O => \N__24236\,
            I => \N__24208\
        );

    \I__5800\ : InMux
    port map (
            O => \N__24235\,
            I => \N__24208\
        );

    \I__5799\ : LocalMux
    port map (
            O => \N__24232\,
            I => \N__24203\
        );

    \I__5798\ : LocalMux
    port map (
            O => \N__24229\,
            I => \N__24203\
        );

    \I__5797\ : InMux
    port map (
            O => \N__24226\,
            I => \N__24200\
        );

    \I__5796\ : InMux
    port map (
            O => \N__24225\,
            I => \N__24197\
        );

    \I__5795\ : Span4Mux_v
    port map (
            O => \N__24222\,
            I => \N__24194\
        );

    \I__5794\ : Span4Mux_v
    port map (
            O => \N__24219\,
            I => \N__24191\
        );

    \I__5793\ : Span4Mux_h
    port map (
            O => \N__24216\,
            I => \N__24188\
        );

    \I__5792\ : Span12Mux_v
    port map (
            O => \N__24213\,
            I => \N__24185\
        );

    \I__5791\ : LocalMux
    port map (
            O => \N__24208\,
            I => \N__24178\
        );

    \I__5790\ : Span4Mux_h
    port map (
            O => \N__24203\,
            I => \N__24178\
        );

    \I__5789\ : LocalMux
    port map (
            O => \N__24200\,
            I => \N__24178\
        );

    \I__5788\ : LocalMux
    port map (
            O => \N__24197\,
            I => \ppm_encoder_1.N_441\
        );

    \I__5787\ : Odrv4
    port map (
            O => \N__24194\,
            I => \ppm_encoder_1.N_441\
        );

    \I__5786\ : Odrv4
    port map (
            O => \N__24191\,
            I => \ppm_encoder_1.N_441\
        );

    \I__5785\ : Odrv4
    port map (
            O => \N__24188\,
            I => \ppm_encoder_1.N_441\
        );

    \I__5784\ : Odrv12
    port map (
            O => \N__24185\,
            I => \ppm_encoder_1.N_441\
        );

    \I__5783\ : Odrv4
    port map (
            O => \N__24178\,
            I => \ppm_encoder_1.N_441\
        );

    \I__5782\ : CascadeMux
    port map (
            O => \N__24165\,
            I => \N__24162\
        );

    \I__5781\ : InMux
    port map (
            O => \N__24162\,
            I => \N__24158\
        );

    \I__5780\ : InMux
    port map (
            O => \N__24161\,
            I => \N__24154\
        );

    \I__5779\ : LocalMux
    port map (
            O => \N__24158\,
            I => \N__24151\
        );

    \I__5778\ : InMux
    port map (
            O => \N__24157\,
            I => \N__24148\
        );

    \I__5777\ : LocalMux
    port map (
            O => \N__24154\,
            I => \N__24144\
        );

    \I__5776\ : Span4Mux_h
    port map (
            O => \N__24151\,
            I => \N__24139\
        );

    \I__5775\ : LocalMux
    port map (
            O => \N__24148\,
            I => \N__24139\
        );

    \I__5774\ : InMux
    port map (
            O => \N__24147\,
            I => \N__24136\
        );

    \I__5773\ : Span4Mux_v
    port map (
            O => \N__24144\,
            I => \N__24131\
        );

    \I__5772\ : Span4Mux_v
    port map (
            O => \N__24139\,
            I => \N__24131\
        );

    \I__5771\ : LocalMux
    port map (
            O => \N__24136\,
            I => \ppm_encoder_1.init_pulsesZ0Z_9\
        );

    \I__5770\ : Odrv4
    port map (
            O => \N__24131\,
            I => \ppm_encoder_1.init_pulsesZ0Z_9\
        );

    \I__5769\ : CascadeMux
    port map (
            O => \N__24126\,
            I => \N__24122\
        );

    \I__5768\ : CascadeMux
    port map (
            O => \N__24125\,
            I => \N__24119\
        );

    \I__5767\ : InMux
    port map (
            O => \N__24122\,
            I => \N__24113\
        );

    \I__5766\ : InMux
    port map (
            O => \N__24119\,
            I => \N__24108\
        );

    \I__5765\ : InMux
    port map (
            O => \N__24118\,
            I => \N__24108\
        );

    \I__5764\ : InMux
    port map (
            O => \N__24117\,
            I => \N__24103\
        );

    \I__5763\ : InMux
    port map (
            O => \N__24116\,
            I => \N__24103\
        );

    \I__5762\ : LocalMux
    port map (
            O => \N__24113\,
            I => \ppm_encoder_1.N_244\
        );

    \I__5761\ : LocalMux
    port map (
            O => \N__24108\,
            I => \ppm_encoder_1.N_244\
        );

    \I__5760\ : LocalMux
    port map (
            O => \N__24103\,
            I => \ppm_encoder_1.N_244\
        );

    \I__5759\ : InMux
    port map (
            O => \N__24096\,
            I => \N__24093\
        );

    \I__5758\ : LocalMux
    port map (
            O => \N__24093\,
            I => \ppm_encoder_1.pulses2count_9_0_1_0\
        );

    \I__5757\ : CascadeMux
    port map (
            O => \N__24090\,
            I => \N__24082\
        );

    \I__5756\ : CascadeMux
    port map (
            O => \N__24089\,
            I => \N__24079\
        );

    \I__5755\ : CascadeMux
    port map (
            O => \N__24088\,
            I => \N__24074\
        );

    \I__5754\ : CascadeMux
    port map (
            O => \N__24087\,
            I => \N__24070\
        );

    \I__5753\ : CascadeMux
    port map (
            O => \N__24086\,
            I => \N__24063\
        );

    \I__5752\ : CascadeMux
    port map (
            O => \N__24085\,
            I => \N__24060\
        );

    \I__5751\ : InMux
    port map (
            O => \N__24082\,
            I => \N__24057\
        );

    \I__5750\ : InMux
    port map (
            O => \N__24079\,
            I => \N__24053\
        );

    \I__5749\ : InMux
    port map (
            O => \N__24078\,
            I => \N__24050\
        );

    \I__5748\ : InMux
    port map (
            O => \N__24077\,
            I => \N__24041\
        );

    \I__5747\ : InMux
    port map (
            O => \N__24074\,
            I => \N__24041\
        );

    \I__5746\ : InMux
    port map (
            O => \N__24073\,
            I => \N__24041\
        );

    \I__5745\ : InMux
    port map (
            O => \N__24070\,
            I => \N__24041\
        );

    \I__5744\ : InMux
    port map (
            O => \N__24069\,
            I => \N__24032\
        );

    \I__5743\ : InMux
    port map (
            O => \N__24068\,
            I => \N__24032\
        );

    \I__5742\ : InMux
    port map (
            O => \N__24067\,
            I => \N__24032\
        );

    \I__5741\ : InMux
    port map (
            O => \N__24066\,
            I => \N__24032\
        );

    \I__5740\ : InMux
    port map (
            O => \N__24063\,
            I => \N__24029\
        );

    \I__5739\ : InMux
    port map (
            O => \N__24060\,
            I => \N__24026\
        );

    \I__5738\ : LocalMux
    port map (
            O => \N__24057\,
            I => \N__24021\
        );

    \I__5737\ : InMux
    port map (
            O => \N__24056\,
            I => \N__24018\
        );

    \I__5736\ : LocalMux
    port map (
            O => \N__24053\,
            I => \N__24014\
        );

    \I__5735\ : LocalMux
    port map (
            O => \N__24050\,
            I => \N__24011\
        );

    \I__5734\ : LocalMux
    port map (
            O => \N__24041\,
            I => \N__24006\
        );

    \I__5733\ : LocalMux
    port map (
            O => \N__24032\,
            I => \N__24006\
        );

    \I__5732\ : LocalMux
    port map (
            O => \N__24029\,
            I => \N__23999\
        );

    \I__5731\ : LocalMux
    port map (
            O => \N__24026\,
            I => \N__23996\
        );

    \I__5730\ : InMux
    port map (
            O => \N__24025\,
            I => \N__23991\
        );

    \I__5729\ : InMux
    port map (
            O => \N__24024\,
            I => \N__23991\
        );

    \I__5728\ : Span4Mux_v
    port map (
            O => \N__24021\,
            I => \N__23986\
        );

    \I__5727\ : LocalMux
    port map (
            O => \N__24018\,
            I => \N__23986\
        );

    \I__5726\ : InMux
    port map (
            O => \N__24017\,
            I => \N__23983\
        );

    \I__5725\ : Span4Mux_h
    port map (
            O => \N__24014\,
            I => \N__23977\
        );

    \I__5724\ : Span4Mux_v
    port map (
            O => \N__24011\,
            I => \N__23972\
        );

    \I__5723\ : Span4Mux_v
    port map (
            O => \N__24006\,
            I => \N__23972\
        );

    \I__5722\ : CascadeMux
    port map (
            O => \N__24005\,
            I => \N__23969\
        );

    \I__5721\ : InMux
    port map (
            O => \N__24004\,
            I => \N__23966\
        );

    \I__5720\ : CascadeMux
    port map (
            O => \N__24003\,
            I => \N__23963\
        );

    \I__5719\ : CascadeMux
    port map (
            O => \N__24002\,
            I => \N__23956\
        );

    \I__5718\ : Span4Mux_v
    port map (
            O => \N__23999\,
            I => \N__23947\
        );

    \I__5717\ : Span4Mux_h
    port map (
            O => \N__23996\,
            I => \N__23947\
        );

    \I__5716\ : LocalMux
    port map (
            O => \N__23991\,
            I => \N__23947\
        );

    \I__5715\ : Span4Mux_h
    port map (
            O => \N__23986\,
            I => \N__23947\
        );

    \I__5714\ : LocalMux
    port map (
            O => \N__23983\,
            I => \N__23944\
        );

    \I__5713\ : InMux
    port map (
            O => \N__23982\,
            I => \N__23937\
        );

    \I__5712\ : InMux
    port map (
            O => \N__23981\,
            I => \N__23937\
        );

    \I__5711\ : InMux
    port map (
            O => \N__23980\,
            I => \N__23937\
        );

    \I__5710\ : Span4Mux_v
    port map (
            O => \N__23977\,
            I => \N__23934\
        );

    \I__5709\ : Span4Mux_h
    port map (
            O => \N__23972\,
            I => \N__23931\
        );

    \I__5708\ : InMux
    port map (
            O => \N__23969\,
            I => \N__23928\
        );

    \I__5707\ : LocalMux
    port map (
            O => \N__23966\,
            I => \N__23925\
        );

    \I__5706\ : InMux
    port map (
            O => \N__23963\,
            I => \N__23920\
        );

    \I__5705\ : InMux
    port map (
            O => \N__23962\,
            I => \N__23920\
        );

    \I__5704\ : InMux
    port map (
            O => \N__23961\,
            I => \N__23911\
        );

    \I__5703\ : InMux
    port map (
            O => \N__23960\,
            I => \N__23911\
        );

    \I__5702\ : InMux
    port map (
            O => \N__23959\,
            I => \N__23911\
        );

    \I__5701\ : InMux
    port map (
            O => \N__23956\,
            I => \N__23911\
        );

    \I__5700\ : Span4Mux_v
    port map (
            O => \N__23947\,
            I => \N__23908\
        );

    \I__5699\ : Odrv4
    port map (
            O => \N__23944\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_2\
        );

    \I__5698\ : LocalMux
    port map (
            O => \N__23937\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_2\
        );

    \I__5697\ : Odrv4
    port map (
            O => \N__23934\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_2\
        );

    \I__5696\ : Odrv4
    port map (
            O => \N__23931\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_2\
        );

    \I__5695\ : LocalMux
    port map (
            O => \N__23928\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_2\
        );

    \I__5694\ : Odrv12
    port map (
            O => \N__23925\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_2\
        );

    \I__5693\ : LocalMux
    port map (
            O => \N__23920\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_2\
        );

    \I__5692\ : LocalMux
    port map (
            O => \N__23911\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_2\
        );

    \I__5691\ : Odrv4
    port map (
            O => \N__23908\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_2\
        );

    \I__5690\ : InMux
    port map (
            O => \N__23889\,
            I => \N__23886\
        );

    \I__5689\ : LocalMux
    port map (
            O => \N__23886\,
            I => \ppm_encoder_1.pulses2countZ0Z_0\
        );

    \I__5688\ : ClkMux
    port map (
            O => \N__23883\,
            I => \N__23577\
        );

    \I__5687\ : ClkMux
    port map (
            O => \N__23882\,
            I => \N__23577\
        );

    \I__5686\ : ClkMux
    port map (
            O => \N__23881\,
            I => \N__23577\
        );

    \I__5685\ : ClkMux
    port map (
            O => \N__23880\,
            I => \N__23577\
        );

    \I__5684\ : ClkMux
    port map (
            O => \N__23879\,
            I => \N__23577\
        );

    \I__5683\ : ClkMux
    port map (
            O => \N__23878\,
            I => \N__23577\
        );

    \I__5682\ : ClkMux
    port map (
            O => \N__23877\,
            I => \N__23577\
        );

    \I__5681\ : ClkMux
    port map (
            O => \N__23876\,
            I => \N__23577\
        );

    \I__5680\ : ClkMux
    port map (
            O => \N__23875\,
            I => \N__23577\
        );

    \I__5679\ : ClkMux
    port map (
            O => \N__23874\,
            I => \N__23577\
        );

    \I__5678\ : ClkMux
    port map (
            O => \N__23873\,
            I => \N__23577\
        );

    \I__5677\ : ClkMux
    port map (
            O => \N__23872\,
            I => \N__23577\
        );

    \I__5676\ : ClkMux
    port map (
            O => \N__23871\,
            I => \N__23577\
        );

    \I__5675\ : ClkMux
    port map (
            O => \N__23870\,
            I => \N__23577\
        );

    \I__5674\ : ClkMux
    port map (
            O => \N__23869\,
            I => \N__23577\
        );

    \I__5673\ : ClkMux
    port map (
            O => \N__23868\,
            I => \N__23577\
        );

    \I__5672\ : ClkMux
    port map (
            O => \N__23867\,
            I => \N__23577\
        );

    \I__5671\ : ClkMux
    port map (
            O => \N__23866\,
            I => \N__23577\
        );

    \I__5670\ : ClkMux
    port map (
            O => \N__23865\,
            I => \N__23577\
        );

    \I__5669\ : ClkMux
    port map (
            O => \N__23864\,
            I => \N__23577\
        );

    \I__5668\ : ClkMux
    port map (
            O => \N__23863\,
            I => \N__23577\
        );

    \I__5667\ : ClkMux
    port map (
            O => \N__23862\,
            I => \N__23577\
        );

    \I__5666\ : ClkMux
    port map (
            O => \N__23861\,
            I => \N__23577\
        );

    \I__5665\ : ClkMux
    port map (
            O => \N__23860\,
            I => \N__23577\
        );

    \I__5664\ : ClkMux
    port map (
            O => \N__23859\,
            I => \N__23577\
        );

    \I__5663\ : ClkMux
    port map (
            O => \N__23858\,
            I => \N__23577\
        );

    \I__5662\ : ClkMux
    port map (
            O => \N__23857\,
            I => \N__23577\
        );

    \I__5661\ : ClkMux
    port map (
            O => \N__23856\,
            I => \N__23577\
        );

    \I__5660\ : ClkMux
    port map (
            O => \N__23855\,
            I => \N__23577\
        );

    \I__5659\ : ClkMux
    port map (
            O => \N__23854\,
            I => \N__23577\
        );

    \I__5658\ : ClkMux
    port map (
            O => \N__23853\,
            I => \N__23577\
        );

    \I__5657\ : ClkMux
    port map (
            O => \N__23852\,
            I => \N__23577\
        );

    \I__5656\ : ClkMux
    port map (
            O => \N__23851\,
            I => \N__23577\
        );

    \I__5655\ : ClkMux
    port map (
            O => \N__23850\,
            I => \N__23577\
        );

    \I__5654\ : ClkMux
    port map (
            O => \N__23849\,
            I => \N__23577\
        );

    \I__5653\ : ClkMux
    port map (
            O => \N__23848\,
            I => \N__23577\
        );

    \I__5652\ : ClkMux
    port map (
            O => \N__23847\,
            I => \N__23577\
        );

    \I__5651\ : ClkMux
    port map (
            O => \N__23846\,
            I => \N__23577\
        );

    \I__5650\ : ClkMux
    port map (
            O => \N__23845\,
            I => \N__23577\
        );

    \I__5649\ : ClkMux
    port map (
            O => \N__23844\,
            I => \N__23577\
        );

    \I__5648\ : ClkMux
    port map (
            O => \N__23843\,
            I => \N__23577\
        );

    \I__5647\ : ClkMux
    port map (
            O => \N__23842\,
            I => \N__23577\
        );

    \I__5646\ : ClkMux
    port map (
            O => \N__23841\,
            I => \N__23577\
        );

    \I__5645\ : ClkMux
    port map (
            O => \N__23840\,
            I => \N__23577\
        );

    \I__5644\ : ClkMux
    port map (
            O => \N__23839\,
            I => \N__23577\
        );

    \I__5643\ : ClkMux
    port map (
            O => \N__23838\,
            I => \N__23577\
        );

    \I__5642\ : ClkMux
    port map (
            O => \N__23837\,
            I => \N__23577\
        );

    \I__5641\ : ClkMux
    port map (
            O => \N__23836\,
            I => \N__23577\
        );

    \I__5640\ : ClkMux
    port map (
            O => \N__23835\,
            I => \N__23577\
        );

    \I__5639\ : ClkMux
    port map (
            O => \N__23834\,
            I => \N__23577\
        );

    \I__5638\ : ClkMux
    port map (
            O => \N__23833\,
            I => \N__23577\
        );

    \I__5637\ : ClkMux
    port map (
            O => \N__23832\,
            I => \N__23577\
        );

    \I__5636\ : ClkMux
    port map (
            O => \N__23831\,
            I => \N__23577\
        );

    \I__5635\ : ClkMux
    port map (
            O => \N__23830\,
            I => \N__23577\
        );

    \I__5634\ : ClkMux
    port map (
            O => \N__23829\,
            I => \N__23577\
        );

    \I__5633\ : ClkMux
    port map (
            O => \N__23828\,
            I => \N__23577\
        );

    \I__5632\ : ClkMux
    port map (
            O => \N__23827\,
            I => \N__23577\
        );

    \I__5631\ : ClkMux
    port map (
            O => \N__23826\,
            I => \N__23577\
        );

    \I__5630\ : ClkMux
    port map (
            O => \N__23825\,
            I => \N__23577\
        );

    \I__5629\ : ClkMux
    port map (
            O => \N__23824\,
            I => \N__23577\
        );

    \I__5628\ : ClkMux
    port map (
            O => \N__23823\,
            I => \N__23577\
        );

    \I__5627\ : ClkMux
    port map (
            O => \N__23822\,
            I => \N__23577\
        );

    \I__5626\ : ClkMux
    port map (
            O => \N__23821\,
            I => \N__23577\
        );

    \I__5625\ : ClkMux
    port map (
            O => \N__23820\,
            I => \N__23577\
        );

    \I__5624\ : ClkMux
    port map (
            O => \N__23819\,
            I => \N__23577\
        );

    \I__5623\ : ClkMux
    port map (
            O => \N__23818\,
            I => \N__23577\
        );

    \I__5622\ : ClkMux
    port map (
            O => \N__23817\,
            I => \N__23577\
        );

    \I__5621\ : ClkMux
    port map (
            O => \N__23816\,
            I => \N__23577\
        );

    \I__5620\ : ClkMux
    port map (
            O => \N__23815\,
            I => \N__23577\
        );

    \I__5619\ : ClkMux
    port map (
            O => \N__23814\,
            I => \N__23577\
        );

    \I__5618\ : ClkMux
    port map (
            O => \N__23813\,
            I => \N__23577\
        );

    \I__5617\ : ClkMux
    port map (
            O => \N__23812\,
            I => \N__23577\
        );

    \I__5616\ : ClkMux
    port map (
            O => \N__23811\,
            I => \N__23577\
        );

    \I__5615\ : ClkMux
    port map (
            O => \N__23810\,
            I => \N__23577\
        );

    \I__5614\ : ClkMux
    port map (
            O => \N__23809\,
            I => \N__23577\
        );

    \I__5613\ : ClkMux
    port map (
            O => \N__23808\,
            I => \N__23577\
        );

    \I__5612\ : ClkMux
    port map (
            O => \N__23807\,
            I => \N__23577\
        );

    \I__5611\ : ClkMux
    port map (
            O => \N__23806\,
            I => \N__23577\
        );

    \I__5610\ : ClkMux
    port map (
            O => \N__23805\,
            I => \N__23577\
        );

    \I__5609\ : ClkMux
    port map (
            O => \N__23804\,
            I => \N__23577\
        );

    \I__5608\ : ClkMux
    port map (
            O => \N__23803\,
            I => \N__23577\
        );

    \I__5607\ : ClkMux
    port map (
            O => \N__23802\,
            I => \N__23577\
        );

    \I__5606\ : ClkMux
    port map (
            O => \N__23801\,
            I => \N__23577\
        );

    \I__5605\ : ClkMux
    port map (
            O => \N__23800\,
            I => \N__23577\
        );

    \I__5604\ : ClkMux
    port map (
            O => \N__23799\,
            I => \N__23577\
        );

    \I__5603\ : ClkMux
    port map (
            O => \N__23798\,
            I => \N__23577\
        );

    \I__5602\ : ClkMux
    port map (
            O => \N__23797\,
            I => \N__23577\
        );

    \I__5601\ : ClkMux
    port map (
            O => \N__23796\,
            I => \N__23577\
        );

    \I__5600\ : ClkMux
    port map (
            O => \N__23795\,
            I => \N__23577\
        );

    \I__5599\ : ClkMux
    port map (
            O => \N__23794\,
            I => \N__23577\
        );

    \I__5598\ : ClkMux
    port map (
            O => \N__23793\,
            I => \N__23577\
        );

    \I__5597\ : ClkMux
    port map (
            O => \N__23792\,
            I => \N__23577\
        );

    \I__5596\ : ClkMux
    port map (
            O => \N__23791\,
            I => \N__23577\
        );

    \I__5595\ : ClkMux
    port map (
            O => \N__23790\,
            I => \N__23577\
        );

    \I__5594\ : ClkMux
    port map (
            O => \N__23789\,
            I => \N__23577\
        );

    \I__5593\ : ClkMux
    port map (
            O => \N__23788\,
            I => \N__23577\
        );

    \I__5592\ : ClkMux
    port map (
            O => \N__23787\,
            I => \N__23577\
        );

    \I__5591\ : ClkMux
    port map (
            O => \N__23786\,
            I => \N__23577\
        );

    \I__5590\ : ClkMux
    port map (
            O => \N__23785\,
            I => \N__23577\
        );

    \I__5589\ : ClkMux
    port map (
            O => \N__23784\,
            I => \N__23577\
        );

    \I__5588\ : ClkMux
    port map (
            O => \N__23783\,
            I => \N__23577\
        );

    \I__5587\ : ClkMux
    port map (
            O => \N__23782\,
            I => \N__23577\
        );

    \I__5586\ : GlobalMux
    port map (
            O => \N__23577\,
            I => \N__23574\
        );

    \I__5585\ : gio2CtrlBuf
    port map (
            O => \N__23574\,
            I => clk_system_c_g
        );

    \I__5584\ : CEMux
    port map (
            O => \N__23571\,
            I => \N__23541\
        );

    \I__5583\ : CEMux
    port map (
            O => \N__23570\,
            I => \N__23541\
        );

    \I__5582\ : CEMux
    port map (
            O => \N__23569\,
            I => \N__23541\
        );

    \I__5581\ : CEMux
    port map (
            O => \N__23568\,
            I => \N__23541\
        );

    \I__5580\ : CEMux
    port map (
            O => \N__23567\,
            I => \N__23541\
        );

    \I__5579\ : CEMux
    port map (
            O => \N__23566\,
            I => \N__23541\
        );

    \I__5578\ : CEMux
    port map (
            O => \N__23565\,
            I => \N__23541\
        );

    \I__5577\ : CEMux
    port map (
            O => \N__23564\,
            I => \N__23541\
        );

    \I__5576\ : CEMux
    port map (
            O => \N__23563\,
            I => \N__23541\
        );

    \I__5575\ : CEMux
    port map (
            O => \N__23562\,
            I => \N__23541\
        );

    \I__5574\ : GlobalMux
    port map (
            O => \N__23541\,
            I => \N__23538\
        );

    \I__5573\ : gio2CtrlBuf
    port map (
            O => \N__23538\,
            I => \ppm_encoder_1.N_238_i_0_g\
        );

    \I__5572\ : CascadeMux
    port map (
            O => \N__23535\,
            I => \N__23527\
        );

    \I__5571\ : CascadeMux
    port map (
            O => \N__23534\,
            I => \N__23524\
        );

    \I__5570\ : CascadeMux
    port map (
            O => \N__23533\,
            I => \N__23517\
        );

    \I__5569\ : CascadeMux
    port map (
            O => \N__23532\,
            I => \N__23514\
        );

    \I__5568\ : CascadeMux
    port map (
            O => \N__23531\,
            I => \N__23508\
        );

    \I__5567\ : InMux
    port map (
            O => \N__23530\,
            I => \N__23487\
        );

    \I__5566\ : InMux
    port map (
            O => \N__23527\,
            I => \N__23482\
        );

    \I__5565\ : InMux
    port map (
            O => \N__23524\,
            I => \N__23482\
        );

    \I__5564\ : InMux
    port map (
            O => \N__23523\,
            I => \N__23479\
        );

    \I__5563\ : InMux
    port map (
            O => \N__23522\,
            I => \N__23476\
        );

    \I__5562\ : InMux
    port map (
            O => \N__23521\,
            I => \N__23473\
        );

    \I__5561\ : InMux
    port map (
            O => \N__23520\,
            I => \N__23470\
        );

    \I__5560\ : InMux
    port map (
            O => \N__23517\,
            I => \N__23463\
        );

    \I__5559\ : InMux
    port map (
            O => \N__23514\,
            I => \N__23463\
        );

    \I__5558\ : InMux
    port map (
            O => \N__23513\,
            I => \N__23463\
        );

    \I__5557\ : InMux
    port map (
            O => \N__23512\,
            I => \N__23460\
        );

    \I__5556\ : InMux
    port map (
            O => \N__23511\,
            I => \N__23457\
        );

    \I__5555\ : InMux
    port map (
            O => \N__23508\,
            I => \N__23450\
        );

    \I__5554\ : InMux
    port map (
            O => \N__23507\,
            I => \N__23450\
        );

    \I__5553\ : InMux
    port map (
            O => \N__23506\,
            I => \N__23450\
        );

    \I__5552\ : InMux
    port map (
            O => \N__23505\,
            I => \N__23445\
        );

    \I__5551\ : InMux
    port map (
            O => \N__23504\,
            I => \N__23445\
        );

    \I__5550\ : InMux
    port map (
            O => \N__23503\,
            I => \N__23442\
        );

    \I__5549\ : InMux
    port map (
            O => \N__23502\,
            I => \N__23439\
        );

    \I__5548\ : InMux
    port map (
            O => \N__23501\,
            I => \N__23436\
        );

    \I__5547\ : InMux
    port map (
            O => \N__23500\,
            I => \N__23433\
        );

    \I__5546\ : InMux
    port map (
            O => \N__23499\,
            I => \N__23428\
        );

    \I__5545\ : InMux
    port map (
            O => \N__23498\,
            I => \N__23428\
        );

    \I__5544\ : InMux
    port map (
            O => \N__23497\,
            I => \N__23425\
        );

    \I__5543\ : InMux
    port map (
            O => \N__23496\,
            I => \N__23422\
        );

    \I__5542\ : InMux
    port map (
            O => \N__23495\,
            I => \N__23415\
        );

    \I__5541\ : InMux
    port map (
            O => \N__23494\,
            I => \N__23415\
        );

    \I__5540\ : InMux
    port map (
            O => \N__23493\,
            I => \N__23415\
        );

    \I__5539\ : InMux
    port map (
            O => \N__23492\,
            I => \N__23412\
        );

    \I__5538\ : InMux
    port map (
            O => \N__23491\,
            I => \N__23409\
        );

    \I__5537\ : InMux
    port map (
            O => \N__23490\,
            I => \N__23406\
        );

    \I__5536\ : LocalMux
    port map (
            O => \N__23487\,
            I => \N__23338\
        );

    \I__5535\ : LocalMux
    port map (
            O => \N__23482\,
            I => \N__23335\
        );

    \I__5534\ : LocalMux
    port map (
            O => \N__23479\,
            I => \N__23332\
        );

    \I__5533\ : LocalMux
    port map (
            O => \N__23476\,
            I => \N__23329\
        );

    \I__5532\ : LocalMux
    port map (
            O => \N__23473\,
            I => \N__23326\
        );

    \I__5531\ : LocalMux
    port map (
            O => \N__23470\,
            I => \N__23323\
        );

    \I__5530\ : LocalMux
    port map (
            O => \N__23463\,
            I => \N__23320\
        );

    \I__5529\ : LocalMux
    port map (
            O => \N__23460\,
            I => \N__23317\
        );

    \I__5528\ : LocalMux
    port map (
            O => \N__23457\,
            I => \N__23314\
        );

    \I__5527\ : LocalMux
    port map (
            O => \N__23450\,
            I => \N__23311\
        );

    \I__5526\ : LocalMux
    port map (
            O => \N__23445\,
            I => \N__23308\
        );

    \I__5525\ : LocalMux
    port map (
            O => \N__23442\,
            I => \N__23305\
        );

    \I__5524\ : LocalMux
    port map (
            O => \N__23439\,
            I => \N__23302\
        );

    \I__5523\ : LocalMux
    port map (
            O => \N__23436\,
            I => \N__23299\
        );

    \I__5522\ : LocalMux
    port map (
            O => \N__23433\,
            I => \N__23296\
        );

    \I__5521\ : LocalMux
    port map (
            O => \N__23428\,
            I => \N__23293\
        );

    \I__5520\ : LocalMux
    port map (
            O => \N__23425\,
            I => \N__23290\
        );

    \I__5519\ : LocalMux
    port map (
            O => \N__23422\,
            I => \N__23287\
        );

    \I__5518\ : LocalMux
    port map (
            O => \N__23415\,
            I => \N__23284\
        );

    \I__5517\ : LocalMux
    port map (
            O => \N__23412\,
            I => \N__23281\
        );

    \I__5516\ : LocalMux
    port map (
            O => \N__23409\,
            I => \N__23278\
        );

    \I__5515\ : LocalMux
    port map (
            O => \N__23406\,
            I => \N__23275\
        );

    \I__5514\ : SRMux
    port map (
            O => \N__23405\,
            I => \N__23100\
        );

    \I__5513\ : SRMux
    port map (
            O => \N__23404\,
            I => \N__23100\
        );

    \I__5512\ : SRMux
    port map (
            O => \N__23403\,
            I => \N__23100\
        );

    \I__5511\ : SRMux
    port map (
            O => \N__23402\,
            I => \N__23100\
        );

    \I__5510\ : SRMux
    port map (
            O => \N__23401\,
            I => \N__23100\
        );

    \I__5509\ : SRMux
    port map (
            O => \N__23400\,
            I => \N__23100\
        );

    \I__5508\ : SRMux
    port map (
            O => \N__23399\,
            I => \N__23100\
        );

    \I__5507\ : SRMux
    port map (
            O => \N__23398\,
            I => \N__23100\
        );

    \I__5506\ : SRMux
    port map (
            O => \N__23397\,
            I => \N__23100\
        );

    \I__5505\ : SRMux
    port map (
            O => \N__23396\,
            I => \N__23100\
        );

    \I__5504\ : SRMux
    port map (
            O => \N__23395\,
            I => \N__23100\
        );

    \I__5503\ : SRMux
    port map (
            O => \N__23394\,
            I => \N__23100\
        );

    \I__5502\ : SRMux
    port map (
            O => \N__23393\,
            I => \N__23100\
        );

    \I__5501\ : SRMux
    port map (
            O => \N__23392\,
            I => \N__23100\
        );

    \I__5500\ : SRMux
    port map (
            O => \N__23391\,
            I => \N__23100\
        );

    \I__5499\ : SRMux
    port map (
            O => \N__23390\,
            I => \N__23100\
        );

    \I__5498\ : SRMux
    port map (
            O => \N__23389\,
            I => \N__23100\
        );

    \I__5497\ : SRMux
    port map (
            O => \N__23388\,
            I => \N__23100\
        );

    \I__5496\ : SRMux
    port map (
            O => \N__23387\,
            I => \N__23100\
        );

    \I__5495\ : SRMux
    port map (
            O => \N__23386\,
            I => \N__23100\
        );

    \I__5494\ : SRMux
    port map (
            O => \N__23385\,
            I => \N__23100\
        );

    \I__5493\ : SRMux
    port map (
            O => \N__23384\,
            I => \N__23100\
        );

    \I__5492\ : SRMux
    port map (
            O => \N__23383\,
            I => \N__23100\
        );

    \I__5491\ : SRMux
    port map (
            O => \N__23382\,
            I => \N__23100\
        );

    \I__5490\ : SRMux
    port map (
            O => \N__23381\,
            I => \N__23100\
        );

    \I__5489\ : SRMux
    port map (
            O => \N__23380\,
            I => \N__23100\
        );

    \I__5488\ : SRMux
    port map (
            O => \N__23379\,
            I => \N__23100\
        );

    \I__5487\ : SRMux
    port map (
            O => \N__23378\,
            I => \N__23100\
        );

    \I__5486\ : SRMux
    port map (
            O => \N__23377\,
            I => \N__23100\
        );

    \I__5485\ : SRMux
    port map (
            O => \N__23376\,
            I => \N__23100\
        );

    \I__5484\ : SRMux
    port map (
            O => \N__23375\,
            I => \N__23100\
        );

    \I__5483\ : SRMux
    port map (
            O => \N__23374\,
            I => \N__23100\
        );

    \I__5482\ : SRMux
    port map (
            O => \N__23373\,
            I => \N__23100\
        );

    \I__5481\ : SRMux
    port map (
            O => \N__23372\,
            I => \N__23100\
        );

    \I__5480\ : SRMux
    port map (
            O => \N__23371\,
            I => \N__23100\
        );

    \I__5479\ : SRMux
    port map (
            O => \N__23370\,
            I => \N__23100\
        );

    \I__5478\ : SRMux
    port map (
            O => \N__23369\,
            I => \N__23100\
        );

    \I__5477\ : SRMux
    port map (
            O => \N__23368\,
            I => \N__23100\
        );

    \I__5476\ : SRMux
    port map (
            O => \N__23367\,
            I => \N__23100\
        );

    \I__5475\ : SRMux
    port map (
            O => \N__23366\,
            I => \N__23100\
        );

    \I__5474\ : SRMux
    port map (
            O => \N__23365\,
            I => \N__23100\
        );

    \I__5473\ : SRMux
    port map (
            O => \N__23364\,
            I => \N__23100\
        );

    \I__5472\ : SRMux
    port map (
            O => \N__23363\,
            I => \N__23100\
        );

    \I__5471\ : SRMux
    port map (
            O => \N__23362\,
            I => \N__23100\
        );

    \I__5470\ : SRMux
    port map (
            O => \N__23361\,
            I => \N__23100\
        );

    \I__5469\ : SRMux
    port map (
            O => \N__23360\,
            I => \N__23100\
        );

    \I__5468\ : SRMux
    port map (
            O => \N__23359\,
            I => \N__23100\
        );

    \I__5467\ : SRMux
    port map (
            O => \N__23358\,
            I => \N__23100\
        );

    \I__5466\ : SRMux
    port map (
            O => \N__23357\,
            I => \N__23100\
        );

    \I__5465\ : SRMux
    port map (
            O => \N__23356\,
            I => \N__23100\
        );

    \I__5464\ : SRMux
    port map (
            O => \N__23355\,
            I => \N__23100\
        );

    \I__5463\ : SRMux
    port map (
            O => \N__23354\,
            I => \N__23100\
        );

    \I__5462\ : SRMux
    port map (
            O => \N__23353\,
            I => \N__23100\
        );

    \I__5461\ : SRMux
    port map (
            O => \N__23352\,
            I => \N__23100\
        );

    \I__5460\ : SRMux
    port map (
            O => \N__23351\,
            I => \N__23100\
        );

    \I__5459\ : SRMux
    port map (
            O => \N__23350\,
            I => \N__23100\
        );

    \I__5458\ : SRMux
    port map (
            O => \N__23349\,
            I => \N__23100\
        );

    \I__5457\ : SRMux
    port map (
            O => \N__23348\,
            I => \N__23100\
        );

    \I__5456\ : SRMux
    port map (
            O => \N__23347\,
            I => \N__23100\
        );

    \I__5455\ : SRMux
    port map (
            O => \N__23346\,
            I => \N__23100\
        );

    \I__5454\ : SRMux
    port map (
            O => \N__23345\,
            I => \N__23100\
        );

    \I__5453\ : SRMux
    port map (
            O => \N__23344\,
            I => \N__23100\
        );

    \I__5452\ : SRMux
    port map (
            O => \N__23343\,
            I => \N__23100\
        );

    \I__5451\ : SRMux
    port map (
            O => \N__23342\,
            I => \N__23100\
        );

    \I__5450\ : SRMux
    port map (
            O => \N__23341\,
            I => \N__23100\
        );

    \I__5449\ : Glb2LocalMux
    port map (
            O => \N__23338\,
            I => \N__23100\
        );

    \I__5448\ : Glb2LocalMux
    port map (
            O => \N__23335\,
            I => \N__23100\
        );

    \I__5447\ : Glb2LocalMux
    port map (
            O => \N__23332\,
            I => \N__23100\
        );

    \I__5446\ : Glb2LocalMux
    port map (
            O => \N__23329\,
            I => \N__23100\
        );

    \I__5445\ : Glb2LocalMux
    port map (
            O => \N__23326\,
            I => \N__23100\
        );

    \I__5444\ : Glb2LocalMux
    port map (
            O => \N__23323\,
            I => \N__23100\
        );

    \I__5443\ : Glb2LocalMux
    port map (
            O => \N__23320\,
            I => \N__23100\
        );

    \I__5442\ : Glb2LocalMux
    port map (
            O => \N__23317\,
            I => \N__23100\
        );

    \I__5441\ : Glb2LocalMux
    port map (
            O => \N__23314\,
            I => \N__23100\
        );

    \I__5440\ : Glb2LocalMux
    port map (
            O => \N__23311\,
            I => \N__23100\
        );

    \I__5439\ : Glb2LocalMux
    port map (
            O => \N__23308\,
            I => \N__23100\
        );

    \I__5438\ : Glb2LocalMux
    port map (
            O => \N__23305\,
            I => \N__23100\
        );

    \I__5437\ : Glb2LocalMux
    port map (
            O => \N__23302\,
            I => \N__23100\
        );

    \I__5436\ : Glb2LocalMux
    port map (
            O => \N__23299\,
            I => \N__23100\
        );

    \I__5435\ : Glb2LocalMux
    port map (
            O => \N__23296\,
            I => \N__23100\
        );

    \I__5434\ : Glb2LocalMux
    port map (
            O => \N__23293\,
            I => \N__23100\
        );

    \I__5433\ : Glb2LocalMux
    port map (
            O => \N__23290\,
            I => \N__23100\
        );

    \I__5432\ : Glb2LocalMux
    port map (
            O => \N__23287\,
            I => \N__23100\
        );

    \I__5431\ : Glb2LocalMux
    port map (
            O => \N__23284\,
            I => \N__23100\
        );

    \I__5430\ : Glb2LocalMux
    port map (
            O => \N__23281\,
            I => \N__23100\
        );

    \I__5429\ : Glb2LocalMux
    port map (
            O => \N__23278\,
            I => \N__23100\
        );

    \I__5428\ : Glb2LocalMux
    port map (
            O => \N__23275\,
            I => \N__23100\
        );

    \I__5427\ : GlobalMux
    port map (
            O => \N__23100\,
            I => \N__23097\
        );

    \I__5426\ : gio2CtrlBuf
    port map (
            O => \N__23097\,
            I => reset_system_g
        );

    \I__5425\ : InMux
    port map (
            O => \N__23094\,
            I => \N__23091\
        );

    \I__5424\ : LocalMux
    port map (
            O => \N__23091\,
            I => \ppm_encoder_1.counter24_0_I_1_c_RNOZ0\
        );

    \I__5423\ : InMux
    port map (
            O => \N__23088\,
            I => \N__23085\
        );

    \I__5422\ : LocalMux
    port map (
            O => \N__23085\,
            I => \N__23082\
        );

    \I__5421\ : Span4Mux_h
    port map (
            O => \N__23082\,
            I => \N__23079\
        );

    \I__5420\ : Odrv4
    port map (
            O => \N__23079\,
            I => \ppm_encoder_1.counter24_0_I_9_c_RNOZ0\
        );

    \I__5419\ : InMux
    port map (
            O => \N__23076\,
            I => \N__23073\
        );

    \I__5418\ : LocalMux
    port map (
            O => \N__23073\,
            I => \ppm_encoder_1.counter24_0_I_15_c_RNOZ0\
        );

    \I__5417\ : InMux
    port map (
            O => \N__23070\,
            I => \N__23067\
        );

    \I__5416\ : LocalMux
    port map (
            O => \N__23067\,
            I => \N__23064\
        );

    \I__5415\ : Odrv4
    port map (
            O => \N__23064\,
            I => \ppm_encoder_1.counter24_0_I_21_c_RNOZ0\
        );

    \I__5414\ : InMux
    port map (
            O => \N__23061\,
            I => \N__23058\
        );

    \I__5413\ : LocalMux
    port map (
            O => \N__23058\,
            I => \ppm_encoder_1.counter24_0_I_33_c_RNOZ0\
        );

    \I__5412\ : InMux
    port map (
            O => \N__23055\,
            I => \N__23052\
        );

    \I__5411\ : LocalMux
    port map (
            O => \N__23052\,
            I => \N__23049\
        );

    \I__5410\ : Odrv4
    port map (
            O => \N__23049\,
            I => \ppm_encoder_1.un1_PPM_STATE_0_sqmuxa_0_i_0_a2_1\
        );

    \I__5409\ : CascadeMux
    port map (
            O => \N__23046\,
            I => \ppm_encoder_1.un1_PPM_STATE_0_sqmuxa_0_i_0_a2_16_4_cascade_\
        );

    \I__5408\ : InMux
    port map (
            O => \N__23043\,
            I => \N__23040\
        );

    \I__5407\ : LocalMux
    port map (
            O => \N__23040\,
            I => \N__23037\
        );

    \I__5406\ : Span4Mux_v
    port map (
            O => \N__23037\,
            I => \N__23034\
        );

    \I__5405\ : Odrv4
    port map (
            O => \N__23034\,
            I => \ppm_encoder_1.pulses2countZ0Z_12\
        );

    \I__5404\ : CascadeMux
    port map (
            O => \N__23031\,
            I => \N__23028\
        );

    \I__5403\ : InMux
    port map (
            O => \N__23028\,
            I => \N__23025\
        );

    \I__5402\ : LocalMux
    port map (
            O => \N__23025\,
            I => \N__23022\
        );

    \I__5401\ : Odrv4
    port map (
            O => \N__23022\,
            I => \ppm_encoder_1.pulses2countZ0Z_13\
        );

    \I__5400\ : InMux
    port map (
            O => \N__23019\,
            I => \N__23014\
        );

    \I__5399\ : InMux
    port map (
            O => \N__23018\,
            I => \N__23009\
        );

    \I__5398\ : InMux
    port map (
            O => \N__23017\,
            I => \N__23009\
        );

    \I__5397\ : LocalMux
    port map (
            O => \N__23014\,
            I => \ppm_encoder_1.counterZ0Z_12\
        );

    \I__5396\ : LocalMux
    port map (
            O => \N__23009\,
            I => \ppm_encoder_1.counterZ0Z_12\
        );

    \I__5395\ : InMux
    port map (
            O => \N__23004\,
            I => \N__23001\
        );

    \I__5394\ : LocalMux
    port map (
            O => \N__23001\,
            I => \N__22998\
        );

    \I__5393\ : Odrv4
    port map (
            O => \N__22998\,
            I => \ppm_encoder_1.pulses2countZ0Z_18\
        );

    \I__5392\ : InMux
    port map (
            O => \N__22995\,
            I => \N__22991\
        );

    \I__5391\ : InMux
    port map (
            O => \N__22994\,
            I => \N__22987\
        );

    \I__5390\ : LocalMux
    port map (
            O => \N__22991\,
            I => \N__22984\
        );

    \I__5389\ : InMux
    port map (
            O => \N__22990\,
            I => \N__22981\
        );

    \I__5388\ : LocalMux
    port map (
            O => \N__22987\,
            I => \ppm_encoder_1.counterZ0Z_18\
        );

    \I__5387\ : Odrv4
    port map (
            O => \N__22984\,
            I => \ppm_encoder_1.counterZ0Z_18\
        );

    \I__5386\ : LocalMux
    port map (
            O => \N__22981\,
            I => \ppm_encoder_1.counterZ0Z_18\
        );

    \I__5385\ : InMux
    port map (
            O => \N__22974\,
            I => \N__22971\
        );

    \I__5384\ : LocalMux
    port map (
            O => \N__22971\,
            I => \ppm_encoder_1.un1_PPM_STATE_0_sqmuxa_0_i_0_a2_2_3\
        );

    \I__5383\ : InMux
    port map (
            O => \N__22968\,
            I => \N__22963\
        );

    \I__5382\ : InMux
    port map (
            O => \N__22967\,
            I => \N__22960\
        );

    \I__5381\ : InMux
    port map (
            O => \N__22966\,
            I => \N__22957\
        );

    \I__5380\ : LocalMux
    port map (
            O => \N__22963\,
            I => \ppm_encoder_1.counterZ0Z_15\
        );

    \I__5379\ : LocalMux
    port map (
            O => \N__22960\,
            I => \ppm_encoder_1.counterZ0Z_15\
        );

    \I__5378\ : LocalMux
    port map (
            O => \N__22957\,
            I => \ppm_encoder_1.counterZ0Z_15\
        );

    \I__5377\ : CascadeMux
    port map (
            O => \N__22950\,
            I => \N__22947\
        );

    \I__5376\ : InMux
    port map (
            O => \N__22947\,
            I => \N__22944\
        );

    \I__5375\ : LocalMux
    port map (
            O => \N__22944\,
            I => \N__22941\
        );

    \I__5374\ : Odrv4
    port map (
            O => \N__22941\,
            I => \ppm_encoder_1.un1_PPM_STATE_0_sqmuxa_0_i_0_a2_2_4\
        );

    \I__5373\ : InMux
    port map (
            O => \N__22938\,
            I => \N__22933\
        );

    \I__5372\ : InMux
    port map (
            O => \N__22937\,
            I => \N__22930\
        );

    \I__5371\ : InMux
    port map (
            O => \N__22936\,
            I => \N__22927\
        );

    \I__5370\ : LocalMux
    port map (
            O => \N__22933\,
            I => \ppm_encoder_1.counterZ0Z_13\
        );

    \I__5369\ : LocalMux
    port map (
            O => \N__22930\,
            I => \ppm_encoder_1.counterZ0Z_13\
        );

    \I__5368\ : LocalMux
    port map (
            O => \N__22927\,
            I => \ppm_encoder_1.counterZ0Z_13\
        );

    \I__5367\ : InMux
    port map (
            O => \N__22920\,
            I => \N__22917\
        );

    \I__5366\ : LocalMux
    port map (
            O => \N__22917\,
            I => \ppm_encoder_1.un1_PPM_STATE_0_sqmuxa_0_i_0_a2_2\
        );

    \I__5365\ : InMux
    port map (
            O => \N__22914\,
            I => \N__22911\
        );

    \I__5364\ : LocalMux
    port map (
            O => \N__22911\,
            I => \N__22908\
        );

    \I__5363\ : Odrv4
    port map (
            O => \N__22908\,
            I => \ppm_encoder_1.un1_PPM_STATE_1_sqmuxa_i_i_a2_0_1\
        );

    \I__5362\ : InMux
    port map (
            O => \N__22905\,
            I => \N__22902\
        );

    \I__5361\ : LocalMux
    port map (
            O => \N__22902\,
            I => \ppm_encoder_1.un1_PPM_STATE_0_sqmuxa_0_i_0_a2_16_4\
        );

    \I__5360\ : CascadeMux
    port map (
            O => \N__22899\,
            I => \ppm_encoder_1.un1_PPM_STATE_0_sqmuxa_0_i_0_a2_2_cascade_\
        );

    \I__5359\ : InMux
    port map (
            O => \N__22896\,
            I => \N__22892\
        );

    \I__5358\ : InMux
    port map (
            O => \N__22895\,
            I => \N__22889\
        );

    \I__5357\ : LocalMux
    port map (
            O => \N__22892\,
            I => \N__22886\
        );

    \I__5356\ : LocalMux
    port map (
            O => \N__22889\,
            I => \N__22883\
        );

    \I__5355\ : Span4Mux_v
    port map (
            O => \N__22886\,
            I => \N__22880\
        );

    \I__5354\ : Span4Mux_h
    port map (
            O => \N__22883\,
            I => \N__22877\
        );

    \I__5353\ : Odrv4
    port map (
            O => \N__22880\,
            I => \ppm_encoder_1.un1_PPM_STATE_0_sqmuxa_0_i_0_a2_16_5\
        );

    \I__5352\ : Odrv4
    port map (
            O => \N__22877\,
            I => \ppm_encoder_1.un1_PPM_STATE_0_sqmuxa_0_i_0_a2_16_5\
        );

    \I__5351\ : CascadeMux
    port map (
            O => \N__22872\,
            I => \N__22869\
        );

    \I__5350\ : InMux
    port map (
            O => \N__22869\,
            I => \N__22863\
        );

    \I__5349\ : InMux
    port map (
            O => \N__22868\,
            I => \N__22863\
        );

    \I__5348\ : LocalMux
    port map (
            O => \N__22863\,
            I => \N__22859\
        );

    \I__5347\ : InMux
    port map (
            O => \N__22862\,
            I => \N__22856\
        );

    \I__5346\ : Odrv12
    port map (
            O => \N__22859\,
            I => \ppm_encoder_1.counter24_0_I_57_c_RNIJMMDZ0\
        );

    \I__5345\ : LocalMux
    port map (
            O => \N__22856\,
            I => \ppm_encoder_1.counter24_0_I_57_c_RNIJMMDZ0\
        );

    \I__5344\ : CascadeMux
    port map (
            O => \N__22851\,
            I => \ppm_encoder_1.N_431_cascade_\
        );

    \I__5343\ : InMux
    port map (
            O => \N__22848\,
            I => \N__22845\
        );

    \I__5342\ : LocalMux
    port map (
            O => \N__22845\,
            I => \N__22842\
        );

    \I__5341\ : Span4Mux_h
    port map (
            O => \N__22842\,
            I => \N__22832\
        );

    \I__5340\ : InMux
    port map (
            O => \N__22841\,
            I => \N__22825\
        );

    \I__5339\ : InMux
    port map (
            O => \N__22840\,
            I => \N__22825\
        );

    \I__5338\ : InMux
    port map (
            O => \N__22839\,
            I => \N__22825\
        );

    \I__5337\ : InMux
    port map (
            O => \N__22838\,
            I => \N__22822\
        );

    \I__5336\ : InMux
    port map (
            O => \N__22837\,
            I => \N__22819\
        );

    \I__5335\ : InMux
    port map (
            O => \N__22836\,
            I => \N__22814\
        );

    \I__5334\ : InMux
    port map (
            O => \N__22835\,
            I => \N__22814\
        );

    \I__5333\ : Odrv4
    port map (
            O => \N__22832\,
            I => \ppm_encoder_1.PPM_STATEZ0Z_1\
        );

    \I__5332\ : LocalMux
    port map (
            O => \N__22825\,
            I => \ppm_encoder_1.PPM_STATEZ0Z_1\
        );

    \I__5331\ : LocalMux
    port map (
            O => \N__22822\,
            I => \ppm_encoder_1.PPM_STATEZ0Z_1\
        );

    \I__5330\ : LocalMux
    port map (
            O => \N__22819\,
            I => \ppm_encoder_1.PPM_STATEZ0Z_1\
        );

    \I__5329\ : LocalMux
    port map (
            O => \N__22814\,
            I => \ppm_encoder_1.PPM_STATEZ0Z_1\
        );

    \I__5328\ : IoInMux
    port map (
            O => \N__22803\,
            I => \N__22800\
        );

    \I__5327\ : LocalMux
    port map (
            O => \N__22800\,
            I => \N__22797\
        );

    \I__5326\ : IoSpan4Mux
    port map (
            O => \N__22797\,
            I => \N__22794\
        );

    \I__5325\ : Span4Mux_s3_v
    port map (
            O => \N__22794\,
            I => \N__22791\
        );

    \I__5324\ : Sp12to4
    port map (
            O => \N__22791\,
            I => \N__22788\
        );

    \I__5323\ : Span12Mux_v
    port map (
            O => \N__22788\,
            I => \N__22784\
        );

    \I__5322\ : InMux
    port map (
            O => \N__22787\,
            I => \N__22781\
        );

    \I__5321\ : Odrv12
    port map (
            O => \N__22784\,
            I => ppm_output_c
        );

    \I__5320\ : LocalMux
    port map (
            O => \N__22781\,
            I => ppm_output_c
        );

    \I__5319\ : InMux
    port map (
            O => \N__22776\,
            I => \N__22773\
        );

    \I__5318\ : LocalMux
    port map (
            O => \N__22773\,
            I => \ppm_encoder_1.pulses2countZ0Z_16\
        );

    \I__5317\ : CascadeMux
    port map (
            O => \N__22770\,
            I => \N__22767\
        );

    \I__5316\ : InMux
    port map (
            O => \N__22767\,
            I => \N__22763\
        );

    \I__5315\ : InMux
    port map (
            O => \N__22766\,
            I => \N__22759\
        );

    \I__5314\ : LocalMux
    port map (
            O => \N__22763\,
            I => \N__22756\
        );

    \I__5313\ : InMux
    port map (
            O => \N__22762\,
            I => \N__22753\
        );

    \I__5312\ : LocalMux
    port map (
            O => \N__22759\,
            I => \ppm_encoder_1.counterZ0Z_17\
        );

    \I__5311\ : Odrv4
    port map (
            O => \N__22756\,
            I => \ppm_encoder_1.counterZ0Z_17\
        );

    \I__5310\ : LocalMux
    port map (
            O => \N__22753\,
            I => \ppm_encoder_1.counterZ0Z_17\
        );

    \I__5309\ : CascadeMux
    port map (
            O => \N__22746\,
            I => \N__22743\
        );

    \I__5308\ : InMux
    port map (
            O => \N__22743\,
            I => \N__22740\
        );

    \I__5307\ : LocalMux
    port map (
            O => \N__22740\,
            I => \N__22737\
        );

    \I__5306\ : Odrv12
    port map (
            O => \N__22737\,
            I => \ppm_encoder_1.pulses2countZ0Z_17\
        );

    \I__5305\ : InMux
    port map (
            O => \N__22734\,
            I => \N__22729\
        );

    \I__5304\ : InMux
    port map (
            O => \N__22733\,
            I => \N__22726\
        );

    \I__5303\ : InMux
    port map (
            O => \N__22732\,
            I => \N__22723\
        );

    \I__5302\ : LocalMux
    port map (
            O => \N__22729\,
            I => \ppm_encoder_1.counterZ0Z_16\
        );

    \I__5301\ : LocalMux
    port map (
            O => \N__22726\,
            I => \ppm_encoder_1.counterZ0Z_16\
        );

    \I__5300\ : LocalMux
    port map (
            O => \N__22723\,
            I => \ppm_encoder_1.counterZ0Z_16\
        );

    \I__5299\ : InMux
    port map (
            O => \N__22716\,
            I => \N__22713\
        );

    \I__5298\ : LocalMux
    port map (
            O => \N__22713\,
            I => \N__22710\
        );

    \I__5297\ : Span4Mux_h
    port map (
            O => \N__22710\,
            I => \N__22707\
        );

    \I__5296\ : Odrv4
    port map (
            O => \N__22707\,
            I => \ppm_encoder_1.pulses2count_9_i_1_8\
        );

    \I__5295\ : InMux
    port map (
            O => \N__22704\,
            I => \N__22699\
        );

    \I__5294\ : CascadeMux
    port map (
            O => \N__22703\,
            I => \N__22696\
        );

    \I__5293\ : CascadeMux
    port map (
            O => \N__22702\,
            I => \N__22693\
        );

    \I__5292\ : LocalMux
    port map (
            O => \N__22699\,
            I => \N__22689\
        );

    \I__5291\ : InMux
    port map (
            O => \N__22696\,
            I => \N__22684\
        );

    \I__5290\ : InMux
    port map (
            O => \N__22693\,
            I => \N__22684\
        );

    \I__5289\ : InMux
    port map (
            O => \N__22692\,
            I => \N__22681\
        );

    \I__5288\ : Span4Mux_v
    port map (
            O => \N__22689\,
            I => \N__22676\
        );

    \I__5287\ : LocalMux
    port map (
            O => \N__22684\,
            I => \N__22676\
        );

    \I__5286\ : LocalMux
    port map (
            O => \N__22681\,
            I => \N__22673\
        );

    \I__5285\ : Span4Mux_h
    port map (
            O => \N__22676\,
            I => \N__22670\
        );

    \I__5284\ : Span4Mux_v
    port map (
            O => \N__22673\,
            I => \N__22667\
        );

    \I__5283\ : Span4Mux_v
    port map (
            O => \N__22670\,
            I => \N__22664\
        );

    \I__5282\ : Span4Mux_v
    port map (
            O => \N__22667\,
            I => \N__22661\
        );

    \I__5281\ : Odrv4
    port map (
            O => \N__22664\,
            I => \ppm_encoder_1.init_pulsesZ0Z_8\
        );

    \I__5280\ : Odrv4
    port map (
            O => \N__22661\,
            I => \ppm_encoder_1.init_pulsesZ0Z_8\
        );

    \I__5279\ : InMux
    port map (
            O => \N__22656\,
            I => \N__22653\
        );

    \I__5278\ : LocalMux
    port map (
            O => \N__22653\,
            I => \N__22650\
        );

    \I__5277\ : Span4Mux_h
    port map (
            O => \N__22650\,
            I => \N__22647\
        );

    \I__5276\ : Odrv4
    port map (
            O => \N__22647\,
            I => \ppm_encoder_1.pulses2count_9_i_1_4\
        );

    \I__5275\ : InMux
    port map (
            O => \N__22644\,
            I => \N__22641\
        );

    \I__5274\ : LocalMux
    port map (
            O => \N__22641\,
            I => \N__22636\
        );

    \I__5273\ : CascadeMux
    port map (
            O => \N__22640\,
            I => \N__22633\
        );

    \I__5272\ : InMux
    port map (
            O => \N__22639\,
            I => \N__22629\
        );

    \I__5271\ : Span12Mux_s8_v
    port map (
            O => \N__22636\,
            I => \N__22626\
        );

    \I__5270\ : InMux
    port map (
            O => \N__22633\,
            I => \N__22623\
        );

    \I__5269\ : InMux
    port map (
            O => \N__22632\,
            I => \N__22620\
        );

    \I__5268\ : LocalMux
    port map (
            O => \N__22629\,
            I => \N__22617\
        );

    \I__5267\ : Odrv12
    port map (
            O => \N__22626\,
            I => \ppm_encoder_1.init_pulsesZ0Z_4\
        );

    \I__5266\ : LocalMux
    port map (
            O => \N__22623\,
            I => \ppm_encoder_1.init_pulsesZ0Z_4\
        );

    \I__5265\ : LocalMux
    port map (
            O => \N__22620\,
            I => \ppm_encoder_1.init_pulsesZ0Z_4\
        );

    \I__5264\ : Odrv4
    port map (
            O => \N__22617\,
            I => \ppm_encoder_1.init_pulsesZ0Z_4\
        );

    \I__5263\ : InMux
    port map (
            O => \N__22608\,
            I => \N__22605\
        );

    \I__5262\ : LocalMux
    port map (
            O => \N__22605\,
            I => \ppm_encoder_1.pulses2countZ0Z_4\
        );

    \I__5261\ : InMux
    port map (
            O => \N__22602\,
            I => \N__22599\
        );

    \I__5260\ : LocalMux
    port map (
            O => \N__22599\,
            I => \N__22596\
        );

    \I__5259\ : Span4Mux_h
    port map (
            O => \N__22596\,
            I => \N__22593\
        );

    \I__5258\ : Odrv4
    port map (
            O => \N__22593\,
            I => \ppm_encoder_1.N_300\
        );

    \I__5257\ : CascadeMux
    port map (
            O => \N__22590\,
            I => \N__22587\
        );

    \I__5256\ : InMux
    port map (
            O => \N__22587\,
            I => \N__22584\
        );

    \I__5255\ : LocalMux
    port map (
            O => \N__22584\,
            I => \N__22581\
        );

    \I__5254\ : Odrv4
    port map (
            O => \N__22581\,
            I => \ppm_encoder_1.pulses2count_9_i_0_5\
        );

    \I__5253\ : InMux
    port map (
            O => \N__22578\,
            I => \N__22573\
        );

    \I__5252\ : CascadeMux
    port map (
            O => \N__22577\,
            I => \N__22570\
        );

    \I__5251\ : CascadeMux
    port map (
            O => \N__22576\,
            I => \N__22566\
        );

    \I__5250\ : LocalMux
    port map (
            O => \N__22573\,
            I => \N__22563\
        );

    \I__5249\ : InMux
    port map (
            O => \N__22570\,
            I => \N__22560\
        );

    \I__5248\ : InMux
    port map (
            O => \N__22569\,
            I => \N__22557\
        );

    \I__5247\ : InMux
    port map (
            O => \N__22566\,
            I => \N__22554\
        );

    \I__5246\ : Span4Mux_h
    port map (
            O => \N__22563\,
            I => \N__22549\
        );

    \I__5245\ : LocalMux
    port map (
            O => \N__22560\,
            I => \N__22549\
        );

    \I__5244\ : LocalMux
    port map (
            O => \N__22557\,
            I => \N__22544\
        );

    \I__5243\ : LocalMux
    port map (
            O => \N__22554\,
            I => \N__22544\
        );

    \I__5242\ : Odrv4
    port map (
            O => \N__22549\,
            I => \ppm_encoder_1.init_pulsesZ0Z_5\
        );

    \I__5241\ : Odrv12
    port map (
            O => \N__22544\,
            I => \ppm_encoder_1.init_pulsesZ0Z_5\
        );

    \I__5240\ : CascadeMux
    port map (
            O => \N__22539\,
            I => \N__22536\
        );

    \I__5239\ : InMux
    port map (
            O => \N__22536\,
            I => \N__22533\
        );

    \I__5238\ : LocalMux
    port map (
            O => \N__22533\,
            I => \ppm_encoder_1.pulses2countZ0Z_5\
        );

    \I__5237\ : CascadeMux
    port map (
            O => \N__22530\,
            I => \N__22527\
        );

    \I__5236\ : InMux
    port map (
            O => \N__22527\,
            I => \N__22522\
        );

    \I__5235\ : InMux
    port map (
            O => \N__22526\,
            I => \N__22519\
        );

    \I__5234\ : InMux
    port map (
            O => \N__22525\,
            I => \N__22516\
        );

    \I__5233\ : LocalMux
    port map (
            O => \N__22522\,
            I => \N__22513\
        );

    \I__5232\ : LocalMux
    port map (
            O => \N__22519\,
            I => \N__22509\
        );

    \I__5231\ : LocalMux
    port map (
            O => \N__22516\,
            I => \N__22506\
        );

    \I__5230\ : Span4Mux_v
    port map (
            O => \N__22513\,
            I => \N__22503\
        );

    \I__5229\ : InMux
    port map (
            O => \N__22512\,
            I => \N__22500\
        );

    \I__5228\ : Span4Mux_h
    port map (
            O => \N__22509\,
            I => \N__22495\
        );

    \I__5227\ : Span4Mux_h
    port map (
            O => \N__22506\,
            I => \N__22495\
        );

    \I__5226\ : Odrv4
    port map (
            O => \N__22503\,
            I => \ppm_encoder_1.init_pulsesZ0Z_10\
        );

    \I__5225\ : LocalMux
    port map (
            O => \N__22500\,
            I => \ppm_encoder_1.init_pulsesZ0Z_10\
        );

    \I__5224\ : Odrv4
    port map (
            O => \N__22495\,
            I => \ppm_encoder_1.init_pulsesZ0Z_10\
        );

    \I__5223\ : InMux
    port map (
            O => \N__22488\,
            I => \N__22485\
        );

    \I__5222\ : LocalMux
    port map (
            O => \N__22485\,
            I => \N__22482\
        );

    \I__5221\ : Span4Mux_h
    port map (
            O => \N__22482\,
            I => \N__22479\
        );

    \I__5220\ : Odrv4
    port map (
            O => \N__22479\,
            I => \ppm_encoder_1.pulses2count_9_i_1_10\
        );

    \I__5219\ : InMux
    port map (
            O => \N__22476\,
            I => \N__22473\
        );

    \I__5218\ : LocalMux
    port map (
            O => \N__22473\,
            I => \ppm_encoder_1.pulses2countZ0Z_10\
        );

    \I__5217\ : CascadeMux
    port map (
            O => \N__22470\,
            I => \N__22465\
        );

    \I__5216\ : CascadeMux
    port map (
            O => \N__22469\,
            I => \N__22462\
        );

    \I__5215\ : InMux
    port map (
            O => \N__22468\,
            I => \N__22458\
        );

    \I__5214\ : InMux
    port map (
            O => \N__22465\,
            I => \N__22455\
        );

    \I__5213\ : InMux
    port map (
            O => \N__22462\,
            I => \N__22452\
        );

    \I__5212\ : InMux
    port map (
            O => \N__22461\,
            I => \N__22449\
        );

    \I__5211\ : LocalMux
    port map (
            O => \N__22458\,
            I => \ppm_encoder_1.counterZ0Z_11\
        );

    \I__5210\ : LocalMux
    port map (
            O => \N__22455\,
            I => \ppm_encoder_1.counterZ0Z_11\
        );

    \I__5209\ : LocalMux
    port map (
            O => \N__22452\,
            I => \ppm_encoder_1.counterZ0Z_11\
        );

    \I__5208\ : LocalMux
    port map (
            O => \N__22449\,
            I => \ppm_encoder_1.counterZ0Z_11\
        );

    \I__5207\ : CascadeMux
    port map (
            O => \N__22440\,
            I => \N__22437\
        );

    \I__5206\ : InMux
    port map (
            O => \N__22437\,
            I => \N__22434\
        );

    \I__5205\ : LocalMux
    port map (
            O => \N__22434\,
            I => \N__22431\
        );

    \I__5204\ : Odrv4
    port map (
            O => \N__22431\,
            I => \ppm_encoder_1.pulses2countZ0Z_11\
        );

    \I__5203\ : CascadeMux
    port map (
            O => \N__22428\,
            I => \N__22424\
        );

    \I__5202\ : InMux
    port map (
            O => \N__22427\,
            I => \N__22420\
        );

    \I__5201\ : InMux
    port map (
            O => \N__22424\,
            I => \N__22417\
        );

    \I__5200\ : InMux
    port map (
            O => \N__22423\,
            I => \N__22414\
        );

    \I__5199\ : LocalMux
    port map (
            O => \N__22420\,
            I => \ppm_encoder_1.counterZ0Z_10\
        );

    \I__5198\ : LocalMux
    port map (
            O => \N__22417\,
            I => \ppm_encoder_1.counterZ0Z_10\
        );

    \I__5197\ : LocalMux
    port map (
            O => \N__22414\,
            I => \ppm_encoder_1.counterZ0Z_10\
        );

    \I__5196\ : InMux
    port map (
            O => \N__22407\,
            I => \N__22404\
        );

    \I__5195\ : LocalMux
    port map (
            O => \N__22404\,
            I => \N__22401\
        );

    \I__5194\ : Odrv4
    port map (
            O => \N__22401\,
            I => \ppm_encoder_1.pulses2countZ0Z_14\
        );

    \I__5193\ : CascadeMux
    port map (
            O => \N__22398\,
            I => \N__22395\
        );

    \I__5192\ : InMux
    port map (
            O => \N__22395\,
            I => \N__22392\
        );

    \I__5191\ : LocalMux
    port map (
            O => \N__22392\,
            I => \N__22389\
        );

    \I__5190\ : Odrv4
    port map (
            O => \N__22389\,
            I => \ppm_encoder_1.pulses2countZ0Z_15\
        );

    \I__5189\ : InMux
    port map (
            O => \N__22386\,
            I => \N__22381\
        );

    \I__5188\ : InMux
    port map (
            O => \N__22385\,
            I => \N__22378\
        );

    \I__5187\ : InMux
    port map (
            O => \N__22384\,
            I => \N__22375\
        );

    \I__5186\ : LocalMux
    port map (
            O => \N__22381\,
            I => \ppm_encoder_1.counterZ0Z_7\
        );

    \I__5185\ : LocalMux
    port map (
            O => \N__22378\,
            I => \ppm_encoder_1.counterZ0Z_7\
        );

    \I__5184\ : LocalMux
    port map (
            O => \N__22375\,
            I => \ppm_encoder_1.counterZ0Z_7\
        );

    \I__5183\ : InMux
    port map (
            O => \N__22368\,
            I => \N__22363\
        );

    \I__5182\ : InMux
    port map (
            O => \N__22367\,
            I => \N__22360\
        );

    \I__5181\ : InMux
    port map (
            O => \N__22366\,
            I => \N__22357\
        );

    \I__5180\ : LocalMux
    port map (
            O => \N__22363\,
            I => \ppm_encoder_1.counterZ0Z_5\
        );

    \I__5179\ : LocalMux
    port map (
            O => \N__22360\,
            I => \ppm_encoder_1.counterZ0Z_5\
        );

    \I__5178\ : LocalMux
    port map (
            O => \N__22357\,
            I => \ppm_encoder_1.counterZ0Z_5\
        );

    \I__5177\ : CascadeMux
    port map (
            O => \N__22350\,
            I => \N__22346\
        );

    \I__5176\ : InMux
    port map (
            O => \N__22349\,
            I => \N__22342\
        );

    \I__5175\ : InMux
    port map (
            O => \N__22346\,
            I => \N__22339\
        );

    \I__5174\ : InMux
    port map (
            O => \N__22345\,
            I => \N__22336\
        );

    \I__5173\ : LocalMux
    port map (
            O => \N__22342\,
            I => \ppm_encoder_1.counterZ0Z_14\
        );

    \I__5172\ : LocalMux
    port map (
            O => \N__22339\,
            I => \ppm_encoder_1.counterZ0Z_14\
        );

    \I__5171\ : LocalMux
    port map (
            O => \N__22336\,
            I => \ppm_encoder_1.counterZ0Z_14\
        );

    \I__5170\ : InMux
    port map (
            O => \N__22329\,
            I => \N__22324\
        );

    \I__5169\ : InMux
    port map (
            O => \N__22328\,
            I => \N__22321\
        );

    \I__5168\ : InMux
    port map (
            O => \N__22327\,
            I => \N__22318\
        );

    \I__5167\ : LocalMux
    port map (
            O => \N__22324\,
            I => \ppm_encoder_1.counterZ0Z_6\
        );

    \I__5166\ : LocalMux
    port map (
            O => \N__22321\,
            I => \ppm_encoder_1.counterZ0Z_6\
        );

    \I__5165\ : LocalMux
    port map (
            O => \N__22318\,
            I => \ppm_encoder_1.counterZ0Z_6\
        );

    \I__5164\ : InMux
    port map (
            O => \N__22311\,
            I => \N__22307\
        );

    \I__5163\ : CascadeMux
    port map (
            O => \N__22310\,
            I => \N__22304\
        );

    \I__5162\ : LocalMux
    port map (
            O => \N__22307\,
            I => \N__22300\
        );

    \I__5161\ : InMux
    port map (
            O => \N__22304\,
            I => \N__22297\
        );

    \I__5160\ : InMux
    port map (
            O => \N__22303\,
            I => \N__22294\
        );

    \I__5159\ : Odrv12
    port map (
            O => \N__22300\,
            I => \ppm_encoder_1.rudderZ0Z_5\
        );

    \I__5158\ : LocalMux
    port map (
            O => \N__22297\,
            I => \ppm_encoder_1.rudderZ0Z_5\
        );

    \I__5157\ : LocalMux
    port map (
            O => \N__22294\,
            I => \ppm_encoder_1.rudderZ0Z_5\
        );

    \I__5156\ : CascadeMux
    port map (
            O => \N__22287\,
            I => \N__22284\
        );

    \I__5155\ : InMux
    port map (
            O => \N__22284\,
            I => \N__22280\
        );

    \I__5154\ : CascadeMux
    port map (
            O => \N__22283\,
            I => \N__22276\
        );

    \I__5153\ : LocalMux
    port map (
            O => \N__22280\,
            I => \N__22273\
        );

    \I__5152\ : CascadeMux
    port map (
            O => \N__22279\,
            I => \N__22270\
        );

    \I__5151\ : InMux
    port map (
            O => \N__22276\,
            I => \N__22266\
        );

    \I__5150\ : Span4Mux_h
    port map (
            O => \N__22273\,
            I => \N__22263\
        );

    \I__5149\ : InMux
    port map (
            O => \N__22270\,
            I => \N__22258\
        );

    \I__5148\ : InMux
    port map (
            O => \N__22269\,
            I => \N__22258\
        );

    \I__5147\ : LocalMux
    port map (
            O => \N__22266\,
            I => \ppm_encoder_1.rudderZ0Z_7\
        );

    \I__5146\ : Odrv4
    port map (
            O => \N__22263\,
            I => \ppm_encoder_1.rudderZ0Z_7\
        );

    \I__5145\ : LocalMux
    port map (
            O => \N__22258\,
            I => \ppm_encoder_1.rudderZ0Z_7\
        );

    \I__5144\ : CascadeMux
    port map (
            O => \N__22251\,
            I => \N__22248\
        );

    \I__5143\ : InMux
    port map (
            O => \N__22248\,
            I => \N__22245\
        );

    \I__5142\ : LocalMux
    port map (
            O => \N__22245\,
            I => \N__22242\
        );

    \I__5141\ : Span4Mux_h
    port map (
            O => \N__22242\,
            I => \N__22239\
        );

    \I__5140\ : Odrv4
    port map (
            O => \N__22239\,
            I => \ppm_encoder_1.pulses2count_9_i_0_7\
        );

    \I__5139\ : InMux
    port map (
            O => \N__22236\,
            I => \N__22232\
        );

    \I__5138\ : CascadeMux
    port map (
            O => \N__22235\,
            I => \N__22228\
        );

    \I__5137\ : LocalMux
    port map (
            O => \N__22232\,
            I => \N__22225\
        );

    \I__5136\ : InMux
    port map (
            O => \N__22231\,
            I => \N__22222\
        );

    \I__5135\ : InMux
    port map (
            O => \N__22228\,
            I => \N__22219\
        );

    \I__5134\ : Span4Mux_h
    port map (
            O => \N__22225\,
            I => \N__22216\
        );

    \I__5133\ : LocalMux
    port map (
            O => \N__22222\,
            I => \N__22213\
        );

    \I__5132\ : LocalMux
    port map (
            O => \N__22219\,
            I => \N__22210\
        );

    \I__5131\ : Span4Mux_h
    port map (
            O => \N__22216\,
            I => \N__22207\
        );

    \I__5130\ : Span4Mux_v
    port map (
            O => \N__22213\,
            I => \N__22204\
        );

    \I__5129\ : Span4Mux_h
    port map (
            O => \N__22210\,
            I => \N__22201\
        );

    \I__5128\ : Odrv4
    port map (
            O => \N__22207\,
            I => \ppm_encoder_1.init_pulsesZ0Z_0\
        );

    \I__5127\ : Odrv4
    port map (
            O => \N__22204\,
            I => \ppm_encoder_1.init_pulsesZ0Z_0\
        );

    \I__5126\ : Odrv4
    port map (
            O => \N__22201\,
            I => \ppm_encoder_1.init_pulsesZ0Z_0\
        );

    \I__5125\ : InMux
    port map (
            O => \N__22194\,
            I => \N__22191\
        );

    \I__5124\ : LocalMux
    port map (
            O => \N__22191\,
            I => \N__22188\
        );

    \I__5123\ : Span4Mux_h
    port map (
            O => \N__22188\,
            I => \N__22182\
        );

    \I__5122\ : InMux
    port map (
            O => \N__22187\,
            I => \N__22179\
        );

    \I__5121\ : InMux
    port map (
            O => \N__22186\,
            I => \N__22176\
        );

    \I__5120\ : InMux
    port map (
            O => \N__22185\,
            I => \N__22173\
        );

    \I__5119\ : Odrv4
    port map (
            O => \N__22182\,
            I => \ppm_encoder_1.counterZ0Z_1\
        );

    \I__5118\ : LocalMux
    port map (
            O => \N__22179\,
            I => \ppm_encoder_1.counterZ0Z_1\
        );

    \I__5117\ : LocalMux
    port map (
            O => \N__22176\,
            I => \ppm_encoder_1.counterZ0Z_1\
        );

    \I__5116\ : LocalMux
    port map (
            O => \N__22173\,
            I => \ppm_encoder_1.counterZ0Z_1\
        );

    \I__5115\ : CascadeMux
    port map (
            O => \N__22164\,
            I => \N__22161\
        );

    \I__5114\ : InMux
    port map (
            O => \N__22161\,
            I => \N__22158\
        );

    \I__5113\ : LocalMux
    port map (
            O => \N__22158\,
            I => \ppm_encoder_1.pulses2countZ0Z_1\
        );

    \I__5112\ : InMux
    port map (
            O => \N__22155\,
            I => \N__22151\
        );

    \I__5111\ : InMux
    port map (
            O => \N__22154\,
            I => \N__22147\
        );

    \I__5110\ : LocalMux
    port map (
            O => \N__22151\,
            I => \N__22144\
        );

    \I__5109\ : InMux
    port map (
            O => \N__22150\,
            I => \N__22141\
        );

    \I__5108\ : LocalMux
    port map (
            O => \N__22147\,
            I => \ppm_encoder_1.counterZ0Z_0\
        );

    \I__5107\ : Odrv4
    port map (
            O => \N__22144\,
            I => \ppm_encoder_1.counterZ0Z_0\
        );

    \I__5106\ : LocalMux
    port map (
            O => \N__22141\,
            I => \ppm_encoder_1.counterZ0Z_0\
        );

    \I__5105\ : CascadeMux
    port map (
            O => \N__22134\,
            I => \N__22129\
        );

    \I__5104\ : CascadeMux
    port map (
            O => \N__22133\,
            I => \N__22126\
        );

    \I__5103\ : InMux
    port map (
            O => \N__22132\,
            I => \N__22111\
        );

    \I__5102\ : InMux
    port map (
            O => \N__22129\,
            I => \N__22111\
        );

    \I__5101\ : InMux
    port map (
            O => \N__22126\,
            I => \N__22105\
        );

    \I__5100\ : InMux
    port map (
            O => \N__22125\,
            I => \N__22105\
        );

    \I__5099\ : InMux
    port map (
            O => \N__22124\,
            I => \N__22102\
        );

    \I__5098\ : InMux
    port map (
            O => \N__22123\,
            I => \N__22099\
        );

    \I__5097\ : InMux
    port map (
            O => \N__22122\,
            I => \N__22091\
        );

    \I__5096\ : InMux
    port map (
            O => \N__22121\,
            I => \N__22091\
        );

    \I__5095\ : InMux
    port map (
            O => \N__22120\,
            I => \N__22084\
        );

    \I__5094\ : InMux
    port map (
            O => \N__22119\,
            I => \N__22084\
        );

    \I__5093\ : InMux
    port map (
            O => \N__22118\,
            I => \N__22084\
        );

    \I__5092\ : InMux
    port map (
            O => \N__22117\,
            I => \N__22079\
        );

    \I__5091\ : InMux
    port map (
            O => \N__22116\,
            I => \N__22079\
        );

    \I__5090\ : LocalMux
    port map (
            O => \N__22111\,
            I => \N__22076\
        );

    \I__5089\ : InMux
    port map (
            O => \N__22110\,
            I => \N__22073\
        );

    \I__5088\ : LocalMux
    port map (
            O => \N__22105\,
            I => \N__22069\
        );

    \I__5087\ : LocalMux
    port map (
            O => \N__22102\,
            I => \N__22063\
        );

    \I__5086\ : LocalMux
    port map (
            O => \N__22099\,
            I => \N__22063\
        );

    \I__5085\ : CascadeMux
    port map (
            O => \N__22098\,
            I => \N__22060\
        );

    \I__5084\ : InMux
    port map (
            O => \N__22097\,
            I => \N__22053\
        );

    \I__5083\ : InMux
    port map (
            O => \N__22096\,
            I => \N__22053\
        );

    \I__5082\ : LocalMux
    port map (
            O => \N__22091\,
            I => \N__22050\
        );

    \I__5081\ : LocalMux
    port map (
            O => \N__22084\,
            I => \N__22045\
        );

    \I__5080\ : LocalMux
    port map (
            O => \N__22079\,
            I => \N__22045\
        );

    \I__5079\ : Span4Mux_v
    port map (
            O => \N__22076\,
            I => \N__22042\
        );

    \I__5078\ : LocalMux
    port map (
            O => \N__22073\,
            I => \N__22039\
        );

    \I__5077\ : InMux
    port map (
            O => \N__22072\,
            I => \N__22036\
        );

    \I__5076\ : Span4Mux_h
    port map (
            O => \N__22069\,
            I => \N__22033\
        );

    \I__5075\ : InMux
    port map (
            O => \N__22068\,
            I => \N__22030\
        );

    \I__5074\ : Span4Mux_v
    port map (
            O => \N__22063\,
            I => \N__22027\
        );

    \I__5073\ : InMux
    port map (
            O => \N__22060\,
            I => \N__22020\
        );

    \I__5072\ : InMux
    port map (
            O => \N__22059\,
            I => \N__22020\
        );

    \I__5071\ : InMux
    port map (
            O => \N__22058\,
            I => \N__22020\
        );

    \I__5070\ : LocalMux
    port map (
            O => \N__22053\,
            I => \N__22015\
        );

    \I__5069\ : Span4Mux_h
    port map (
            O => \N__22050\,
            I => \N__22015\
        );

    \I__5068\ : Span4Mux_v
    port map (
            O => \N__22045\,
            I => \N__22008\
        );

    \I__5067\ : Span4Mux_h
    port map (
            O => \N__22042\,
            I => \N__22008\
        );

    \I__5066\ : Span4Mux_h
    port map (
            O => \N__22039\,
            I => \N__22008\
        );

    \I__5065\ : LocalMux
    port map (
            O => \N__22036\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_1\
        );

    \I__5064\ : Odrv4
    port map (
            O => \N__22033\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_1\
        );

    \I__5063\ : LocalMux
    port map (
            O => \N__22030\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_1\
        );

    \I__5062\ : Odrv4
    port map (
            O => \N__22027\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_1\
        );

    \I__5061\ : LocalMux
    port map (
            O => \N__22020\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_1\
        );

    \I__5060\ : Odrv4
    port map (
            O => \N__22015\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_1\
        );

    \I__5059\ : Odrv4
    port map (
            O => \N__22008\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_1\
        );

    \I__5058\ : InMux
    port map (
            O => \N__21993\,
            I => \N__21982\
        );

    \I__5057\ : InMux
    port map (
            O => \N__21992\,
            I => \N__21982\
        );

    \I__5056\ : InMux
    port map (
            O => \N__21991\,
            I => \N__21982\
        );

    \I__5055\ : InMux
    port map (
            O => \N__21990\,
            I => \N__21968\
        );

    \I__5054\ : InMux
    port map (
            O => \N__21989\,
            I => \N__21968\
        );

    \I__5053\ : LocalMux
    port map (
            O => \N__21982\,
            I => \N__21961\
        );

    \I__5052\ : InMux
    port map (
            O => \N__21981\,
            I => \N__21954\
        );

    \I__5051\ : InMux
    port map (
            O => \N__21980\,
            I => \N__21954\
        );

    \I__5050\ : InMux
    port map (
            O => \N__21979\,
            I => \N__21954\
        );

    \I__5049\ : InMux
    port map (
            O => \N__21978\,
            I => \N__21951\
        );

    \I__5048\ : InMux
    port map (
            O => \N__21977\,
            I => \N__21948\
        );

    \I__5047\ : InMux
    port map (
            O => \N__21976\,
            I => \N__21943\
        );

    \I__5046\ : InMux
    port map (
            O => \N__21975\,
            I => \N__21943\
        );

    \I__5045\ : InMux
    port map (
            O => \N__21974\,
            I => \N__21939\
        );

    \I__5044\ : InMux
    port map (
            O => \N__21973\,
            I => \N__21936\
        );

    \I__5043\ : LocalMux
    port map (
            O => \N__21968\,
            I => \N__21933\
        );

    \I__5042\ : InMux
    port map (
            O => \N__21967\,
            I => \N__21930\
        );

    \I__5041\ : InMux
    port map (
            O => \N__21966\,
            I => \N__21925\
        );

    \I__5040\ : InMux
    port map (
            O => \N__21965\,
            I => \N__21920\
        );

    \I__5039\ : InMux
    port map (
            O => \N__21964\,
            I => \N__21920\
        );

    \I__5038\ : Span4Mux_v
    port map (
            O => \N__21961\,
            I => \N__21915\
        );

    \I__5037\ : LocalMux
    port map (
            O => \N__21954\,
            I => \N__21915\
        );

    \I__5036\ : LocalMux
    port map (
            O => \N__21951\,
            I => \N__21908\
        );

    \I__5035\ : LocalMux
    port map (
            O => \N__21948\,
            I => \N__21908\
        );

    \I__5034\ : LocalMux
    port map (
            O => \N__21943\,
            I => \N__21908\
        );

    \I__5033\ : InMux
    port map (
            O => \N__21942\,
            I => \N__21904\
        );

    \I__5032\ : LocalMux
    port map (
            O => \N__21939\,
            I => \N__21901\
        );

    \I__5031\ : LocalMux
    port map (
            O => \N__21936\,
            I => \N__21896\
        );

    \I__5030\ : Span4Mux_v
    port map (
            O => \N__21933\,
            I => \N__21896\
        );

    \I__5029\ : LocalMux
    port map (
            O => \N__21930\,
            I => \N__21893\
        );

    \I__5028\ : InMux
    port map (
            O => \N__21929\,
            I => \N__21888\
        );

    \I__5027\ : InMux
    port map (
            O => \N__21928\,
            I => \N__21888\
        );

    \I__5026\ : LocalMux
    port map (
            O => \N__21925\,
            I => \N__21883\
        );

    \I__5025\ : LocalMux
    port map (
            O => \N__21920\,
            I => \N__21883\
        );

    \I__5024\ : Span4Mux_v
    port map (
            O => \N__21915\,
            I => \N__21875\
        );

    \I__5023\ : Span4Mux_v
    port map (
            O => \N__21908\,
            I => \N__21875\
        );

    \I__5022\ : InMux
    port map (
            O => \N__21907\,
            I => \N__21872\
        );

    \I__5021\ : LocalMux
    port map (
            O => \N__21904\,
            I => \N__21869\
        );

    \I__5020\ : Span4Mux_v
    port map (
            O => \N__21901\,
            I => \N__21864\
        );

    \I__5019\ : Span4Mux_h
    port map (
            O => \N__21896\,
            I => \N__21864\
        );

    \I__5018\ : Span4Mux_h
    port map (
            O => \N__21893\,
            I => \N__21861\
        );

    \I__5017\ : LocalMux
    port map (
            O => \N__21888\,
            I => \N__21856\
        );

    \I__5016\ : Span4Mux_v
    port map (
            O => \N__21883\,
            I => \N__21856\
        );

    \I__5015\ : InMux
    port map (
            O => \N__21882\,
            I => \N__21849\
        );

    \I__5014\ : InMux
    port map (
            O => \N__21881\,
            I => \N__21849\
        );

    \I__5013\ : InMux
    port map (
            O => \N__21880\,
            I => \N__21849\
        );

    \I__5012\ : Span4Mux_h
    port map (
            O => \N__21875\,
            I => \N__21844\
        );

    \I__5011\ : LocalMux
    port map (
            O => \N__21872\,
            I => \N__21844\
        );

    \I__5010\ : Odrv4
    port map (
            O => \N__21869\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_0\
        );

    \I__5009\ : Odrv4
    port map (
            O => \N__21864\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_0\
        );

    \I__5008\ : Odrv4
    port map (
            O => \N__21861\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_0\
        );

    \I__5007\ : Odrv4
    port map (
            O => \N__21856\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_0\
        );

    \I__5006\ : LocalMux
    port map (
            O => \N__21849\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_0\
        );

    \I__5005\ : Odrv4
    port map (
            O => \N__21844\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_0\
        );

    \I__5004\ : CascadeMux
    port map (
            O => \N__21831\,
            I => \N__21827\
        );

    \I__5003\ : CascadeMux
    port map (
            O => \N__21830\,
            I => \N__21824\
        );

    \I__5002\ : InMux
    port map (
            O => \N__21827\,
            I => \N__21821\
        );

    \I__5001\ : InMux
    port map (
            O => \N__21824\,
            I => \N__21818\
        );

    \I__5000\ : LocalMux
    port map (
            O => \N__21821\,
            I => \N__21814\
        );

    \I__4999\ : LocalMux
    port map (
            O => \N__21818\,
            I => \N__21810\
        );

    \I__4998\ : CascadeMux
    port map (
            O => \N__21817\,
            I => \N__21807\
        );

    \I__4997\ : Span4Mux_h
    port map (
            O => \N__21814\,
            I => \N__21804\
        );

    \I__4996\ : InMux
    port map (
            O => \N__21813\,
            I => \N__21801\
        );

    \I__4995\ : Span4Mux_h
    port map (
            O => \N__21810\,
            I => \N__21798\
        );

    \I__4994\ : InMux
    port map (
            O => \N__21807\,
            I => \N__21795\
        );

    \I__4993\ : Odrv4
    port map (
            O => \N__21804\,
            I => \ppm_encoder_1.init_pulsesZ0Z_15\
        );

    \I__4992\ : LocalMux
    port map (
            O => \N__21801\,
            I => \ppm_encoder_1.init_pulsesZ0Z_15\
        );

    \I__4991\ : Odrv4
    port map (
            O => \N__21798\,
            I => \ppm_encoder_1.init_pulsesZ0Z_15\
        );

    \I__4990\ : LocalMux
    port map (
            O => \N__21795\,
            I => \ppm_encoder_1.init_pulsesZ0Z_15\
        );

    \I__4989\ : CascadeMux
    port map (
            O => \N__21786\,
            I => \N__21782\
        );

    \I__4988\ : InMux
    port map (
            O => \N__21785\,
            I => \N__21769\
        );

    \I__4987\ : InMux
    port map (
            O => \N__21782\,
            I => \N__21766\
        );

    \I__4986\ : InMux
    port map (
            O => \N__21781\,
            I => \N__21763\
        );

    \I__4985\ : InMux
    port map (
            O => \N__21780\,
            I => \N__21753\
        );

    \I__4984\ : InMux
    port map (
            O => \N__21779\,
            I => \N__21753\
        );

    \I__4983\ : InMux
    port map (
            O => \N__21778\,
            I => \N__21753\
        );

    \I__4982\ : InMux
    port map (
            O => \N__21777\,
            I => \N__21744\
        );

    \I__4981\ : InMux
    port map (
            O => \N__21776\,
            I => \N__21744\
        );

    \I__4980\ : InMux
    port map (
            O => \N__21775\,
            I => \N__21744\
        );

    \I__4979\ : InMux
    port map (
            O => \N__21774\,
            I => \N__21744\
        );

    \I__4978\ : CascadeMux
    port map (
            O => \N__21773\,
            I => \N__21741\
        );

    \I__4977\ : InMux
    port map (
            O => \N__21772\,
            I => \N__21738\
        );

    \I__4976\ : LocalMux
    port map (
            O => \N__21769\,
            I => \N__21735\
        );

    \I__4975\ : LocalMux
    port map (
            O => \N__21766\,
            I => \N__21730\
        );

    \I__4974\ : LocalMux
    port map (
            O => \N__21763\,
            I => \N__21727\
        );

    \I__4973\ : InMux
    port map (
            O => \N__21762\,
            I => \N__21722\
        );

    \I__4972\ : InMux
    port map (
            O => \N__21761\,
            I => \N__21722\
        );

    \I__4971\ : InMux
    port map (
            O => \N__21760\,
            I => \N__21719\
        );

    \I__4970\ : LocalMux
    port map (
            O => \N__21753\,
            I => \N__21716\
        );

    \I__4969\ : LocalMux
    port map (
            O => \N__21744\,
            I => \N__21713\
        );

    \I__4968\ : InMux
    port map (
            O => \N__21741\,
            I => \N__21710\
        );

    \I__4967\ : LocalMux
    port map (
            O => \N__21738\,
            I => \N__21707\
        );

    \I__4966\ : Span4Mux_h
    port map (
            O => \N__21735\,
            I => \N__21704\
        );

    \I__4965\ : CascadeMux
    port map (
            O => \N__21734\,
            I => \N__21699\
        );

    \I__4964\ : CascadeMux
    port map (
            O => \N__21733\,
            I => \N__21696\
        );

    \I__4963\ : Span4Mux_v
    port map (
            O => \N__21730\,
            I => \N__21691\
        );

    \I__4962\ : Span4Mux_h
    port map (
            O => \N__21727\,
            I => \N__21691\
        );

    \I__4961\ : LocalMux
    port map (
            O => \N__21722\,
            I => \N__21688\
        );

    \I__4960\ : LocalMux
    port map (
            O => \N__21719\,
            I => \N__21679\
        );

    \I__4959\ : Span4Mux_v
    port map (
            O => \N__21716\,
            I => \N__21679\
        );

    \I__4958\ : Span4Mux_v
    port map (
            O => \N__21713\,
            I => \N__21676\
        );

    \I__4957\ : LocalMux
    port map (
            O => \N__21710\,
            I => \N__21669\
        );

    \I__4956\ : Span4Mux_h
    port map (
            O => \N__21707\,
            I => \N__21669\
        );

    \I__4955\ : Span4Mux_v
    port map (
            O => \N__21704\,
            I => \N__21669\
        );

    \I__4954\ : InMux
    port map (
            O => \N__21703\,
            I => \N__21666\
        );

    \I__4953\ : InMux
    port map (
            O => \N__21702\,
            I => \N__21659\
        );

    \I__4952\ : InMux
    port map (
            O => \N__21699\,
            I => \N__21659\
        );

    \I__4951\ : InMux
    port map (
            O => \N__21696\,
            I => \N__21659\
        );

    \I__4950\ : Span4Mux_v
    port map (
            O => \N__21691\,
            I => \N__21654\
        );

    \I__4949\ : Span4Mux_h
    port map (
            O => \N__21688\,
            I => \N__21654\
        );

    \I__4948\ : InMux
    port map (
            O => \N__21687\,
            I => \N__21651\
        );

    \I__4947\ : InMux
    port map (
            O => \N__21686\,
            I => \N__21644\
        );

    \I__4946\ : InMux
    port map (
            O => \N__21685\,
            I => \N__21644\
        );

    \I__4945\ : InMux
    port map (
            O => \N__21684\,
            I => \N__21644\
        );

    \I__4944\ : Span4Mux_v
    port map (
            O => \N__21679\,
            I => \N__21637\
        );

    \I__4943\ : Span4Mux_v
    port map (
            O => \N__21676\,
            I => \N__21637\
        );

    \I__4942\ : Span4Mux_v
    port map (
            O => \N__21669\,
            I => \N__21637\
        );

    \I__4941\ : LocalMux
    port map (
            O => \N__21666\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_3\
        );

    \I__4940\ : LocalMux
    port map (
            O => \N__21659\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_3\
        );

    \I__4939\ : Odrv4
    port map (
            O => \N__21654\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_3\
        );

    \I__4938\ : LocalMux
    port map (
            O => \N__21651\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_3\
        );

    \I__4937\ : LocalMux
    port map (
            O => \N__21644\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_3\
        );

    \I__4936\ : Odrv4
    port map (
            O => \N__21637\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_3\
        );

    \I__4935\ : CascadeMux
    port map (
            O => \N__21624\,
            I => \N__21615\
        );

    \I__4934\ : CascadeMux
    port map (
            O => \N__21623\,
            I => \N__21611\
        );

    \I__4933\ : InMux
    port map (
            O => \N__21622\,
            I => \N__21606\
        );

    \I__4932\ : CascadeMux
    port map (
            O => \N__21621\,
            I => \N__21603\
        );

    \I__4931\ : CascadeMux
    port map (
            O => \N__21620\,
            I => \N__21599\
        );

    \I__4930\ : InMux
    port map (
            O => \N__21619\,
            I => \N__21594\
        );

    \I__4929\ : InMux
    port map (
            O => \N__21618\,
            I => \N__21594\
        );

    \I__4928\ : InMux
    port map (
            O => \N__21615\,
            I => \N__21585\
        );

    \I__4927\ : InMux
    port map (
            O => \N__21614\,
            I => \N__21585\
        );

    \I__4926\ : InMux
    port map (
            O => \N__21611\,
            I => \N__21585\
        );

    \I__4925\ : InMux
    port map (
            O => \N__21610\,
            I => \N__21585\
        );

    \I__4924\ : CascadeMux
    port map (
            O => \N__21609\,
            I => \N__21582\
        );

    \I__4923\ : LocalMux
    port map (
            O => \N__21606\,
            I => \N__21579\
        );

    \I__4922\ : InMux
    port map (
            O => \N__21603\,
            I => \N__21576\
        );

    \I__4921\ : InMux
    port map (
            O => \N__21602\,
            I => \N__21571\
        );

    \I__4920\ : InMux
    port map (
            O => \N__21599\,
            I => \N__21571\
        );

    \I__4919\ : LocalMux
    port map (
            O => \N__21594\,
            I => \N__21566\
        );

    \I__4918\ : LocalMux
    port map (
            O => \N__21585\,
            I => \N__21566\
        );

    \I__4917\ : InMux
    port map (
            O => \N__21582\,
            I => \N__21563\
        );

    \I__4916\ : Span4Mux_s3_v
    port map (
            O => \N__21579\,
            I => \N__21558\
        );

    \I__4915\ : LocalMux
    port map (
            O => \N__21576\,
            I => \N__21558\
        );

    \I__4914\ : LocalMux
    port map (
            O => \N__21571\,
            I => \N__21555\
        );

    \I__4913\ : Span4Mux_v
    port map (
            O => \N__21566\,
            I => \N__21552\
        );

    \I__4912\ : LocalMux
    port map (
            O => \N__21563\,
            I => \N__21545\
        );

    \I__4911\ : Span4Mux_v
    port map (
            O => \N__21558\,
            I => \N__21545\
        );

    \I__4910\ : Span4Mux_v
    port map (
            O => \N__21555\,
            I => \N__21545\
        );

    \I__4909\ : Odrv4
    port map (
            O => \N__21552\,
            I => \ppm_encoder_1.N_235\
        );

    \I__4908\ : Odrv4
    port map (
            O => \N__21545\,
            I => \ppm_encoder_1.N_235\
        );

    \I__4907\ : InMux
    port map (
            O => \N__21540\,
            I => \N__21536\
        );

    \I__4906\ : InMux
    port map (
            O => \N__21539\,
            I => \N__21533\
        );

    \I__4905\ : LocalMux
    port map (
            O => \N__21536\,
            I => \N__21530\
        );

    \I__4904\ : LocalMux
    port map (
            O => \N__21533\,
            I => \N__21527\
        );

    \I__4903\ : Span4Mux_v
    port map (
            O => \N__21530\,
            I => \N__21524\
        );

    \I__4902\ : Span12Mux_h
    port map (
            O => \N__21527\,
            I => \N__21521\
        );

    \I__4901\ : Span4Mux_h
    port map (
            O => \N__21524\,
            I => \N__21518\
        );

    \I__4900\ : Odrv12
    port map (
            O => \N__21521\,
            I => \ppm_encoder_1.rudderZ0Z_14\
        );

    \I__4899\ : Odrv4
    port map (
            O => \N__21518\,
            I => \ppm_encoder_1.rudderZ0Z_14\
        );

    \I__4898\ : InMux
    port map (
            O => \N__21513\,
            I => \N__21508\
        );

    \I__4897\ : CascadeMux
    port map (
            O => \N__21512\,
            I => \N__21504\
        );

    \I__4896\ : InMux
    port map (
            O => \N__21511\,
            I => \N__21501\
        );

    \I__4895\ : LocalMux
    port map (
            O => \N__21508\,
            I => \N__21498\
        );

    \I__4894\ : InMux
    port map (
            O => \N__21507\,
            I => \N__21495\
        );

    \I__4893\ : InMux
    port map (
            O => \N__21504\,
            I => \N__21492\
        );

    \I__4892\ : LocalMux
    port map (
            O => \N__21501\,
            I => \N__21489\
        );

    \I__4891\ : Span4Mux_h
    port map (
            O => \N__21498\,
            I => \N__21484\
        );

    \I__4890\ : LocalMux
    port map (
            O => \N__21495\,
            I => \N__21484\
        );

    \I__4889\ : LocalMux
    port map (
            O => \N__21492\,
            I => \N__21481\
        );

    \I__4888\ : Span4Mux_s3_v
    port map (
            O => \N__21489\,
            I => \N__21476\
        );

    \I__4887\ : Span4Mux_v
    port map (
            O => \N__21484\,
            I => \N__21476\
        );

    \I__4886\ : Odrv4
    port map (
            O => \N__21481\,
            I => \ppm_encoder_1.init_pulsesZ0Z_14\
        );

    \I__4885\ : Odrv4
    port map (
            O => \N__21476\,
            I => \ppm_encoder_1.init_pulsesZ0Z_14\
        );

    \I__4884\ : CascadeMux
    port map (
            O => \N__21471\,
            I => \ppm_encoder_1.pulses2count_9_i_0_14_cascade_\
        );

    \I__4883\ : InMux
    port map (
            O => \N__21468\,
            I => \N__21465\
        );

    \I__4882\ : LocalMux
    port map (
            O => \N__21465\,
            I => \N__21462\
        );

    \I__4881\ : Span12Mux_h
    port map (
            O => \N__21462\,
            I => \N__21458\
        );

    \I__4880\ : InMux
    port map (
            O => \N__21461\,
            I => \N__21455\
        );

    \I__4879\ : Odrv12
    port map (
            O => \N__21458\,
            I => \ppm_encoder_1.N_304\
        );

    \I__4878\ : LocalMux
    port map (
            O => \N__21455\,
            I => \ppm_encoder_1.N_304\
        );

    \I__4877\ : InMux
    port map (
            O => \N__21450\,
            I => \N__21446\
        );

    \I__4876\ : InMux
    port map (
            O => \N__21449\,
            I => \N__21442\
        );

    \I__4875\ : LocalMux
    port map (
            O => \N__21446\,
            I => \N__21439\
        );

    \I__4874\ : InMux
    port map (
            O => \N__21445\,
            I => \N__21436\
        );

    \I__4873\ : LocalMux
    port map (
            O => \N__21442\,
            I => \ppm_encoder_1.counterZ0Z_4\
        );

    \I__4872\ : Odrv4
    port map (
            O => \N__21439\,
            I => \ppm_encoder_1.counterZ0Z_4\
        );

    \I__4871\ : LocalMux
    port map (
            O => \N__21436\,
            I => \ppm_encoder_1.counterZ0Z_4\
        );

    \I__4870\ : InMux
    port map (
            O => \N__21429\,
            I => \ppm_encoder_1.un1_counter_13_cry_16\
        );

    \I__4869\ : InMux
    port map (
            O => \N__21426\,
            I => \ppm_encoder_1.un1_counter_13_cry_17\
        );

    \I__4868\ : SRMux
    port map (
            O => \N__21423\,
            I => \N__21414\
        );

    \I__4867\ : SRMux
    port map (
            O => \N__21422\,
            I => \N__21414\
        );

    \I__4866\ : SRMux
    port map (
            O => \N__21421\,
            I => \N__21414\
        );

    \I__4865\ : GlobalMux
    port map (
            O => \N__21414\,
            I => \N__21411\
        );

    \I__4864\ : gio2CtrlBuf
    port map (
            O => \N__21411\,
            I => \ppm_encoder_1.N_512_g\
        );

    \I__4863\ : InMux
    port map (
            O => \N__21408\,
            I => \N__21404\
        );

    \I__4862\ : InMux
    port map (
            O => \N__21407\,
            I => \N__21401\
        );

    \I__4861\ : LocalMux
    port map (
            O => \N__21404\,
            I => \N__21398\
        );

    \I__4860\ : LocalMux
    port map (
            O => \N__21401\,
            I => \N__21395\
        );

    \I__4859\ : Span4Mux_v
    port map (
            O => \N__21398\,
            I => \N__21389\
        );

    \I__4858\ : Span4Mux_h
    port map (
            O => \N__21395\,
            I => \N__21389\
        );

    \I__4857\ : InMux
    port map (
            O => \N__21394\,
            I => \N__21386\
        );

    \I__4856\ : Odrv4
    port map (
            O => \N__21389\,
            I => \ppm_encoder_1.N_247\
        );

    \I__4855\ : LocalMux
    port map (
            O => \N__21386\,
            I => \ppm_encoder_1.N_247\
        );

    \I__4854\ : InMux
    port map (
            O => \N__21381\,
            I => \N__21378\
        );

    \I__4853\ : LocalMux
    port map (
            O => \N__21378\,
            I => \ppm_encoder_1.pulses2count_9_0_2_11\
        );

    \I__4852\ : CascadeMux
    port map (
            O => \N__21375\,
            I => \N__21372\
        );

    \I__4851\ : InMux
    port map (
            O => \N__21372\,
            I => \N__21369\
        );

    \I__4850\ : LocalMux
    port map (
            O => \N__21369\,
            I => \ppm_encoder_1.N_388\
        );

    \I__4849\ : InMux
    port map (
            O => \N__21366\,
            I => \N__21363\
        );

    \I__4848\ : LocalMux
    port map (
            O => \N__21363\,
            I => \N__21360\
        );

    \I__4847\ : Span4Mux_h
    port map (
            O => \N__21360\,
            I => \N__21357\
        );

    \I__4846\ : Span4Mux_v
    port map (
            O => \N__21357\,
            I => \N__21354\
        );

    \I__4845\ : Odrv4
    port map (
            O => \N__21354\,
            I => \ppm_encoder_1.pulses2count_9_0_0_11\
        );

    \I__4844\ : CascadeMux
    port map (
            O => \N__21351\,
            I => \N__21346\
        );

    \I__4843\ : InMux
    port map (
            O => \N__21350\,
            I => \N__21343\
        );

    \I__4842\ : InMux
    port map (
            O => \N__21349\,
            I => \N__21340\
        );

    \I__4841\ : InMux
    port map (
            O => \N__21346\,
            I => \N__21337\
        );

    \I__4840\ : LocalMux
    port map (
            O => \N__21343\,
            I => \N__21333\
        );

    \I__4839\ : LocalMux
    port map (
            O => \N__21340\,
            I => \N__21330\
        );

    \I__4838\ : LocalMux
    port map (
            O => \N__21337\,
            I => \N__21327\
        );

    \I__4837\ : CascadeMux
    port map (
            O => \N__21336\,
            I => \N__21324\
        );

    \I__4836\ : Span4Mux_h
    port map (
            O => \N__21333\,
            I => \N__21321\
        );

    \I__4835\ : Sp12to4
    port map (
            O => \N__21330\,
            I => \N__21318\
        );

    \I__4834\ : Span4Mux_h
    port map (
            O => \N__21327\,
            I => \N__21315\
        );

    \I__4833\ : InMux
    port map (
            O => \N__21324\,
            I => \N__21312\
        );

    \I__4832\ : Odrv4
    port map (
            O => \N__21321\,
            I => \ppm_encoder_1.init_pulsesZ0Z_13\
        );

    \I__4831\ : Odrv12
    port map (
            O => \N__21318\,
            I => \ppm_encoder_1.init_pulsesZ0Z_13\
        );

    \I__4830\ : Odrv4
    port map (
            O => \N__21315\,
            I => \ppm_encoder_1.init_pulsesZ0Z_13\
        );

    \I__4829\ : LocalMux
    port map (
            O => \N__21312\,
            I => \ppm_encoder_1.init_pulsesZ0Z_13\
        );

    \I__4828\ : CascadeMux
    port map (
            O => \N__21303\,
            I => \N__21300\
        );

    \I__4827\ : InMux
    port map (
            O => \N__21300\,
            I => \N__21297\
        );

    \I__4826\ : LocalMux
    port map (
            O => \N__21297\,
            I => \ppm_encoder_1.pulses2count_9_0_0_13\
        );

    \I__4825\ : InMux
    port map (
            O => \N__21294\,
            I => \N__21291\
        );

    \I__4824\ : LocalMux
    port map (
            O => \N__21291\,
            I => \N__21288\
        );

    \I__4823\ : Span4Mux_v
    port map (
            O => \N__21288\,
            I => \N__21284\
        );

    \I__4822\ : InMux
    port map (
            O => \N__21287\,
            I => \N__21281\
        );

    \I__4821\ : Odrv4
    port map (
            O => \N__21284\,
            I => \ppm_encoder_1.N_303\
        );

    \I__4820\ : LocalMux
    port map (
            O => \N__21281\,
            I => \ppm_encoder_1.N_303\
        );

    \I__4819\ : CascadeMux
    port map (
            O => \N__21276\,
            I => \N__21273\
        );

    \I__4818\ : InMux
    port map (
            O => \N__21273\,
            I => \N__21268\
        );

    \I__4817\ : CascadeMux
    port map (
            O => \N__21272\,
            I => \N__21265\
        );

    \I__4816\ : CascadeMux
    port map (
            O => \N__21271\,
            I => \N__21262\
        );

    \I__4815\ : LocalMux
    port map (
            O => \N__21268\,
            I => \N__21259\
        );

    \I__4814\ : InMux
    port map (
            O => \N__21265\,
            I => \N__21256\
        );

    \I__4813\ : InMux
    port map (
            O => \N__21262\,
            I => \N__21253\
        );

    \I__4812\ : Span4Mux_h
    port map (
            O => \N__21259\,
            I => \N__21248\
        );

    \I__4811\ : LocalMux
    port map (
            O => \N__21256\,
            I => \N__21248\
        );

    \I__4810\ : LocalMux
    port map (
            O => \N__21253\,
            I => \N__21245\
        );

    \I__4809\ : Span4Mux_h
    port map (
            O => \N__21248\,
            I => \N__21242\
        );

    \I__4808\ : Span4Mux_h
    port map (
            O => \N__21245\,
            I => \N__21239\
        );

    \I__4807\ : Odrv4
    port map (
            O => \N__21242\,
            I => \ppm_encoder_1.init_pulsesZ0Z_16\
        );

    \I__4806\ : Odrv4
    port map (
            O => \N__21239\,
            I => \ppm_encoder_1.init_pulsesZ0Z_16\
        );

    \I__4805\ : InMux
    port map (
            O => \N__21234\,
            I => \N__21224\
        );

    \I__4804\ : InMux
    port map (
            O => \N__21233\,
            I => \N__21192\
        );

    \I__4803\ : InMux
    port map (
            O => \N__21232\,
            I => \N__21192\
        );

    \I__4802\ : InMux
    port map (
            O => \N__21231\,
            I => \N__21192\
        );

    \I__4801\ : InMux
    port map (
            O => \N__21230\,
            I => \N__21192\
        );

    \I__4800\ : InMux
    port map (
            O => \N__21229\,
            I => \N__21187\
        );

    \I__4799\ : InMux
    port map (
            O => \N__21228\,
            I => \N__21187\
        );

    \I__4798\ : CascadeMux
    port map (
            O => \N__21227\,
            I => \N__21184\
        );

    \I__4797\ : LocalMux
    port map (
            O => \N__21224\,
            I => \N__21181\
        );

    \I__4796\ : InMux
    port map (
            O => \N__21223\,
            I => \N__21178\
        );

    \I__4795\ : InMux
    port map (
            O => \N__21222\,
            I => \N__21173\
        );

    \I__4794\ : InMux
    port map (
            O => \N__21221\,
            I => \N__21173\
        );

    \I__4793\ : InMux
    port map (
            O => \N__21220\,
            I => \N__21170\
        );

    \I__4792\ : InMux
    port map (
            O => \N__21219\,
            I => \N__21164\
        );

    \I__4791\ : InMux
    port map (
            O => \N__21218\,
            I => \N__21155\
        );

    \I__4790\ : InMux
    port map (
            O => \N__21217\,
            I => \N__21155\
        );

    \I__4789\ : InMux
    port map (
            O => \N__21216\,
            I => \N__21155\
        );

    \I__4788\ : InMux
    port map (
            O => \N__21215\,
            I => \N__21155\
        );

    \I__4787\ : InMux
    port map (
            O => \N__21214\,
            I => \N__21146\
        );

    \I__4786\ : InMux
    port map (
            O => \N__21213\,
            I => \N__21146\
        );

    \I__4785\ : InMux
    port map (
            O => \N__21212\,
            I => \N__21146\
        );

    \I__4784\ : InMux
    port map (
            O => \N__21211\,
            I => \N__21146\
        );

    \I__4783\ : InMux
    port map (
            O => \N__21210\,
            I => \N__21140\
        );

    \I__4782\ : InMux
    port map (
            O => \N__21209\,
            I => \N__21140\
        );

    \I__4781\ : InMux
    port map (
            O => \N__21208\,
            I => \N__21131\
        );

    \I__4780\ : InMux
    port map (
            O => \N__21207\,
            I => \N__21131\
        );

    \I__4779\ : InMux
    port map (
            O => \N__21206\,
            I => \N__21131\
        );

    \I__4778\ : InMux
    port map (
            O => \N__21205\,
            I => \N__21131\
        );

    \I__4777\ : InMux
    port map (
            O => \N__21204\,
            I => \N__21123\
        );

    \I__4776\ : InMux
    port map (
            O => \N__21203\,
            I => \N__21123\
        );

    \I__4775\ : InMux
    port map (
            O => \N__21202\,
            I => \N__21123\
        );

    \I__4774\ : InMux
    port map (
            O => \N__21201\,
            I => \N__21120\
        );

    \I__4773\ : LocalMux
    port map (
            O => \N__21192\,
            I => \N__21115\
        );

    \I__4772\ : LocalMux
    port map (
            O => \N__21187\,
            I => \N__21115\
        );

    \I__4771\ : InMux
    port map (
            O => \N__21184\,
            I => \N__21112\
        );

    \I__4770\ : Span4Mux_h
    port map (
            O => \N__21181\,
            I => \N__21109\
        );

    \I__4769\ : LocalMux
    port map (
            O => \N__21178\,
            I => \N__21106\
        );

    \I__4768\ : LocalMux
    port map (
            O => \N__21173\,
            I => \N__21101\
        );

    \I__4767\ : LocalMux
    port map (
            O => \N__21170\,
            I => \N__21101\
        );

    \I__4766\ : CascadeMux
    port map (
            O => \N__21169\,
            I => \N__21094\
        );

    \I__4765\ : CascadeMux
    port map (
            O => \N__21168\,
            I => \N__21091\
        );

    \I__4764\ : InMux
    port map (
            O => \N__21167\,
            I => \N__21080\
        );

    \I__4763\ : LocalMux
    port map (
            O => \N__21164\,
            I => \N__21073\
        );

    \I__4762\ : LocalMux
    port map (
            O => \N__21155\,
            I => \N__21073\
        );

    \I__4761\ : LocalMux
    port map (
            O => \N__21146\,
            I => \N__21073\
        );

    \I__4760\ : InMux
    port map (
            O => \N__21145\,
            I => \N__21070\
        );

    \I__4759\ : LocalMux
    port map (
            O => \N__21140\,
            I => \N__21065\
        );

    \I__4758\ : LocalMux
    port map (
            O => \N__21131\,
            I => \N__21065\
        );

    \I__4757\ : CascadeMux
    port map (
            O => \N__21130\,
            I => \N__21057\
        );

    \I__4756\ : LocalMux
    port map (
            O => \N__21123\,
            I => \N__21044\
        );

    \I__4755\ : LocalMux
    port map (
            O => \N__21120\,
            I => \N__21044\
        );

    \I__4754\ : Span4Mux_v
    port map (
            O => \N__21115\,
            I => \N__21044\
        );

    \I__4753\ : LocalMux
    port map (
            O => \N__21112\,
            I => \N__21044\
        );

    \I__4752\ : Sp12to4
    port map (
            O => \N__21109\,
            I => \N__21041\
        );

    \I__4751\ : Span4Mux_v
    port map (
            O => \N__21106\,
            I => \N__21038\
        );

    \I__4750\ : Span4Mux_v
    port map (
            O => \N__21101\,
            I => \N__21035\
        );

    \I__4749\ : InMux
    port map (
            O => \N__21100\,
            I => \N__21032\
        );

    \I__4748\ : InMux
    port map (
            O => \N__21099\,
            I => \N__21021\
        );

    \I__4747\ : InMux
    port map (
            O => \N__21098\,
            I => \N__21021\
        );

    \I__4746\ : InMux
    port map (
            O => \N__21097\,
            I => \N__21021\
        );

    \I__4745\ : InMux
    port map (
            O => \N__21094\,
            I => \N__21021\
        );

    \I__4744\ : InMux
    port map (
            O => \N__21091\,
            I => \N__21021\
        );

    \I__4743\ : InMux
    port map (
            O => \N__21090\,
            I => \N__21010\
        );

    \I__4742\ : InMux
    port map (
            O => \N__21089\,
            I => \N__21010\
        );

    \I__4741\ : InMux
    port map (
            O => \N__21088\,
            I => \N__21010\
        );

    \I__4740\ : InMux
    port map (
            O => \N__21087\,
            I => \N__21010\
        );

    \I__4739\ : InMux
    port map (
            O => \N__21086\,
            I => \N__21010\
        );

    \I__4738\ : InMux
    port map (
            O => \N__21085\,
            I => \N__21005\
        );

    \I__4737\ : InMux
    port map (
            O => \N__21084\,
            I => \N__21005\
        );

    \I__4736\ : InMux
    port map (
            O => \N__21083\,
            I => \N__21002\
        );

    \I__4735\ : LocalMux
    port map (
            O => \N__21080\,
            I => \N__20993\
        );

    \I__4734\ : Span4Mux_v
    port map (
            O => \N__21073\,
            I => \N__20993\
        );

    \I__4733\ : LocalMux
    port map (
            O => \N__21070\,
            I => \N__20993\
        );

    \I__4732\ : Span4Mux_h
    port map (
            O => \N__21065\,
            I => \N__20993\
        );

    \I__4731\ : InMux
    port map (
            O => \N__21064\,
            I => \N__20984\
        );

    \I__4730\ : InMux
    port map (
            O => \N__21063\,
            I => \N__20984\
        );

    \I__4729\ : InMux
    port map (
            O => \N__21062\,
            I => \N__20984\
        );

    \I__4728\ : InMux
    port map (
            O => \N__21061\,
            I => \N__20984\
        );

    \I__4727\ : InMux
    port map (
            O => \N__21060\,
            I => \N__20979\
        );

    \I__4726\ : InMux
    port map (
            O => \N__21057\,
            I => \N__20979\
        );

    \I__4725\ : InMux
    port map (
            O => \N__21056\,
            I => \N__20970\
        );

    \I__4724\ : InMux
    port map (
            O => \N__21055\,
            I => \N__20970\
        );

    \I__4723\ : InMux
    port map (
            O => \N__21054\,
            I => \N__20970\
        );

    \I__4722\ : InMux
    port map (
            O => \N__21053\,
            I => \N__20970\
        );

    \I__4721\ : Odrv4
    port map (
            O => \N__21044\,
            I => \ppm_encoder_1.PPM_STATE_fast_RNICIABZ0Z_0\
        );

    \I__4720\ : Odrv12
    port map (
            O => \N__21041\,
            I => \ppm_encoder_1.PPM_STATE_fast_RNICIABZ0Z_0\
        );

    \I__4719\ : Odrv4
    port map (
            O => \N__21038\,
            I => \ppm_encoder_1.PPM_STATE_fast_RNICIABZ0Z_0\
        );

    \I__4718\ : Odrv4
    port map (
            O => \N__21035\,
            I => \ppm_encoder_1.PPM_STATE_fast_RNICIABZ0Z_0\
        );

    \I__4717\ : LocalMux
    port map (
            O => \N__21032\,
            I => \ppm_encoder_1.PPM_STATE_fast_RNICIABZ0Z_0\
        );

    \I__4716\ : LocalMux
    port map (
            O => \N__21021\,
            I => \ppm_encoder_1.PPM_STATE_fast_RNICIABZ0Z_0\
        );

    \I__4715\ : LocalMux
    port map (
            O => \N__21010\,
            I => \ppm_encoder_1.PPM_STATE_fast_RNICIABZ0Z_0\
        );

    \I__4714\ : LocalMux
    port map (
            O => \N__21005\,
            I => \ppm_encoder_1.PPM_STATE_fast_RNICIABZ0Z_0\
        );

    \I__4713\ : LocalMux
    port map (
            O => \N__21002\,
            I => \ppm_encoder_1.PPM_STATE_fast_RNICIABZ0Z_0\
        );

    \I__4712\ : Odrv4
    port map (
            O => \N__20993\,
            I => \ppm_encoder_1.PPM_STATE_fast_RNICIABZ0Z_0\
        );

    \I__4711\ : LocalMux
    port map (
            O => \N__20984\,
            I => \ppm_encoder_1.PPM_STATE_fast_RNICIABZ0Z_0\
        );

    \I__4710\ : LocalMux
    port map (
            O => \N__20979\,
            I => \ppm_encoder_1.PPM_STATE_fast_RNICIABZ0Z_0\
        );

    \I__4709\ : LocalMux
    port map (
            O => \N__20970\,
            I => \ppm_encoder_1.PPM_STATE_fast_RNICIABZ0Z_0\
        );

    \I__4708\ : IoInMux
    port map (
            O => \N__20943\,
            I => \N__20940\
        );

    \I__4707\ : LocalMux
    port map (
            O => \N__20940\,
            I => \N__20937\
        );

    \I__4706\ : Span12Mux_s6_v
    port map (
            O => \N__20937\,
            I => \N__20934\
        );

    \I__4705\ : Odrv12
    port map (
            O => \N__20934\,
            I => \ppm_encoder_1.N_238_i_0\
        );

    \I__4704\ : CascadeMux
    port map (
            O => \N__20931\,
            I => \N__20927\
        );

    \I__4703\ : InMux
    port map (
            O => \N__20930\,
            I => \N__20923\
        );

    \I__4702\ : InMux
    port map (
            O => \N__20927\,
            I => \N__20920\
        );

    \I__4701\ : CascadeMux
    port map (
            O => \N__20926\,
            I => \N__20917\
        );

    \I__4700\ : LocalMux
    port map (
            O => \N__20923\,
            I => \N__20914\
        );

    \I__4699\ : LocalMux
    port map (
            O => \N__20920\,
            I => \N__20911\
        );

    \I__4698\ : InMux
    port map (
            O => \N__20917\,
            I => \N__20908\
        );

    \I__4697\ : Span4Mux_h
    port map (
            O => \N__20914\,
            I => \N__20905\
        );

    \I__4696\ : Span4Mux_v
    port map (
            O => \N__20911\,
            I => \N__20902\
        );

    \I__4695\ : LocalMux
    port map (
            O => \N__20908\,
            I => \N__20899\
        );

    \I__4694\ : Span4Mux_v
    port map (
            O => \N__20905\,
            I => \N__20894\
        );

    \I__4693\ : Span4Mux_v
    port map (
            O => \N__20902\,
            I => \N__20894\
        );

    \I__4692\ : Odrv4
    port map (
            O => \N__20899\,
            I => \ppm_encoder_1.init_pulsesZ0Z_17\
        );

    \I__4691\ : Odrv4
    port map (
            O => \N__20894\,
            I => \ppm_encoder_1.init_pulsesZ0Z_17\
        );

    \I__4690\ : CascadeMux
    port map (
            O => \N__20889\,
            I => \N__20886\
        );

    \I__4689\ : InMux
    port map (
            O => \N__20886\,
            I => \N__20882\
        );

    \I__4688\ : InMux
    port map (
            O => \N__20885\,
            I => \N__20879\
        );

    \I__4687\ : LocalMux
    port map (
            O => \N__20882\,
            I => \N__20876\
        );

    \I__4686\ : LocalMux
    port map (
            O => \N__20879\,
            I => \N__20872\
        );

    \I__4685\ : Span4Mux_h
    port map (
            O => \N__20876\,
            I => \N__20869\
        );

    \I__4684\ : InMux
    port map (
            O => \N__20875\,
            I => \N__20866\
        );

    \I__4683\ : Span4Mux_v
    port map (
            O => \N__20872\,
            I => \N__20863\
        );

    \I__4682\ : Odrv4
    port map (
            O => \N__20869\,
            I => \ppm_encoder_1.init_pulsesZ0Z_18\
        );

    \I__4681\ : LocalMux
    port map (
            O => \N__20866\,
            I => \ppm_encoder_1.init_pulsesZ0Z_18\
        );

    \I__4680\ : Odrv4
    port map (
            O => \N__20863\,
            I => \ppm_encoder_1.init_pulsesZ0Z_18\
        );

    \I__4679\ : InMux
    port map (
            O => \N__20856\,
            I => \bfn_11_25_0_\
        );

    \I__4678\ : InMux
    port map (
            O => \N__20853\,
            I => \ppm_encoder_1.un1_counter_13_cry_8\
        );

    \I__4677\ : InMux
    port map (
            O => \N__20850\,
            I => \ppm_encoder_1.un1_counter_13_cry_9\
        );

    \I__4676\ : InMux
    port map (
            O => \N__20847\,
            I => \ppm_encoder_1.un1_counter_13_cry_10\
        );

    \I__4675\ : InMux
    port map (
            O => \N__20844\,
            I => \ppm_encoder_1.un1_counter_13_cry_11\
        );

    \I__4674\ : InMux
    port map (
            O => \N__20841\,
            I => \ppm_encoder_1.un1_counter_13_cry_12\
        );

    \I__4673\ : InMux
    port map (
            O => \N__20838\,
            I => \ppm_encoder_1.un1_counter_13_cry_13\
        );

    \I__4672\ : InMux
    port map (
            O => \N__20835\,
            I => \ppm_encoder_1.un1_counter_13_cry_14\
        );

    \I__4671\ : InMux
    port map (
            O => \N__20832\,
            I => \bfn_11_26_0_\
        );

    \I__4670\ : InMux
    port map (
            O => \N__20829\,
            I => \N__20825\
        );

    \I__4669\ : InMux
    port map (
            O => \N__20828\,
            I => \N__20822\
        );

    \I__4668\ : LocalMux
    port map (
            O => \N__20825\,
            I => \N__20817\
        );

    \I__4667\ : LocalMux
    port map (
            O => \N__20822\,
            I => \N__20817\
        );

    \I__4666\ : Span4Mux_v
    port map (
            O => \N__20817\,
            I => \N__20812\
        );

    \I__4665\ : InMux
    port map (
            O => \N__20816\,
            I => \N__20809\
        );

    \I__4664\ : CascadeMux
    port map (
            O => \N__20815\,
            I => \N__20806\
        );

    \I__4663\ : Span4Mux_h
    port map (
            O => \N__20812\,
            I => \N__20801\
        );

    \I__4662\ : LocalMux
    port map (
            O => \N__20809\,
            I => \N__20801\
        );

    \I__4661\ : InMux
    port map (
            O => \N__20806\,
            I => \N__20798\
        );

    \I__4660\ : Odrv4
    port map (
            O => \N__20801\,
            I => \ppm_encoder_1.N_443\
        );

    \I__4659\ : LocalMux
    port map (
            O => \N__20798\,
            I => \ppm_encoder_1.N_443\
        );

    \I__4658\ : CascadeMux
    port map (
            O => \N__20793\,
            I => \N__20790\
        );

    \I__4657\ : InMux
    port map (
            O => \N__20790\,
            I => \N__20787\
        );

    \I__4656\ : LocalMux
    port map (
            O => \N__20787\,
            I => \N__20784\
        );

    \I__4655\ : Span12Mux_s8_v
    port map (
            O => \N__20784\,
            I => \N__20781\
        );

    \I__4654\ : Odrv12
    port map (
            O => \N__20781\,
            I => \ppm_encoder_1.pulses2count_9_0_2_1\
        );

    \I__4653\ : InMux
    port map (
            O => \N__20778\,
            I => \N__20772\
        );

    \I__4652\ : InMux
    port map (
            O => \N__20777\,
            I => \N__20772\
        );

    \I__4651\ : LocalMux
    port map (
            O => \N__20772\,
            I => \N__20767\
        );

    \I__4650\ : InMux
    port map (
            O => \N__20771\,
            I => \N__20762\
        );

    \I__4649\ : InMux
    port map (
            O => \N__20770\,
            I => \N__20762\
        );

    \I__4648\ : Odrv4
    port map (
            O => \N__20767\,
            I => \ppm_encoder_1.throttleZ0Z_1\
        );

    \I__4647\ : LocalMux
    port map (
            O => \N__20762\,
            I => \ppm_encoder_1.throttleZ0Z_1\
        );

    \I__4646\ : InMux
    port map (
            O => \N__20757\,
            I => \ppm_encoder_1.un1_counter_13_cry_0\
        );

    \I__4645\ : InMux
    port map (
            O => \N__20754\,
            I => \N__20749\
        );

    \I__4644\ : InMux
    port map (
            O => \N__20753\,
            I => \N__20746\
        );

    \I__4643\ : InMux
    port map (
            O => \N__20752\,
            I => \N__20743\
        );

    \I__4642\ : LocalMux
    port map (
            O => \N__20749\,
            I => \ppm_encoder_1.counterZ0Z_2\
        );

    \I__4641\ : LocalMux
    port map (
            O => \N__20746\,
            I => \ppm_encoder_1.counterZ0Z_2\
        );

    \I__4640\ : LocalMux
    port map (
            O => \N__20743\,
            I => \ppm_encoder_1.counterZ0Z_2\
        );

    \I__4639\ : InMux
    port map (
            O => \N__20736\,
            I => \ppm_encoder_1.un1_counter_13_cry_1\
        );

    \I__4638\ : InMux
    port map (
            O => \N__20733\,
            I => \N__20728\
        );

    \I__4637\ : InMux
    port map (
            O => \N__20732\,
            I => \N__20725\
        );

    \I__4636\ : InMux
    port map (
            O => \N__20731\,
            I => \N__20722\
        );

    \I__4635\ : LocalMux
    port map (
            O => \N__20728\,
            I => \ppm_encoder_1.counterZ0Z_3\
        );

    \I__4634\ : LocalMux
    port map (
            O => \N__20725\,
            I => \ppm_encoder_1.counterZ0Z_3\
        );

    \I__4633\ : LocalMux
    port map (
            O => \N__20722\,
            I => \ppm_encoder_1.counterZ0Z_3\
        );

    \I__4632\ : InMux
    port map (
            O => \N__20715\,
            I => \ppm_encoder_1.un1_counter_13_cry_2\
        );

    \I__4631\ : InMux
    port map (
            O => \N__20712\,
            I => \ppm_encoder_1.un1_counter_13_cry_3\
        );

    \I__4630\ : InMux
    port map (
            O => \N__20709\,
            I => \ppm_encoder_1.un1_counter_13_cry_4\
        );

    \I__4629\ : InMux
    port map (
            O => \N__20706\,
            I => \ppm_encoder_1.un1_counter_13_cry_5\
        );

    \I__4628\ : InMux
    port map (
            O => \N__20703\,
            I => \ppm_encoder_1.un1_counter_13_cry_6\
        );

    \I__4627\ : InMux
    port map (
            O => \N__20700\,
            I => \N__20697\
        );

    \I__4626\ : LocalMux
    port map (
            O => \N__20697\,
            I => \N__20694\
        );

    \I__4625\ : Span12Mux_h
    port map (
            O => \N__20694\,
            I => \N__20691\
        );

    \I__4624\ : Odrv12
    port map (
            O => \N__20691\,
            I => \ppm_encoder_1.N_369\
        );

    \I__4623\ : CascadeMux
    port map (
            O => \N__20688\,
            I => \ppm_encoder_1.N_371_cascade_\
        );

    \I__4622\ : InMux
    port map (
            O => \N__20685\,
            I => \N__20682\
        );

    \I__4621\ : LocalMux
    port map (
            O => \N__20682\,
            I => \N__20679\
        );

    \I__4620\ : Span4Mux_v
    port map (
            O => \N__20679\,
            I => \N__20676\
        );

    \I__4619\ : Span4Mux_v
    port map (
            O => \N__20676\,
            I => \N__20672\
        );

    \I__4618\ : InMux
    port map (
            O => \N__20675\,
            I => \N__20669\
        );

    \I__4617\ : Odrv4
    port map (
            O => \N__20672\,
            I => \ppm_encoder_1.rudderZ0Z_4\
        );

    \I__4616\ : LocalMux
    port map (
            O => \N__20669\,
            I => \ppm_encoder_1.rudderZ0Z_4\
        );

    \I__4615\ : InMux
    port map (
            O => \N__20664\,
            I => \N__20660\
        );

    \I__4614\ : CascadeMux
    port map (
            O => \N__20663\,
            I => \N__20656\
        );

    \I__4613\ : LocalMux
    port map (
            O => \N__20660\,
            I => \N__20653\
        );

    \I__4612\ : InMux
    port map (
            O => \N__20659\,
            I => \N__20650\
        );

    \I__4611\ : InMux
    port map (
            O => \N__20656\,
            I => \N__20647\
        );

    \I__4610\ : Span4Mux_v
    port map (
            O => \N__20653\,
            I => \N__20644\
        );

    \I__4609\ : LocalMux
    port map (
            O => \N__20650\,
            I => \N__20641\
        );

    \I__4608\ : LocalMux
    port map (
            O => \N__20647\,
            I => \N__20638\
        );

    \I__4607\ : Span4Mux_h
    port map (
            O => \N__20644\,
            I => \N__20635\
        );

    \I__4606\ : Span4Mux_h
    port map (
            O => \N__20641\,
            I => \N__20632\
        );

    \I__4605\ : Odrv4
    port map (
            O => \N__20638\,
            I => \ppm_encoder_1.rudderZ0Z_13\
        );

    \I__4604\ : Odrv4
    port map (
            O => \N__20635\,
            I => \ppm_encoder_1.rudderZ0Z_13\
        );

    \I__4603\ : Odrv4
    port map (
            O => \N__20632\,
            I => \ppm_encoder_1.rudderZ0Z_13\
        );

    \I__4602\ : InMux
    port map (
            O => \N__20625\,
            I => \N__20622\
        );

    \I__4601\ : LocalMux
    port map (
            O => \N__20622\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_15\
        );

    \I__4600\ : InMux
    port map (
            O => \N__20619\,
            I => \N__20616\
        );

    \I__4599\ : LocalMux
    port map (
            O => \N__20616\,
            I => \N__20611\
        );

    \I__4598\ : InMux
    port map (
            O => \N__20615\,
            I => \N__20608\
        );

    \I__4597\ : InMux
    port map (
            O => \N__20614\,
            I => \N__20605\
        );

    \I__4596\ : Span4Mux_v
    port map (
            O => \N__20611\,
            I => \N__20602\
        );

    \I__4595\ : LocalMux
    port map (
            O => \N__20608\,
            I => \N__20599\
        );

    \I__4594\ : LocalMux
    port map (
            O => \N__20605\,
            I => \ppm_encoder_1.throttleZ0Z_2\
        );

    \I__4593\ : Odrv4
    port map (
            O => \N__20602\,
            I => \ppm_encoder_1.throttleZ0Z_2\
        );

    \I__4592\ : Odrv12
    port map (
            O => \N__20599\,
            I => \ppm_encoder_1.throttleZ0Z_2\
        );

    \I__4591\ : InMux
    port map (
            O => \N__20592\,
            I => \N__20588\
        );

    \I__4590\ : CascadeMux
    port map (
            O => \N__20591\,
            I => \N__20583\
        );

    \I__4589\ : LocalMux
    port map (
            O => \N__20588\,
            I => \N__20580\
        );

    \I__4588\ : InMux
    port map (
            O => \N__20587\,
            I => \N__20577\
        );

    \I__4587\ : InMux
    port map (
            O => \N__20586\,
            I => \N__20574\
        );

    \I__4586\ : InMux
    port map (
            O => \N__20583\,
            I => \N__20571\
        );

    \I__4585\ : Span4Mux_h
    port map (
            O => \N__20580\,
            I => \N__20562\
        );

    \I__4584\ : LocalMux
    port map (
            O => \N__20577\,
            I => \N__20562\
        );

    \I__4583\ : LocalMux
    port map (
            O => \N__20574\,
            I => \N__20562\
        );

    \I__4582\ : LocalMux
    port map (
            O => \N__20571\,
            I => \N__20562\
        );

    \I__4581\ : Span4Mux_v
    port map (
            O => \N__20562\,
            I => \N__20559\
        );

    \I__4580\ : Odrv4
    port map (
            O => \N__20559\,
            I => \ppm_encoder_1.init_pulsesZ0Z_3\
        );

    \I__4579\ : InMux
    port map (
            O => \N__20556\,
            I => \N__20553\
        );

    \I__4578\ : LocalMux
    port map (
            O => \N__20553\,
            I => \N__20550\
        );

    \I__4577\ : Odrv4
    port map (
            O => \N__20550\,
            I => \ppm_encoder_1.N_360\
        );

    \I__4576\ : CascadeMux
    port map (
            O => \N__20547\,
            I => \N__20544\
        );

    \I__4575\ : InMux
    port map (
            O => \N__20544\,
            I => \N__20541\
        );

    \I__4574\ : LocalMux
    port map (
            O => \N__20541\,
            I => \N__20536\
        );

    \I__4573\ : InMux
    port map (
            O => \N__20540\,
            I => \N__20533\
        );

    \I__4572\ : CascadeMux
    port map (
            O => \N__20539\,
            I => \N__20528\
        );

    \I__4571\ : Span4Mux_v
    port map (
            O => \N__20536\,
            I => \N__20525\
        );

    \I__4570\ : LocalMux
    port map (
            O => \N__20533\,
            I => \N__20522\
        );

    \I__4569\ : InMux
    port map (
            O => \N__20532\,
            I => \N__20515\
        );

    \I__4568\ : InMux
    port map (
            O => \N__20531\,
            I => \N__20515\
        );

    \I__4567\ : InMux
    port map (
            O => \N__20528\,
            I => \N__20515\
        );

    \I__4566\ : Span4Mux_h
    port map (
            O => \N__20525\,
            I => \N__20512\
        );

    \I__4565\ : Span4Mux_h
    port map (
            O => \N__20522\,
            I => \N__20507\
        );

    \I__4564\ : LocalMux
    port map (
            O => \N__20515\,
            I => \N__20507\
        );

    \I__4563\ : Odrv4
    port map (
            O => \N__20512\,
            I => \ppm_encoder_1.init_pulsesZ0Z_2\
        );

    \I__4562\ : Odrv4
    port map (
            O => \N__20507\,
            I => \ppm_encoder_1.init_pulsesZ0Z_2\
        );

    \I__4561\ : CascadeMux
    port map (
            O => \N__20502\,
            I => \N__20498\
        );

    \I__4560\ : InMux
    port map (
            O => \N__20501\,
            I => \N__20495\
        );

    \I__4559\ : InMux
    port map (
            O => \N__20498\,
            I => \N__20492\
        );

    \I__4558\ : LocalMux
    port map (
            O => \N__20495\,
            I => \ppm_encoder_1.pulses2count_9_0_0_3\
        );

    \I__4557\ : LocalMux
    port map (
            O => \N__20492\,
            I => \ppm_encoder_1.pulses2count_9_0_0_3\
        );

    \I__4556\ : InMux
    port map (
            O => \N__20487\,
            I => \N__20484\
        );

    \I__4555\ : LocalMux
    port map (
            O => \N__20484\,
            I => \ppm_encoder_1.pulses2countZ0Z_2\
        );

    \I__4554\ : CascadeMux
    port map (
            O => \N__20481\,
            I => \N__20478\
        );

    \I__4553\ : InMux
    port map (
            O => \N__20478\,
            I => \N__20475\
        );

    \I__4552\ : LocalMux
    port map (
            O => \N__20475\,
            I => \ppm_encoder_1.pulses2countZ0Z_3\
        );

    \I__4551\ : InMux
    port map (
            O => \N__20472\,
            I => \N__20469\
        );

    \I__4550\ : LocalMux
    port map (
            O => \N__20469\,
            I => \ppm_encoder_1.N_365\
        );

    \I__4549\ : InMux
    port map (
            O => \N__20466\,
            I => \N__20463\
        );

    \I__4548\ : LocalMux
    port map (
            O => \N__20463\,
            I => \ppm_encoder_1.init_pulses_RNILB4MZ0Z_0\
        );

    \I__4547\ : InMux
    port map (
            O => \N__20460\,
            I => \N__20455\
        );

    \I__4546\ : InMux
    port map (
            O => \N__20459\,
            I => \N__20450\
        );

    \I__4545\ : InMux
    port map (
            O => \N__20458\,
            I => \N__20450\
        );

    \I__4544\ : LocalMux
    port map (
            O => \N__20455\,
            I => \N__20444\
        );

    \I__4543\ : LocalMux
    port map (
            O => \N__20450\,
            I => \N__20444\
        );

    \I__4542\ : InMux
    port map (
            O => \N__20449\,
            I => \N__20441\
        );

    \I__4541\ : Span4Mux_h
    port map (
            O => \N__20444\,
            I => \N__20435\
        );

    \I__4540\ : LocalMux
    port map (
            O => \N__20441\,
            I => \N__20435\
        );

    \I__4539\ : CascadeMux
    port map (
            O => \N__20440\,
            I => \N__20432\
        );

    \I__4538\ : Span4Mux_v
    port map (
            O => \N__20435\,
            I => \N__20429\
        );

    \I__4537\ : InMux
    port map (
            O => \N__20432\,
            I => \N__20426\
        );

    \I__4536\ : Odrv4
    port map (
            O => \N__20429\,
            I => \ppm_encoder_1.N_247_i_i\
        );

    \I__4535\ : LocalMux
    port map (
            O => \N__20426\,
            I => \ppm_encoder_1.N_247_i_i\
        );

    \I__4534\ : CascadeMux
    port map (
            O => \N__20421\,
            I => \N__20415\
        );

    \I__4533\ : InMux
    port map (
            O => \N__20420\,
            I => \N__20409\
        );

    \I__4532\ : InMux
    port map (
            O => \N__20419\,
            I => \N__20409\
        );

    \I__4531\ : InMux
    port map (
            O => \N__20418\,
            I => \N__20403\
        );

    \I__4530\ : InMux
    port map (
            O => \N__20415\,
            I => \N__20400\
        );

    \I__4529\ : InMux
    port map (
            O => \N__20414\,
            I => \N__20392\
        );

    \I__4528\ : LocalMux
    port map (
            O => \N__20409\,
            I => \N__20388\
        );

    \I__4527\ : InMux
    port map (
            O => \N__20408\,
            I => \N__20381\
        );

    \I__4526\ : InMux
    port map (
            O => \N__20407\,
            I => \N__20381\
        );

    \I__4525\ : InMux
    port map (
            O => \N__20406\,
            I => \N__20381\
        );

    \I__4524\ : LocalMux
    port map (
            O => \N__20403\,
            I => \N__20376\
        );

    \I__4523\ : LocalMux
    port map (
            O => \N__20400\,
            I => \N__20376\
        );

    \I__4522\ : InMux
    port map (
            O => \N__20399\,
            I => \N__20371\
        );

    \I__4521\ : InMux
    port map (
            O => \N__20398\,
            I => \N__20371\
        );

    \I__4520\ : InMux
    port map (
            O => \N__20397\,
            I => \N__20368\
        );

    \I__4519\ : InMux
    port map (
            O => \N__20396\,
            I => \N__20363\
        );

    \I__4518\ : InMux
    port map (
            O => \N__20395\,
            I => \N__20363\
        );

    \I__4517\ : LocalMux
    port map (
            O => \N__20392\,
            I => \N__20359\
        );

    \I__4516\ : InMux
    port map (
            O => \N__20391\,
            I => \N__20356\
        );

    \I__4515\ : Span4Mux_v
    port map (
            O => \N__20388\,
            I => \N__20351\
        );

    \I__4514\ : LocalMux
    port map (
            O => \N__20381\,
            I => \N__20351\
        );

    \I__4513\ : Span4Mux_v
    port map (
            O => \N__20376\,
            I => \N__20337\
        );

    \I__4512\ : LocalMux
    port map (
            O => \N__20371\,
            I => \N__20337\
        );

    \I__4511\ : LocalMux
    port map (
            O => \N__20368\,
            I => \N__20334\
        );

    \I__4510\ : LocalMux
    port map (
            O => \N__20363\,
            I => \N__20331\
        );

    \I__4509\ : InMux
    port map (
            O => \N__20362\,
            I => \N__20328\
        );

    \I__4508\ : Span4Mux_v
    port map (
            O => \N__20359\,
            I => \N__20321\
        );

    \I__4507\ : LocalMux
    port map (
            O => \N__20356\,
            I => \N__20321\
        );

    \I__4506\ : Span4Mux_v
    port map (
            O => \N__20351\,
            I => \N__20321\
        );

    \I__4505\ : InMux
    port map (
            O => \N__20350\,
            I => \N__20316\
        );

    \I__4504\ : InMux
    port map (
            O => \N__20349\,
            I => \N__20316\
        );

    \I__4503\ : InMux
    port map (
            O => \N__20348\,
            I => \N__20311\
        );

    \I__4502\ : InMux
    port map (
            O => \N__20347\,
            I => \N__20311\
        );

    \I__4501\ : InMux
    port map (
            O => \N__20346\,
            I => \N__20302\
        );

    \I__4500\ : InMux
    port map (
            O => \N__20345\,
            I => \N__20302\
        );

    \I__4499\ : InMux
    port map (
            O => \N__20344\,
            I => \N__20302\
        );

    \I__4498\ : InMux
    port map (
            O => \N__20343\,
            I => \N__20302\
        );

    \I__4497\ : InMux
    port map (
            O => \N__20342\,
            I => \N__20299\
        );

    \I__4496\ : Span4Mux_h
    port map (
            O => \N__20337\,
            I => \N__20294\
        );

    \I__4495\ : Span4Mux_v
    port map (
            O => \N__20334\,
            I => \N__20294\
        );

    \I__4494\ : Span4Mux_h
    port map (
            O => \N__20331\,
            I => \N__20287\
        );

    \I__4493\ : LocalMux
    port map (
            O => \N__20328\,
            I => \N__20287\
        );

    \I__4492\ : Span4Mux_h
    port map (
            O => \N__20321\,
            I => \N__20287\
        );

    \I__4491\ : LocalMux
    port map (
            O => \N__20316\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z2\
        );

    \I__4490\ : LocalMux
    port map (
            O => \N__20311\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z2\
        );

    \I__4489\ : LocalMux
    port map (
            O => \N__20302\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z2\
        );

    \I__4488\ : LocalMux
    port map (
            O => \N__20299\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z2\
        );

    \I__4487\ : Odrv4
    port map (
            O => \N__20294\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z2\
        );

    \I__4486\ : Odrv4
    port map (
            O => \N__20287\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z2\
        );

    \I__4485\ : CascadeMux
    port map (
            O => \N__20274\,
            I => \N__20269\
        );

    \I__4484\ : CascadeMux
    port map (
            O => \N__20273\,
            I => \N__20266\
        );

    \I__4483\ : InMux
    port map (
            O => \N__20272\,
            I => \N__20263\
        );

    \I__4482\ : InMux
    port map (
            O => \N__20269\,
            I => \N__20258\
        );

    \I__4481\ : InMux
    port map (
            O => \N__20266\,
            I => \N__20258\
        );

    \I__4480\ : LocalMux
    port map (
            O => \N__20263\,
            I => \N__20250\
        );

    \I__4479\ : LocalMux
    port map (
            O => \N__20258\,
            I => \N__20250\
        );

    \I__4478\ : InMux
    port map (
            O => \N__20257\,
            I => \N__20247\
        );

    \I__4477\ : InMux
    port map (
            O => \N__20256\,
            I => \N__20244\
        );

    \I__4476\ : InMux
    port map (
            O => \N__20255\,
            I => \N__20237\
        );

    \I__4475\ : Span4Mux_v
    port map (
            O => \N__20250\,
            I => \N__20232\
        );

    \I__4474\ : LocalMux
    port map (
            O => \N__20247\,
            I => \N__20229\
        );

    \I__4473\ : LocalMux
    port map (
            O => \N__20244\,
            I => \N__20226\
        );

    \I__4472\ : InMux
    port map (
            O => \N__20243\,
            I => \N__20223\
        );

    \I__4471\ : InMux
    port map (
            O => \N__20242\,
            I => \N__20219\
        );

    \I__4470\ : InMux
    port map (
            O => \N__20241\,
            I => \N__20214\
        );

    \I__4469\ : InMux
    port map (
            O => \N__20240\,
            I => \N__20211\
        );

    \I__4468\ : LocalMux
    port map (
            O => \N__20237\,
            I => \N__20208\
        );

    \I__4467\ : InMux
    port map (
            O => \N__20236\,
            I => \N__20203\
        );

    \I__4466\ : InMux
    port map (
            O => \N__20235\,
            I => \N__20203\
        );

    \I__4465\ : Span4Mux_h
    port map (
            O => \N__20232\,
            I => \N__20200\
        );

    \I__4464\ : Span4Mux_h
    port map (
            O => \N__20229\,
            I => \N__20193\
        );

    \I__4463\ : Span4Mux_h
    port map (
            O => \N__20226\,
            I => \N__20193\
        );

    \I__4462\ : LocalMux
    port map (
            O => \N__20223\,
            I => \N__20193\
        );

    \I__4461\ : InMux
    port map (
            O => \N__20222\,
            I => \N__20190\
        );

    \I__4460\ : LocalMux
    port map (
            O => \N__20219\,
            I => \N__20187\
        );

    \I__4459\ : InMux
    port map (
            O => \N__20218\,
            I => \N__20182\
        );

    \I__4458\ : InMux
    port map (
            O => \N__20217\,
            I => \N__20182\
        );

    \I__4457\ : LocalMux
    port map (
            O => \N__20214\,
            I => \N__20177\
        );

    \I__4456\ : LocalMux
    port map (
            O => \N__20211\,
            I => \N__20177\
        );

    \I__4455\ : Odrv4
    port map (
            O => \N__20208\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z2\
        );

    \I__4454\ : LocalMux
    port map (
            O => \N__20203\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z2\
        );

    \I__4453\ : Odrv4
    port map (
            O => \N__20200\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z2\
        );

    \I__4452\ : Odrv4
    port map (
            O => \N__20193\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z2\
        );

    \I__4451\ : LocalMux
    port map (
            O => \N__20190\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z2\
        );

    \I__4450\ : Odrv12
    port map (
            O => \N__20187\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z2\
        );

    \I__4449\ : LocalMux
    port map (
            O => \N__20182\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z2\
        );

    \I__4448\ : Odrv4
    port map (
            O => \N__20177\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z2\
        );

    \I__4447\ : InMux
    port map (
            O => \N__20160\,
            I => \N__20152\
        );

    \I__4446\ : InMux
    port map (
            O => \N__20159\,
            I => \N__20152\
        );

    \I__4445\ : InMux
    port map (
            O => \N__20158\,
            I => \N__20147\
        );

    \I__4444\ : InMux
    port map (
            O => \N__20157\,
            I => \N__20144\
        );

    \I__4443\ : LocalMux
    port map (
            O => \N__20152\,
            I => \N__20140\
        );

    \I__4442\ : InMux
    port map (
            O => \N__20151\,
            I => \N__20137\
        );

    \I__4441\ : InMux
    port map (
            O => \N__20150\,
            I => \N__20134\
        );

    \I__4440\ : LocalMux
    port map (
            O => \N__20147\,
            I => \N__20129\
        );

    \I__4439\ : LocalMux
    port map (
            O => \N__20144\,
            I => \N__20124\
        );

    \I__4438\ : InMux
    port map (
            O => \N__20143\,
            I => \N__20121\
        );

    \I__4437\ : Span4Mux_h
    port map (
            O => \N__20140\,
            I => \N__20116\
        );

    \I__4436\ : LocalMux
    port map (
            O => \N__20137\,
            I => \N__20110\
        );

    \I__4435\ : LocalMux
    port map (
            O => \N__20134\,
            I => \N__20110\
        );

    \I__4434\ : InMux
    port map (
            O => \N__20133\,
            I => \N__20105\
        );

    \I__4433\ : InMux
    port map (
            O => \N__20132\,
            I => \N__20105\
        );

    \I__4432\ : Span4Mux_h
    port map (
            O => \N__20129\,
            I => \N__20100\
        );

    \I__4431\ : InMux
    port map (
            O => \N__20128\,
            I => \N__20097\
        );

    \I__4430\ : InMux
    port map (
            O => \N__20127\,
            I => \N__20094\
        );

    \I__4429\ : Span4Mux_h
    port map (
            O => \N__20124\,
            I => \N__20091\
        );

    \I__4428\ : LocalMux
    port map (
            O => \N__20121\,
            I => \N__20088\
        );

    \I__4427\ : InMux
    port map (
            O => \N__20120\,
            I => \N__20083\
        );

    \I__4426\ : InMux
    port map (
            O => \N__20119\,
            I => \N__20083\
        );

    \I__4425\ : Span4Mux_v
    port map (
            O => \N__20116\,
            I => \N__20080\
        );

    \I__4424\ : InMux
    port map (
            O => \N__20115\,
            I => \N__20077\
        );

    \I__4423\ : Span4Mux_h
    port map (
            O => \N__20110\,
            I => \N__20072\
        );

    \I__4422\ : LocalMux
    port map (
            O => \N__20105\,
            I => \N__20072\
        );

    \I__4421\ : InMux
    port map (
            O => \N__20104\,
            I => \N__20067\
        );

    \I__4420\ : InMux
    port map (
            O => \N__20103\,
            I => \N__20067\
        );

    \I__4419\ : Span4Mux_v
    port map (
            O => \N__20100\,
            I => \N__20060\
        );

    \I__4418\ : LocalMux
    port map (
            O => \N__20097\,
            I => \N__20060\
        );

    \I__4417\ : LocalMux
    port map (
            O => \N__20094\,
            I => \N__20060\
        );

    \I__4416\ : Odrv4
    port map (
            O => \N__20091\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z2\
        );

    \I__4415\ : Odrv4
    port map (
            O => \N__20088\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z2\
        );

    \I__4414\ : LocalMux
    port map (
            O => \N__20083\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z2\
        );

    \I__4413\ : Odrv4
    port map (
            O => \N__20080\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z2\
        );

    \I__4412\ : LocalMux
    port map (
            O => \N__20077\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z2\
        );

    \I__4411\ : Odrv4
    port map (
            O => \N__20072\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z2\
        );

    \I__4410\ : LocalMux
    port map (
            O => \N__20067\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z2\
        );

    \I__4409\ : Odrv4
    port map (
            O => \N__20060\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z2\
        );

    \I__4408\ : CascadeMux
    port map (
            O => \N__20043\,
            I => \N__20040\
        );

    \I__4407\ : InMux
    port map (
            O => \N__20040\,
            I => \N__20036\
        );

    \I__4406\ : CascadeMux
    port map (
            O => \N__20039\,
            I => \N__20033\
        );

    \I__4405\ : LocalMux
    port map (
            O => \N__20036\,
            I => \N__20029\
        );

    \I__4404\ : InMux
    port map (
            O => \N__20033\,
            I => \N__20026\
        );

    \I__4403\ : InMux
    port map (
            O => \N__20032\,
            I => \N__20023\
        );

    \I__4402\ : Span4Mux_v
    port map (
            O => \N__20029\,
            I => \N__20018\
        );

    \I__4401\ : LocalMux
    port map (
            O => \N__20026\,
            I => \N__20018\
        );

    \I__4400\ : LocalMux
    port map (
            O => \N__20023\,
            I => \N__20015\
        );

    \I__4399\ : Span4Mux_h
    port map (
            O => \N__20018\,
            I => \N__20011\
        );

    \I__4398\ : Span4Mux_h
    port map (
            O => \N__20015\,
            I => \N__20008\
        );

    \I__4397\ : InMux
    port map (
            O => \N__20014\,
            I => \N__20005\
        );

    \I__4396\ : Span4Mux_v
    port map (
            O => \N__20011\,
            I => \N__20002\
        );

    \I__4395\ : Odrv4
    port map (
            O => \N__20008\,
            I => \ppm_encoder_1.init_pulsesZ0Z_11\
        );

    \I__4394\ : LocalMux
    port map (
            O => \N__20005\,
            I => \ppm_encoder_1.init_pulsesZ0Z_11\
        );

    \I__4393\ : Odrv4
    port map (
            O => \N__20002\,
            I => \ppm_encoder_1.init_pulsesZ0Z_11\
        );

    \I__4392\ : CascadeMux
    port map (
            O => \N__19995\,
            I => \ppm_encoder_1.N_441_cascade_\
        );

    \I__4391\ : InMux
    port map (
            O => \N__19992\,
            I => \N__19989\
        );

    \I__4390\ : LocalMux
    port map (
            O => \N__19989\,
            I => \N__19985\
        );

    \I__4389\ : CascadeMux
    port map (
            O => \N__19988\,
            I => \N__19981\
        );

    \I__4388\ : Span4Mux_h
    port map (
            O => \N__19985\,
            I => \N__19978\
        );

    \I__4387\ : InMux
    port map (
            O => \N__19984\,
            I => \N__19973\
        );

    \I__4386\ : InMux
    port map (
            O => \N__19981\,
            I => \N__19973\
        );

    \I__4385\ : Odrv4
    port map (
            O => \N__19978\,
            I => \ppm_encoder_1.throttleZ0Z_11\
        );

    \I__4384\ : LocalMux
    port map (
            O => \N__19973\,
            I => \ppm_encoder_1.throttleZ0Z_11\
        );

    \I__4383\ : InMux
    port map (
            O => \N__19968\,
            I => \N__19965\
        );

    \I__4382\ : LocalMux
    port map (
            O => \N__19965\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_18\
        );

    \I__4381\ : InMux
    port map (
            O => \N__19962\,
            I => \N__19959\
        );

    \I__4380\ : LocalMux
    port map (
            O => \N__19959\,
            I => \N__19955\
        );

    \I__4379\ : CascadeMux
    port map (
            O => \N__19958\,
            I => \N__19951\
        );

    \I__4378\ : Span4Mux_h
    port map (
            O => \N__19955\,
            I => \N__19948\
        );

    \I__4377\ : InMux
    port map (
            O => \N__19954\,
            I => \N__19945\
        );

    \I__4376\ : InMux
    port map (
            O => \N__19951\,
            I => \N__19942\
        );

    \I__4375\ : Span4Mux_h
    port map (
            O => \N__19948\,
            I => \N__19937\
        );

    \I__4374\ : LocalMux
    port map (
            O => \N__19945\,
            I => \N__19937\
        );

    \I__4373\ : LocalMux
    port map (
            O => \N__19942\,
            I => \ppm_encoder_1.throttleZ0Z_10\
        );

    \I__4372\ : Odrv4
    port map (
            O => \N__19937\,
            I => \ppm_encoder_1.throttleZ0Z_10\
        );

    \I__4371\ : InMux
    port map (
            O => \N__19932\,
            I => \N__19928\
        );

    \I__4370\ : CascadeMux
    port map (
            O => \N__19931\,
            I => \N__19924\
        );

    \I__4369\ : LocalMux
    port map (
            O => \N__19928\,
            I => \N__19921\
        );

    \I__4368\ : InMux
    port map (
            O => \N__19927\,
            I => \N__19918\
        );

    \I__4367\ : InMux
    port map (
            O => \N__19924\,
            I => \N__19915\
        );

    \I__4366\ : Span12Mux_s4_v
    port map (
            O => \N__19921\,
            I => \N__19912\
        );

    \I__4365\ : LocalMux
    port map (
            O => \N__19918\,
            I => \N__19909\
        );

    \I__4364\ : LocalMux
    port map (
            O => \N__19915\,
            I => \ppm_encoder_1.rudderZ0Z_10\
        );

    \I__4363\ : Odrv12
    port map (
            O => \N__19912\,
            I => \ppm_encoder_1.rudderZ0Z_10\
        );

    \I__4362\ : Odrv4
    port map (
            O => \N__19909\,
            I => \ppm_encoder_1.rudderZ0Z_10\
        );

    \I__4361\ : InMux
    port map (
            O => \N__19902\,
            I => \N__19899\
        );

    \I__4360\ : LocalMux
    port map (
            O => \N__19899\,
            I => \N__19896\
        );

    \I__4359\ : Span4Mux_h
    port map (
            O => \N__19896\,
            I => \N__19893\
        );

    \I__4358\ : Odrv4
    port map (
            O => \N__19893\,
            I => \ppm_encoder_1.N_383\
        );

    \I__4357\ : CascadeMux
    port map (
            O => \N__19890\,
            I => \ppm_encoder_1.N_385_cascade_\
        );

    \I__4356\ : InMux
    port map (
            O => \N__19887\,
            I => \N__19884\
        );

    \I__4355\ : LocalMux
    port map (
            O => \N__19884\,
            I => \N__19881\
        );

    \I__4354\ : Span4Mux_v
    port map (
            O => \N__19881\,
            I => \N__19878\
        );

    \I__4353\ : Span4Mux_v
    port map (
            O => \N__19878\,
            I => \N__19874\
        );

    \I__4352\ : InMux
    port map (
            O => \N__19877\,
            I => \N__19871\
        );

    \I__4351\ : Odrv4
    port map (
            O => \N__19874\,
            I => \ppm_encoder_1.throttleZ0Z_4\
        );

    \I__4350\ : LocalMux
    port map (
            O => \N__19871\,
            I => \ppm_encoder_1.throttleZ0Z_4\
        );

    \I__4349\ : CascadeMux
    port map (
            O => \N__19866\,
            I => \N__19863\
        );

    \I__4348\ : InMux
    port map (
            O => \N__19863\,
            I => \N__19855\
        );

    \I__4347\ : InMux
    port map (
            O => \N__19862\,
            I => \N__19852\
        );

    \I__4346\ : InMux
    port map (
            O => \N__19861\,
            I => \N__19849\
        );

    \I__4345\ : InMux
    port map (
            O => \N__19860\,
            I => \N__19844\
        );

    \I__4344\ : InMux
    port map (
            O => \N__19859\,
            I => \N__19844\
        );

    \I__4343\ : InMux
    port map (
            O => \N__19858\,
            I => \N__19841\
        );

    \I__4342\ : LocalMux
    port map (
            O => \N__19855\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_3\
        );

    \I__4341\ : LocalMux
    port map (
            O => \N__19852\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_3\
        );

    \I__4340\ : LocalMux
    port map (
            O => \N__19849\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_3\
        );

    \I__4339\ : LocalMux
    port map (
            O => \N__19844\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_3\
        );

    \I__4338\ : LocalMux
    port map (
            O => \N__19841\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_3\
        );

    \I__4337\ : InMux
    port map (
            O => \N__19830\,
            I => \N__19827\
        );

    \I__4336\ : LocalMux
    port map (
            O => \N__19827\,
            I => \N__19823\
        );

    \I__4335\ : CascadeMux
    port map (
            O => \N__19826\,
            I => \N__19812\
        );

    \I__4334\ : Span4Mux_h
    port map (
            O => \N__19823\,
            I => \N__19809\
        );

    \I__4333\ : InMux
    port map (
            O => \N__19822\,
            I => \N__19806\
        );

    \I__4332\ : InMux
    port map (
            O => \N__19821\,
            I => \N__19801\
        );

    \I__4331\ : InMux
    port map (
            O => \N__19820\,
            I => \N__19801\
        );

    \I__4330\ : InMux
    port map (
            O => \N__19819\,
            I => \N__19798\
        );

    \I__4329\ : InMux
    port map (
            O => \N__19818\,
            I => \N__19795\
        );

    \I__4328\ : InMux
    port map (
            O => \N__19817\,
            I => \N__19790\
        );

    \I__4327\ : InMux
    port map (
            O => \N__19816\,
            I => \N__19790\
        );

    \I__4326\ : InMux
    port map (
            O => \N__19815\,
            I => \N__19785\
        );

    \I__4325\ : InMux
    port map (
            O => \N__19812\,
            I => \N__19785\
        );

    \I__4324\ : Odrv4
    port map (
            O => \N__19809\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2\
        );

    \I__4323\ : LocalMux
    port map (
            O => \N__19806\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2\
        );

    \I__4322\ : LocalMux
    port map (
            O => \N__19801\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2\
        );

    \I__4321\ : LocalMux
    port map (
            O => \N__19798\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2\
        );

    \I__4320\ : LocalMux
    port map (
            O => \N__19795\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2\
        );

    \I__4319\ : LocalMux
    port map (
            O => \N__19790\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2\
        );

    \I__4318\ : LocalMux
    port map (
            O => \N__19785\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2\
        );

    \I__4317\ : InMux
    port map (
            O => \N__19770\,
            I => \N__19762\
        );

    \I__4316\ : InMux
    port map (
            O => \N__19769\,
            I => \N__19759\
        );

    \I__4315\ : CascadeMux
    port map (
            O => \N__19768\,
            I => \N__19756\
        );

    \I__4314\ : CascadeMux
    port map (
            O => \N__19767\,
            I => \N__19753\
        );

    \I__4313\ : CascadeMux
    port map (
            O => \N__19766\,
            I => \N__19750\
        );

    \I__4312\ : CascadeMux
    port map (
            O => \N__19765\,
            I => \N__19747\
        );

    \I__4311\ : LocalMux
    port map (
            O => \N__19762\,
            I => \N__19742\
        );

    \I__4310\ : LocalMux
    port map (
            O => \N__19759\,
            I => \N__19739\
        );

    \I__4309\ : InMux
    port map (
            O => \N__19756\,
            I => \N__19730\
        );

    \I__4308\ : InMux
    port map (
            O => \N__19753\,
            I => \N__19730\
        );

    \I__4307\ : InMux
    port map (
            O => \N__19750\,
            I => \N__19730\
        );

    \I__4306\ : InMux
    port map (
            O => \N__19747\,
            I => \N__19730\
        );

    \I__4305\ : InMux
    port map (
            O => \N__19746\,
            I => \N__19727\
        );

    \I__4304\ : InMux
    port map (
            O => \N__19745\,
            I => \N__19724\
        );

    \I__4303\ : Span4Mux_h
    port map (
            O => \N__19742\,
            I => \N__19715\
        );

    \I__4302\ : Span4Mux_h
    port map (
            O => \N__19739\,
            I => \N__19715\
        );

    \I__4301\ : LocalMux
    port map (
            O => \N__19730\,
            I => \N__19715\
        );

    \I__4300\ : LocalMux
    port map (
            O => \N__19727\,
            I => \N__19715\
        );

    \I__4299\ : LocalMux
    port map (
            O => \N__19724\,
            I => \N__19710\
        );

    \I__4298\ : Span4Mux_v
    port map (
            O => \N__19715\,
            I => \N__19707\
        );

    \I__4297\ : CascadeMux
    port map (
            O => \N__19714\,
            I => \N__19702\
        );

    \I__4296\ : InMux
    port map (
            O => \N__19713\,
            I => \N__19698\
        );

    \I__4295\ : Span4Mux_v
    port map (
            O => \N__19710\,
            I => \N__19695\
        );

    \I__4294\ : Span4Mux_h
    port map (
            O => \N__19707\,
            I => \N__19692\
        );

    \I__4293\ : CascadeMux
    port map (
            O => \N__19706\,
            I => \N__19683\
        );

    \I__4292\ : InMux
    port map (
            O => \N__19705\,
            I => \N__19680\
        );

    \I__4291\ : InMux
    port map (
            O => \N__19702\,
            I => \N__19675\
        );

    \I__4290\ : InMux
    port map (
            O => \N__19701\,
            I => \N__19675\
        );

    \I__4289\ : LocalMux
    port map (
            O => \N__19698\,
            I => \N__19672\
        );

    \I__4288\ : Span4Mux_h
    port map (
            O => \N__19695\,
            I => \N__19669\
        );

    \I__4287\ : Span4Mux_h
    port map (
            O => \N__19692\,
            I => \N__19666\
        );

    \I__4286\ : InMux
    port map (
            O => \N__19691\,
            I => \N__19655\
        );

    \I__4285\ : InMux
    port map (
            O => \N__19690\,
            I => \N__19655\
        );

    \I__4284\ : InMux
    port map (
            O => \N__19689\,
            I => \N__19655\
        );

    \I__4283\ : InMux
    port map (
            O => \N__19688\,
            I => \N__19655\
        );

    \I__4282\ : InMux
    port map (
            O => \N__19687\,
            I => \N__19655\
        );

    \I__4281\ : InMux
    port map (
            O => \N__19686\,
            I => \N__19650\
        );

    \I__4280\ : InMux
    port map (
            O => \N__19683\,
            I => \N__19650\
        );

    \I__4279\ : LocalMux
    port map (
            O => \N__19680\,
            I => \N__19643\
        );

    \I__4278\ : LocalMux
    port map (
            O => \N__19675\,
            I => \N__19643\
        );

    \I__4277\ : Span4Mux_h
    port map (
            O => \N__19672\,
            I => \N__19643\
        );

    \I__4276\ : Odrv4
    port map (
            O => \N__19669\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_3_repZ0Z2\
        );

    \I__4275\ : Odrv4
    port map (
            O => \N__19666\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_3_repZ0Z2\
        );

    \I__4274\ : LocalMux
    port map (
            O => \N__19655\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_3_repZ0Z2\
        );

    \I__4273\ : LocalMux
    port map (
            O => \N__19650\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_3_repZ0Z2\
        );

    \I__4272\ : Odrv4
    port map (
            O => \N__19643\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_3_repZ0Z2\
        );

    \I__4271\ : CascadeMux
    port map (
            O => \N__19632\,
            I => \N__19627\
        );

    \I__4270\ : InMux
    port map (
            O => \N__19631\,
            I => \N__19615\
        );

    \I__4269\ : InMux
    port map (
            O => \N__19630\,
            I => \N__19615\
        );

    \I__4268\ : InMux
    port map (
            O => \N__19627\,
            I => \N__19610\
        );

    \I__4267\ : InMux
    port map (
            O => \N__19626\,
            I => \N__19610\
        );

    \I__4266\ : InMux
    port map (
            O => \N__19625\,
            I => \N__19607\
        );

    \I__4265\ : InMux
    port map (
            O => \N__19624\,
            I => \N__19604\
        );

    \I__4264\ : InMux
    port map (
            O => \N__19623\,
            I => \N__19598\
        );

    \I__4263\ : InMux
    port map (
            O => \N__19622\,
            I => \N__19598\
        );

    \I__4262\ : InMux
    port map (
            O => \N__19621\,
            I => \N__19594\
        );

    \I__4261\ : CascadeMux
    port map (
            O => \N__19620\,
            I => \N__19588\
        );

    \I__4260\ : LocalMux
    port map (
            O => \N__19615\,
            I => \N__19582\
        );

    \I__4259\ : LocalMux
    port map (
            O => \N__19610\,
            I => \N__19582\
        );

    \I__4258\ : LocalMux
    port map (
            O => \N__19607\,
            I => \N__19577\
        );

    \I__4257\ : LocalMux
    port map (
            O => \N__19604\,
            I => \N__19577\
        );

    \I__4256\ : InMux
    port map (
            O => \N__19603\,
            I => \N__19574\
        );

    \I__4255\ : LocalMux
    port map (
            O => \N__19598\,
            I => \N__19571\
        );

    \I__4254\ : InMux
    port map (
            O => \N__19597\,
            I => \N__19568\
        );

    \I__4253\ : LocalMux
    port map (
            O => \N__19594\,
            I => \N__19565\
        );

    \I__4252\ : InMux
    port map (
            O => \N__19593\,
            I => \N__19558\
        );

    \I__4251\ : InMux
    port map (
            O => \N__19592\,
            I => \N__19558\
        );

    \I__4250\ : InMux
    port map (
            O => \N__19591\,
            I => \N__19558\
        );

    \I__4249\ : InMux
    port map (
            O => \N__19588\,
            I => \N__19555\
        );

    \I__4248\ : InMux
    port map (
            O => \N__19587\,
            I => \N__19548\
        );

    \I__4247\ : Span4Mux_v
    port map (
            O => \N__19582\,
            I => \N__19541\
        );

    \I__4246\ : Span4Mux_v
    port map (
            O => \N__19577\,
            I => \N__19541\
        );

    \I__4245\ : LocalMux
    port map (
            O => \N__19574\,
            I => \N__19541\
        );

    \I__4244\ : Span4Mux_v
    port map (
            O => \N__19571\,
            I => \N__19533\
        );

    \I__4243\ : LocalMux
    port map (
            O => \N__19568\,
            I => \N__19533\
        );

    \I__4242\ : Span4Mux_v
    port map (
            O => \N__19565\,
            I => \N__19526\
        );

    \I__4241\ : LocalMux
    port map (
            O => \N__19558\,
            I => \N__19526\
        );

    \I__4240\ : LocalMux
    port map (
            O => \N__19555\,
            I => \N__19526\
        );

    \I__4239\ : InMux
    port map (
            O => \N__19554\,
            I => \N__19521\
        );

    \I__4238\ : InMux
    port map (
            O => \N__19553\,
            I => \N__19521\
        );

    \I__4237\ : InMux
    port map (
            O => \N__19552\,
            I => \N__19516\
        );

    \I__4236\ : InMux
    port map (
            O => \N__19551\,
            I => \N__19516\
        );

    \I__4235\ : LocalMux
    port map (
            O => \N__19548\,
            I => \N__19513\
        );

    \I__4234\ : Span4Mux_h
    port map (
            O => \N__19541\,
            I => \N__19510\
        );

    \I__4233\ : InMux
    port map (
            O => \N__19540\,
            I => \N__19507\
        );

    \I__4232\ : InMux
    port map (
            O => \N__19539\,
            I => \N__19502\
        );

    \I__4231\ : InMux
    port map (
            O => \N__19538\,
            I => \N__19502\
        );

    \I__4230\ : Span4Mux_h
    port map (
            O => \N__19533\,
            I => \N__19497\
        );

    \I__4229\ : Span4Mux_h
    port map (
            O => \N__19526\,
            I => \N__19497\
        );

    \I__4228\ : LocalMux
    port map (
            O => \N__19521\,
            I => \N__19492\
        );

    \I__4227\ : LocalMux
    port map (
            O => \N__19516\,
            I => \N__19492\
        );

    \I__4226\ : Odrv4
    port map (
            O => \N__19513\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z1\
        );

    \I__4225\ : Odrv4
    port map (
            O => \N__19510\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z1\
        );

    \I__4224\ : LocalMux
    port map (
            O => \N__19507\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z1\
        );

    \I__4223\ : LocalMux
    port map (
            O => \N__19502\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z1\
        );

    \I__4222\ : Odrv4
    port map (
            O => \N__19497\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z1\
        );

    \I__4221\ : Odrv12
    port map (
            O => \N__19492\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z1\
        );

    \I__4220\ : CascadeMux
    port map (
            O => \N__19479\,
            I => \N__19476\
        );

    \I__4219\ : InMux
    port map (
            O => \N__19476\,
            I => \N__19472\
        );

    \I__4218\ : CascadeMux
    port map (
            O => \N__19475\,
            I => \N__19468\
        );

    \I__4217\ : LocalMux
    port map (
            O => \N__19472\,
            I => \N__19464\
        );

    \I__4216\ : InMux
    port map (
            O => \N__19471\,
            I => \N__19461\
        );

    \I__4215\ : InMux
    port map (
            O => \N__19468\,
            I => \N__19458\
        );

    \I__4214\ : InMux
    port map (
            O => \N__19467\,
            I => \N__19455\
        );

    \I__4213\ : Span4Mux_v
    port map (
            O => \N__19464\,
            I => \N__19452\
        );

    \I__4212\ : LocalMux
    port map (
            O => \N__19461\,
            I => \N__19449\
        );

    \I__4211\ : LocalMux
    port map (
            O => \N__19458\,
            I => \N__19444\
        );

    \I__4210\ : LocalMux
    port map (
            O => \N__19455\,
            I => \N__19444\
        );

    \I__4209\ : Span4Mux_s2_v
    port map (
            O => \N__19452\,
            I => \N__19441\
        );

    \I__4208\ : Span4Mux_h
    port map (
            O => \N__19449\,
            I => \N__19436\
        );

    \I__4207\ : Span4Mux_v
    port map (
            O => \N__19444\,
            I => \N__19436\
        );

    \I__4206\ : Odrv4
    port map (
            O => \N__19441\,
            I => \ppm_encoder_1.init_pulsesZ0Z_7\
        );

    \I__4205\ : Odrv4
    port map (
            O => \N__19436\,
            I => \ppm_encoder_1.init_pulsesZ0Z_7\
        );

    \I__4204\ : InMux
    port map (
            O => \N__19431\,
            I => \N__19428\
        );

    \I__4203\ : LocalMux
    port map (
            O => \N__19428\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_7\
        );

    \I__4202\ : CascadeMux
    port map (
            O => \N__19425\,
            I => \N__19421\
        );

    \I__4201\ : InMux
    port map (
            O => \N__19424\,
            I => \N__19418\
        );

    \I__4200\ : InMux
    port map (
            O => \N__19421\,
            I => \N__19415\
        );

    \I__4199\ : LocalMux
    port map (
            O => \N__19418\,
            I => \ppm_encoder_1.PPM_STATE_fastZ0Z_0\
        );

    \I__4198\ : LocalMux
    port map (
            O => \N__19415\,
            I => \ppm_encoder_1.PPM_STATE_fastZ0Z_0\
        );

    \I__4197\ : InMux
    port map (
            O => \N__19410\,
            I => \N__19407\
        );

    \I__4196\ : LocalMux
    port map (
            O => \N__19407\,
            I => \N__19402\
        );

    \I__4195\ : InMux
    port map (
            O => \N__19406\,
            I => \N__19399\
        );

    \I__4194\ : CascadeMux
    port map (
            O => \N__19405\,
            I => \N__19396\
        );

    \I__4193\ : Span4Mux_v
    port map (
            O => \N__19402\,
            I => \N__19393\
        );

    \I__4192\ : LocalMux
    port map (
            O => \N__19399\,
            I => \N__19390\
        );

    \I__4191\ : InMux
    port map (
            O => \N__19396\,
            I => \N__19387\
        );

    \I__4190\ : Span4Mux_h
    port map (
            O => \N__19393\,
            I => \N__19384\
        );

    \I__4189\ : Span4Mux_h
    port map (
            O => \N__19390\,
            I => \N__19381\
        );

    \I__4188\ : LocalMux
    port map (
            O => \N__19387\,
            I => \ppm_encoder_1.aileronZ0Z_11\
        );

    \I__4187\ : Odrv4
    port map (
            O => \N__19384\,
            I => \ppm_encoder_1.aileronZ0Z_11\
        );

    \I__4186\ : Odrv4
    port map (
            O => \N__19381\,
            I => \ppm_encoder_1.aileronZ0Z_11\
        );

    \I__4185\ : InMux
    port map (
            O => \N__19374\,
            I => \N__19370\
        );

    \I__4184\ : CascadeMux
    port map (
            O => \N__19373\,
            I => \N__19367\
        );

    \I__4183\ : LocalMux
    port map (
            O => \N__19370\,
            I => \N__19364\
        );

    \I__4182\ : InMux
    port map (
            O => \N__19367\,
            I => \N__19361\
        );

    \I__4181\ : Span4Mux_v
    port map (
            O => \N__19364\,
            I => \N__19357\
        );

    \I__4180\ : LocalMux
    port map (
            O => \N__19361\,
            I => \N__19354\
        );

    \I__4179\ : InMux
    port map (
            O => \N__19360\,
            I => \N__19351\
        );

    \I__4178\ : Span4Mux_h
    port map (
            O => \N__19357\,
            I => \N__19348\
        );

    \I__4177\ : Span4Mux_h
    port map (
            O => \N__19354\,
            I => \N__19345\
        );

    \I__4176\ : LocalMux
    port map (
            O => \N__19351\,
            I => \ppm_encoder_1.throttleZ0Z_12\
        );

    \I__4175\ : Odrv4
    port map (
            O => \N__19348\,
            I => \ppm_encoder_1.throttleZ0Z_12\
        );

    \I__4174\ : Odrv4
    port map (
            O => \N__19345\,
            I => \ppm_encoder_1.throttleZ0Z_12\
        );

    \I__4173\ : CascadeMux
    port map (
            O => \N__19338\,
            I => \N__19333\
        );

    \I__4172\ : CascadeMux
    port map (
            O => \N__19337\,
            I => \N__19330\
        );

    \I__4171\ : InMux
    port map (
            O => \N__19336\,
            I => \N__19325\
        );

    \I__4170\ : InMux
    port map (
            O => \N__19333\,
            I => \N__19325\
        );

    \I__4169\ : InMux
    port map (
            O => \N__19330\,
            I => \N__19322\
        );

    \I__4168\ : LocalMux
    port map (
            O => \N__19325\,
            I => \N__19319\
        );

    \I__4167\ : LocalMux
    port map (
            O => \N__19322\,
            I => \N__19315\
        );

    \I__4166\ : Span4Mux_h
    port map (
            O => \N__19319\,
            I => \N__19312\
        );

    \I__4165\ : InMux
    port map (
            O => \N__19318\,
            I => \N__19309\
        );

    \I__4164\ : Span4Mux_h
    port map (
            O => \N__19315\,
            I => \N__19306\
        );

    \I__4163\ : Span4Mux_v
    port map (
            O => \N__19312\,
            I => \N__19303\
        );

    \I__4162\ : LocalMux
    port map (
            O => \N__19309\,
            I => \ppm_encoder_1.init_pulsesZ0Z_12\
        );

    \I__4161\ : Odrv4
    port map (
            O => \N__19306\,
            I => \ppm_encoder_1.init_pulsesZ0Z_12\
        );

    \I__4160\ : Odrv4
    port map (
            O => \N__19303\,
            I => \ppm_encoder_1.init_pulsesZ0Z_12\
        );

    \I__4159\ : CascadeMux
    port map (
            O => \N__19296\,
            I => \N__19292\
        );

    \I__4158\ : InMux
    port map (
            O => \N__19295\,
            I => \N__19289\
        );

    \I__4157\ : InMux
    port map (
            O => \N__19292\,
            I => \N__19286\
        );

    \I__4156\ : LocalMux
    port map (
            O => \N__19289\,
            I => \N__19283\
        );

    \I__4155\ : LocalMux
    port map (
            O => \N__19286\,
            I => \N__19280\
        );

    \I__4154\ : Span4Mux_h
    port map (
            O => \N__19283\,
            I => \N__19277\
        );

    \I__4153\ : Span4Mux_v
    port map (
            O => \N__19280\,
            I => \N__19274\
        );

    \I__4152\ : Span4Mux_h
    port map (
            O => \N__19277\,
            I => \N__19271\
        );

    \I__4151\ : Odrv4
    port map (
            O => \N__19274\,
            I => \ppm_encoder_1.N_258_i_i\
        );

    \I__4150\ : Odrv4
    port map (
            O => \N__19271\,
            I => \ppm_encoder_1.N_258_i_i\
        );

    \I__4149\ : CascadeMux
    port map (
            O => \N__19266\,
            I => \N__19263\
        );

    \I__4148\ : InMux
    port map (
            O => \N__19263\,
            I => \N__19259\
        );

    \I__4147\ : InMux
    port map (
            O => \N__19262\,
            I => \N__19256\
        );

    \I__4146\ : LocalMux
    port map (
            O => \N__19259\,
            I => \N__19253\
        );

    \I__4145\ : LocalMux
    port map (
            O => \N__19256\,
            I => \N__19250\
        );

    \I__4144\ : Span4Mux_h
    port map (
            O => \N__19253\,
            I => \N__19247\
        );

    \I__4143\ : Span4Mux_h
    port map (
            O => \N__19250\,
            I => \N__19244\
        );

    \I__4142\ : Odrv4
    port map (
            O => \N__19247\,
            I => \ppm_encoder_1.N_257_i_i\
        );

    \I__4141\ : Odrv4
    port map (
            O => \N__19244\,
            I => \ppm_encoder_1.N_257_i_i\
        );

    \I__4140\ : InMux
    port map (
            O => \N__19239\,
            I => \N__19236\
        );

    \I__4139\ : LocalMux
    port map (
            O => \N__19236\,
            I => \N__19232\
        );

    \I__4138\ : InMux
    port map (
            O => \N__19235\,
            I => \N__19227\
        );

    \I__4137\ : Span4Mux_h
    port map (
            O => \N__19232\,
            I => \N__19224\
        );

    \I__4136\ : InMux
    port map (
            O => \N__19231\,
            I => \N__19221\
        );

    \I__4135\ : InMux
    port map (
            O => \N__19230\,
            I => \N__19218\
        );

    \I__4134\ : LocalMux
    port map (
            O => \N__19227\,
            I => \ppm_encoder_1.rudderZ0Z_6\
        );

    \I__4133\ : Odrv4
    port map (
            O => \N__19224\,
            I => \ppm_encoder_1.rudderZ0Z_6\
        );

    \I__4132\ : LocalMux
    port map (
            O => \N__19221\,
            I => \ppm_encoder_1.rudderZ0Z_6\
        );

    \I__4131\ : LocalMux
    port map (
            O => \N__19218\,
            I => \ppm_encoder_1.rudderZ0Z_6\
        );

    \I__4130\ : InMux
    port map (
            O => \N__19209\,
            I => \N__19206\
        );

    \I__4129\ : LocalMux
    port map (
            O => \N__19206\,
            I => \ppm_encoder_1.pulses2count_9_0_0_6\
        );

    \I__4128\ : InMux
    port map (
            O => \N__19203\,
            I => \N__19200\
        );

    \I__4127\ : LocalMux
    port map (
            O => \N__19200\,
            I => \N__19197\
        );

    \I__4126\ : Span4Mux_h
    port map (
            O => \N__19197\,
            I => \N__19194\
        );

    \I__4125\ : Span4Mux_v
    port map (
            O => \N__19194\,
            I => \N__19191\
        );

    \I__4124\ : Odrv4
    port map (
            O => \N__19191\,
            I => \ppm_encoder_1.N_301\
        );

    \I__4123\ : CascadeMux
    port map (
            O => \N__19188\,
            I => \N__19184\
        );

    \I__4122\ : InMux
    port map (
            O => \N__19187\,
            I => \N__19181\
        );

    \I__4121\ : InMux
    port map (
            O => \N__19184\,
            I => \N__19177\
        );

    \I__4120\ : LocalMux
    port map (
            O => \N__19181\,
            I => \N__19174\
        );

    \I__4119\ : CascadeMux
    port map (
            O => \N__19180\,
            I => \N__19171\
        );

    \I__4118\ : LocalMux
    port map (
            O => \N__19177\,
            I => \N__19167\
        );

    \I__4117\ : Span4Mux_h
    port map (
            O => \N__19174\,
            I => \N__19164\
        );

    \I__4116\ : InMux
    port map (
            O => \N__19171\,
            I => \N__19159\
        );

    \I__4115\ : InMux
    port map (
            O => \N__19170\,
            I => \N__19159\
        );

    \I__4114\ : Span4Mux_h
    port map (
            O => \N__19167\,
            I => \N__19156\
        );

    \I__4113\ : Span4Mux_v
    port map (
            O => \N__19164\,
            I => \N__19153\
        );

    \I__4112\ : LocalMux
    port map (
            O => \N__19159\,
            I => \N__19150\
        );

    \I__4111\ : Odrv4
    port map (
            O => \N__19156\,
            I => \ppm_encoder_1.init_pulsesZ0Z_6\
        );

    \I__4110\ : Odrv4
    port map (
            O => \N__19153\,
            I => \ppm_encoder_1.init_pulsesZ0Z_6\
        );

    \I__4109\ : Odrv4
    port map (
            O => \N__19150\,
            I => \ppm_encoder_1.init_pulsesZ0Z_6\
        );

    \I__4108\ : InMux
    port map (
            O => \N__19143\,
            I => \N__19140\
        );

    \I__4107\ : LocalMux
    port map (
            O => \N__19140\,
            I => \ppm_encoder_1.pulses2countZ0Z_6\
        );

    \I__4106\ : InMux
    port map (
            O => \N__19137\,
            I => \N__19134\
        );

    \I__4105\ : LocalMux
    port map (
            O => \N__19134\,
            I => \N__19131\
        );

    \I__4104\ : Odrv12
    port map (
            O => \N__19131\,
            I => \ppm_encoder_1.N_302\
        );

    \I__4103\ : CascadeMux
    port map (
            O => \N__19128\,
            I => \N__19125\
        );

    \I__4102\ : InMux
    port map (
            O => \N__19125\,
            I => \N__19122\
        );

    \I__4101\ : LocalMux
    port map (
            O => \N__19122\,
            I => \ppm_encoder_1.pulses2countZ0Z_7\
        );

    \I__4100\ : InMux
    port map (
            O => \N__19119\,
            I => \N__19116\
        );

    \I__4099\ : LocalMux
    port map (
            O => \N__19116\,
            I => \ppm_encoder_1.pulses2count_9_0_2_12\
        );

    \I__4098\ : CascadeMux
    port map (
            O => \N__19113\,
            I => \N__19110\
        );

    \I__4097\ : InMux
    port map (
            O => \N__19110\,
            I => \N__19107\
        );

    \I__4096\ : LocalMux
    port map (
            O => \N__19107\,
            I => \N__19104\
        );

    \I__4095\ : Odrv4
    port map (
            O => \N__19104\,
            I => \ppm_encoder_1.N_393\
        );

    \I__4094\ : InMux
    port map (
            O => \N__19101\,
            I => \N__19098\
        );

    \I__4093\ : LocalMux
    port map (
            O => \N__19098\,
            I => \N__19095\
        );

    \I__4092\ : Odrv4
    port map (
            O => \N__19095\,
            I => \ppm_encoder_1.pulses2count_9_0_0_12\
        );

    \I__4091\ : CascadeMux
    port map (
            O => \N__19092\,
            I => \N__19089\
        );

    \I__4090\ : InMux
    port map (
            O => \N__19089\,
            I => \N__19085\
        );

    \I__4089\ : CascadeMux
    port map (
            O => \N__19088\,
            I => \N__19082\
        );

    \I__4088\ : LocalMux
    port map (
            O => \N__19085\,
            I => \N__19078\
        );

    \I__4087\ : InMux
    port map (
            O => \N__19082\,
            I => \N__19075\
        );

    \I__4086\ : InMux
    port map (
            O => \N__19081\,
            I => \N__19072\
        );

    \I__4085\ : Span4Mux_v
    port map (
            O => \N__19078\,
            I => \N__19069\
        );

    \I__4084\ : LocalMux
    port map (
            O => \N__19075\,
            I => \N__19066\
        );

    \I__4083\ : LocalMux
    port map (
            O => \N__19072\,
            I => \ppm_encoder_1.aileronZ0Z_12\
        );

    \I__4082\ : Odrv4
    port map (
            O => \N__19069\,
            I => \ppm_encoder_1.aileronZ0Z_12\
        );

    \I__4081\ : Odrv12
    port map (
            O => \N__19066\,
            I => \ppm_encoder_1.aileronZ0Z_12\
        );

    \I__4080\ : CascadeMux
    port map (
            O => \N__19059\,
            I => \N__19056\
        );

    \I__4079\ : InMux
    port map (
            O => \N__19056\,
            I => \N__19053\
        );

    \I__4078\ : LocalMux
    port map (
            O => \N__19053\,
            I => \N__19050\
        );

    \I__4077\ : Odrv4
    port map (
            O => \N__19050\,
            I => \ppm_encoder_1.N_396\
        );

    \I__4076\ : InMux
    port map (
            O => \N__19047\,
            I => \N__19044\
        );

    \I__4075\ : LocalMux
    port map (
            O => \N__19044\,
            I => \N__19040\
        );

    \I__4074\ : InMux
    port map (
            O => \N__19043\,
            I => \N__19037\
        );

    \I__4073\ : Span4Mux_h
    port map (
            O => \N__19040\,
            I => \N__19033\
        );

    \I__4072\ : LocalMux
    port map (
            O => \N__19037\,
            I => \N__19030\
        );

    \I__4071\ : InMux
    port map (
            O => \N__19036\,
            I => \N__19027\
        );

    \I__4070\ : Span4Mux_h
    port map (
            O => \N__19033\,
            I => \N__19024\
        );

    \I__4069\ : Span4Mux_h
    port map (
            O => \N__19030\,
            I => \N__19021\
        );

    \I__4068\ : LocalMux
    port map (
            O => \N__19027\,
            I => \ppm_encoder_1.elevatorZ0Z_12\
        );

    \I__4067\ : Odrv4
    port map (
            O => \N__19024\,
            I => \ppm_encoder_1.elevatorZ0Z_12\
        );

    \I__4066\ : Odrv4
    port map (
            O => \N__19021\,
            I => \ppm_encoder_1.elevatorZ0Z_12\
        );

    \I__4065\ : InMux
    port map (
            O => \N__19014\,
            I => \N__19011\
        );

    \I__4064\ : LocalMux
    port map (
            O => \N__19011\,
            I => \N__19007\
        );

    \I__4063\ : CascadeMux
    port map (
            O => \N__19010\,
            I => \N__19004\
        );

    \I__4062\ : Span4Mux_h
    port map (
            O => \N__19007\,
            I => \N__19001\
        );

    \I__4061\ : InMux
    port map (
            O => \N__19004\,
            I => \N__18997\
        );

    \I__4060\ : Span4Mux_v
    port map (
            O => \N__19001\,
            I => \N__18994\
        );

    \I__4059\ : InMux
    port map (
            O => \N__19000\,
            I => \N__18991\
        );

    \I__4058\ : LocalMux
    port map (
            O => \N__18997\,
            I => \ppm_encoder_1.throttleZ0Z_9\
        );

    \I__4057\ : Odrv4
    port map (
            O => \N__18994\,
            I => \ppm_encoder_1.throttleZ0Z_9\
        );

    \I__4056\ : LocalMux
    port map (
            O => \N__18991\,
            I => \ppm_encoder_1.throttleZ0Z_9\
        );

    \I__4055\ : InMux
    port map (
            O => \N__18984\,
            I => \N__18981\
        );

    \I__4054\ : LocalMux
    port map (
            O => \N__18981\,
            I => \N__18978\
        );

    \I__4053\ : Span4Mux_h
    port map (
            O => \N__18978\,
            I => \N__18975\
        );

    \I__4052\ : Odrv4
    port map (
            O => \N__18975\,
            I => \ppm_encoder_1.N_325\
        );

    \I__4051\ : CascadeMux
    port map (
            O => \N__18972\,
            I => \ppm_encoder_1.N_327_cascade_\
        );

    \I__4050\ : InMux
    port map (
            O => \N__18969\,
            I => \N__18966\
        );

    \I__4049\ : LocalMux
    port map (
            O => \N__18966\,
            I => \N__18962\
        );

    \I__4048\ : CascadeMux
    port map (
            O => \N__18965\,
            I => \N__18959\
        );

    \I__4047\ : Span4Mux_h
    port map (
            O => \N__18962\,
            I => \N__18956\
        );

    \I__4046\ : InMux
    port map (
            O => \N__18959\,
            I => \N__18952\
        );

    \I__4045\ : Span4Mux_h
    port map (
            O => \N__18956\,
            I => \N__18949\
        );

    \I__4044\ : InMux
    port map (
            O => \N__18955\,
            I => \N__18946\
        );

    \I__4043\ : LocalMux
    port map (
            O => \N__18952\,
            I => \ppm_encoder_1.rudderZ0Z_9\
        );

    \I__4042\ : Odrv4
    port map (
            O => \N__18949\,
            I => \ppm_encoder_1.rudderZ0Z_9\
        );

    \I__4041\ : LocalMux
    port map (
            O => \N__18946\,
            I => \ppm_encoder_1.rudderZ0Z_9\
        );

    \I__4040\ : InMux
    port map (
            O => \N__18939\,
            I => \N__18936\
        );

    \I__4039\ : LocalMux
    port map (
            O => \N__18936\,
            I => \N__18933\
        );

    \I__4038\ : Span4Mux_h
    port map (
            O => \N__18933\,
            I => \N__18929\
        );

    \I__4037\ : InMux
    port map (
            O => \N__18932\,
            I => \N__18926\
        );

    \I__4036\ : Odrv4
    port map (
            O => \N__18929\,
            I => \ppm_encoder_1.throttleZ0Z_5\
        );

    \I__4035\ : LocalMux
    port map (
            O => \N__18926\,
            I => \ppm_encoder_1.throttleZ0Z_5\
        );

    \I__4034\ : InMux
    port map (
            O => \N__18921\,
            I => \N__18917\
        );

    \I__4033\ : InMux
    port map (
            O => \N__18920\,
            I => \N__18914\
        );

    \I__4032\ : LocalMux
    port map (
            O => \N__18917\,
            I => \N__18911\
        );

    \I__4031\ : LocalMux
    port map (
            O => \N__18914\,
            I => \N__18908\
        );

    \I__4030\ : Odrv4
    port map (
            O => \N__18911\,
            I => \ppm_encoder_1.pulses2count_9_i_o2_0_5\
        );

    \I__4029\ : Odrv4
    port map (
            O => \N__18908\,
            I => \ppm_encoder_1.pulses2count_9_i_o2_0_5\
        );

    \I__4028\ : InMux
    port map (
            O => \N__18903\,
            I => \N__18894\
        );

    \I__4027\ : InMux
    port map (
            O => \N__18902\,
            I => \N__18890\
        );

    \I__4026\ : InMux
    port map (
            O => \N__18901\,
            I => \N__18887\
        );

    \I__4025\ : CascadeMux
    port map (
            O => \N__18900\,
            I => \N__18882\
        );

    \I__4024\ : InMux
    port map (
            O => \N__18899\,
            I => \N__18878\
        );

    \I__4023\ : InMux
    port map (
            O => \N__18898\,
            I => \N__18871\
        );

    \I__4022\ : InMux
    port map (
            O => \N__18897\,
            I => \N__18871\
        );

    \I__4021\ : LocalMux
    port map (
            O => \N__18894\,
            I => \N__18868\
        );

    \I__4020\ : InMux
    port map (
            O => \N__18893\,
            I => \N__18865\
        );

    \I__4019\ : LocalMux
    port map (
            O => \N__18890\,
            I => \N__18860\
        );

    \I__4018\ : LocalMux
    port map (
            O => \N__18887\,
            I => \N__18860\
        );

    \I__4017\ : InMux
    port map (
            O => \N__18886\,
            I => \N__18855\
        );

    \I__4016\ : InMux
    port map (
            O => \N__18885\,
            I => \N__18855\
        );

    \I__4015\ : InMux
    port map (
            O => \N__18882\,
            I => \N__18851\
        );

    \I__4014\ : CascadeMux
    port map (
            O => \N__18881\,
            I => \N__18848\
        );

    \I__4013\ : LocalMux
    port map (
            O => \N__18878\,
            I => \N__18845\
        );

    \I__4012\ : InMux
    port map (
            O => \N__18877\,
            I => \N__18842\
        );

    \I__4011\ : InMux
    port map (
            O => \N__18876\,
            I => \N__18839\
        );

    \I__4010\ : LocalMux
    port map (
            O => \N__18871\,
            I => \N__18836\
        );

    \I__4009\ : Span4Mux_h
    port map (
            O => \N__18868\,
            I => \N__18827\
        );

    \I__4008\ : LocalMux
    port map (
            O => \N__18865\,
            I => \N__18827\
        );

    \I__4007\ : Span4Mux_v
    port map (
            O => \N__18860\,
            I => \N__18827\
        );

    \I__4006\ : LocalMux
    port map (
            O => \N__18855\,
            I => \N__18827\
        );

    \I__4005\ : InMux
    port map (
            O => \N__18854\,
            I => \N__18823\
        );

    \I__4004\ : LocalMux
    port map (
            O => \N__18851\,
            I => \N__18820\
        );

    \I__4003\ : InMux
    port map (
            O => \N__18848\,
            I => \N__18817\
        );

    \I__4002\ : Span4Mux_h
    port map (
            O => \N__18845\,
            I => \N__18814\
        );

    \I__4001\ : LocalMux
    port map (
            O => \N__18842\,
            I => \N__18805\
        );

    \I__4000\ : LocalMux
    port map (
            O => \N__18839\,
            I => \N__18805\
        );

    \I__3999\ : Span4Mux_v
    port map (
            O => \N__18836\,
            I => \N__18805\
        );

    \I__3998\ : Span4Mux_h
    port map (
            O => \N__18827\,
            I => \N__18805\
        );

    \I__3997\ : InMux
    port map (
            O => \N__18826\,
            I => \N__18802\
        );

    \I__3996\ : LocalMux
    port map (
            O => \N__18823\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1\
        );

    \I__3995\ : Odrv12
    port map (
            O => \N__18820\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1\
        );

    \I__3994\ : LocalMux
    port map (
            O => \N__18817\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1\
        );

    \I__3993\ : Odrv4
    port map (
            O => \N__18814\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1\
        );

    \I__3992\ : Odrv4
    port map (
            O => \N__18805\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1\
        );

    \I__3991\ : LocalMux
    port map (
            O => \N__18802\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1\
        );

    \I__3990\ : CascadeMux
    port map (
            O => \N__18789\,
            I => \N__18784\
        );

    \I__3989\ : CascadeMux
    port map (
            O => \N__18788\,
            I => \N__18777\
        );

    \I__3988\ : InMux
    port map (
            O => \N__18787\,
            I => \N__18772\
        );

    \I__3987\ : InMux
    port map (
            O => \N__18784\,
            I => \N__18769\
        );

    \I__3986\ : InMux
    port map (
            O => \N__18783\,
            I => \N__18764\
        );

    \I__3985\ : InMux
    port map (
            O => \N__18782\,
            I => \N__18764\
        );

    \I__3984\ : CascadeMux
    port map (
            O => \N__18781\,
            I => \N__18760\
        );

    \I__3983\ : InMux
    port map (
            O => \N__18780\,
            I => \N__18756\
        );

    \I__3982\ : InMux
    port map (
            O => \N__18777\,
            I => \N__18751\
        );

    \I__3981\ : InMux
    port map (
            O => \N__18776\,
            I => \N__18751\
        );

    \I__3980\ : InMux
    port map (
            O => \N__18775\,
            I => \N__18748\
        );

    \I__3979\ : LocalMux
    port map (
            O => \N__18772\,
            I => \N__18745\
        );

    \I__3978\ : LocalMux
    port map (
            O => \N__18769\,
            I => \N__18742\
        );

    \I__3977\ : LocalMux
    port map (
            O => \N__18764\,
            I => \N__18736\
        );

    \I__3976\ : InMux
    port map (
            O => \N__18763\,
            I => \N__18732\
        );

    \I__3975\ : InMux
    port map (
            O => \N__18760\,
            I => \N__18727\
        );

    \I__3974\ : InMux
    port map (
            O => \N__18759\,
            I => \N__18727\
        );

    \I__3973\ : LocalMux
    port map (
            O => \N__18756\,
            I => \N__18724\
        );

    \I__3972\ : LocalMux
    port map (
            O => \N__18751\,
            I => \N__18721\
        );

    \I__3971\ : LocalMux
    port map (
            O => \N__18748\,
            I => \N__18716\
        );

    \I__3970\ : Span4Mux_v
    port map (
            O => \N__18745\,
            I => \N__18716\
        );

    \I__3969\ : Span4Mux_h
    port map (
            O => \N__18742\,
            I => \N__18713\
        );

    \I__3968\ : InMux
    port map (
            O => \N__18741\,
            I => \N__18710\
        );

    \I__3967\ : InMux
    port map (
            O => \N__18740\,
            I => \N__18707\
        );

    \I__3966\ : InMux
    port map (
            O => \N__18739\,
            I => \N__18704\
        );

    \I__3965\ : Span4Mux_h
    port map (
            O => \N__18736\,
            I => \N__18701\
        );

    \I__3964\ : InMux
    port map (
            O => \N__18735\,
            I => \N__18698\
        );

    \I__3963\ : LocalMux
    port map (
            O => \N__18732\,
            I => \N__18695\
        );

    \I__3962\ : LocalMux
    port map (
            O => \N__18727\,
            I => \N__18692\
        );

    \I__3961\ : Span4Mux_v
    port map (
            O => \N__18724\,
            I => \N__18687\
        );

    \I__3960\ : Span4Mux_h
    port map (
            O => \N__18721\,
            I => \N__18687\
        );

    \I__3959\ : Odrv4
    port map (
            O => \N__18716\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1\
        );

    \I__3958\ : Odrv4
    port map (
            O => \N__18713\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1\
        );

    \I__3957\ : LocalMux
    port map (
            O => \N__18710\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1\
        );

    \I__3956\ : LocalMux
    port map (
            O => \N__18707\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1\
        );

    \I__3955\ : LocalMux
    port map (
            O => \N__18704\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1\
        );

    \I__3954\ : Odrv4
    port map (
            O => \N__18701\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1\
        );

    \I__3953\ : LocalMux
    port map (
            O => \N__18698\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1\
        );

    \I__3952\ : Odrv12
    port map (
            O => \N__18695\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1\
        );

    \I__3951\ : Odrv4
    port map (
            O => \N__18692\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1\
        );

    \I__3950\ : Odrv4
    port map (
            O => \N__18687\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1\
        );

    \I__3949\ : InMux
    port map (
            O => \N__18666\,
            I => \N__18663\
        );

    \I__3948\ : LocalMux
    port map (
            O => \N__18663\,
            I => \N__18660\
        );

    \I__3947\ : Span4Mux_v
    port map (
            O => \N__18660\,
            I => \N__18657\
        );

    \I__3946\ : Odrv4
    port map (
            O => \N__18657\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_8\
        );

    \I__3945\ : CascadeMux
    port map (
            O => \N__18654\,
            I => \N__18650\
        );

    \I__3944\ : CascadeMux
    port map (
            O => \N__18653\,
            I => \N__18647\
        );

    \I__3943\ : InMux
    port map (
            O => \N__18650\,
            I => \N__18644\
        );

    \I__3942\ : InMux
    port map (
            O => \N__18647\,
            I => \N__18641\
        );

    \I__3941\ : LocalMux
    port map (
            O => \N__18644\,
            I => \N__18637\
        );

    \I__3940\ : LocalMux
    port map (
            O => \N__18641\,
            I => \N__18634\
        );

    \I__3939\ : InMux
    port map (
            O => \N__18640\,
            I => \N__18631\
        );

    \I__3938\ : Span4Mux_v
    port map (
            O => \N__18637\,
            I => \N__18628\
        );

    \I__3937\ : Span12Mux_h
    port map (
            O => \N__18634\,
            I => \N__18623\
        );

    \I__3936\ : LocalMux
    port map (
            O => \N__18631\,
            I => \N__18623\
        );

    \I__3935\ : Odrv4
    port map (
            O => \N__18628\,
            I => \ppm_encoder_1.N_204\
        );

    \I__3934\ : Odrv12
    port map (
            O => \N__18623\,
            I => \ppm_encoder_1.N_204\
        );

    \I__3933\ : CascadeMux
    port map (
            O => \N__18618\,
            I => \N__18615\
        );

    \I__3932\ : InMux
    port map (
            O => \N__18615\,
            I => \N__18612\
        );

    \I__3931\ : LocalMux
    port map (
            O => \N__18612\,
            I => \N__18608\
        );

    \I__3930\ : InMux
    port map (
            O => \N__18611\,
            I => \N__18605\
        );

    \I__3929\ : Span4Mux_v
    port map (
            O => \N__18608\,
            I => \N__18600\
        );

    \I__3928\ : LocalMux
    port map (
            O => \N__18605\,
            I => \N__18600\
        );

    \I__3927\ : Odrv4
    port map (
            O => \N__18600\,
            I => \ppm_encoder_1.N_255_i_i\
        );

    \I__3926\ : CascadeMux
    port map (
            O => \N__18597\,
            I => \ppm_encoder_1.N_204_cascade_\
        );

    \I__3925\ : InMux
    port map (
            O => \N__18594\,
            I => \N__18591\
        );

    \I__3924\ : LocalMux
    port map (
            O => \N__18591\,
            I => \N__18586\
        );

    \I__3923\ : InMux
    port map (
            O => \N__18590\,
            I => \N__18581\
        );

    \I__3922\ : InMux
    port map (
            O => \N__18589\,
            I => \N__18581\
        );

    \I__3921\ : Odrv4
    port map (
            O => \N__18586\,
            I => \ppm_encoder_1.elevatorZ0Z_8\
        );

    \I__3920\ : LocalMux
    port map (
            O => \N__18581\,
            I => \ppm_encoder_1.elevatorZ0Z_8\
        );

    \I__3919\ : InMux
    port map (
            O => \N__18576\,
            I => \N__18573\
        );

    \I__3918\ : LocalMux
    port map (
            O => \N__18573\,
            I => \N__18568\
        );

    \I__3917\ : InMux
    port map (
            O => \N__18572\,
            I => \N__18563\
        );

    \I__3916\ : InMux
    port map (
            O => \N__18571\,
            I => \N__18563\
        );

    \I__3915\ : Odrv4
    port map (
            O => \N__18568\,
            I => \ppm_encoder_1.aileronZ0Z_8\
        );

    \I__3914\ : LocalMux
    port map (
            O => \N__18563\,
            I => \ppm_encoder_1.aileronZ0Z_8\
        );

    \I__3913\ : CascadeMux
    port map (
            O => \N__18558\,
            I => \ppm_encoder_1.N_379_cascade_\
        );

    \I__3912\ : CascadeMux
    port map (
            O => \N__18555\,
            I => \N__18552\
        );

    \I__3911\ : InMux
    port map (
            O => \N__18552\,
            I => \N__18547\
        );

    \I__3910\ : InMux
    port map (
            O => \N__18551\,
            I => \N__18544\
        );

    \I__3909\ : InMux
    port map (
            O => \N__18550\,
            I => \N__18541\
        );

    \I__3908\ : LocalMux
    port map (
            O => \N__18547\,
            I => \ppm_encoder_1.rudderZ0Z_8\
        );

    \I__3907\ : LocalMux
    port map (
            O => \N__18544\,
            I => \ppm_encoder_1.rudderZ0Z_8\
        );

    \I__3906\ : LocalMux
    port map (
            O => \N__18541\,
            I => \ppm_encoder_1.rudderZ0Z_8\
        );

    \I__3905\ : InMux
    port map (
            O => \N__18534\,
            I => \N__18529\
        );

    \I__3904\ : InMux
    port map (
            O => \N__18533\,
            I => \N__18526\
        );

    \I__3903\ : InMux
    port map (
            O => \N__18532\,
            I => \N__18523\
        );

    \I__3902\ : LocalMux
    port map (
            O => \N__18529\,
            I => \ppm_encoder_1.throttleZ0Z_7\
        );

    \I__3901\ : LocalMux
    port map (
            O => \N__18526\,
            I => \ppm_encoder_1.throttleZ0Z_7\
        );

    \I__3900\ : LocalMux
    port map (
            O => \N__18523\,
            I => \ppm_encoder_1.throttleZ0Z_7\
        );

    \I__3899\ : InMux
    port map (
            O => \N__18516\,
            I => \N__18513\
        );

    \I__3898\ : LocalMux
    port map (
            O => \N__18513\,
            I => \N__18509\
        );

    \I__3897\ : InMux
    port map (
            O => \N__18512\,
            I => \N__18506\
        );

    \I__3896\ : Odrv4
    port map (
            O => \N__18509\,
            I => \ppm_encoder_1.pulses2count_9_i_o2_0_7\
        );

    \I__3895\ : LocalMux
    port map (
            O => \N__18506\,
            I => \ppm_encoder_1.pulses2count_9_i_o2_0_7\
        );

    \I__3894\ : InMux
    port map (
            O => \N__18501\,
            I => \N__18498\
        );

    \I__3893\ : LocalMux
    port map (
            O => \N__18498\,
            I => \N__18495\
        );

    \I__3892\ : Span4Mux_h
    port map (
            O => \N__18495\,
            I => \N__18490\
        );

    \I__3891\ : InMux
    port map (
            O => \N__18494\,
            I => \N__18487\
        );

    \I__3890\ : CascadeMux
    port map (
            O => \N__18493\,
            I => \N__18484\
        );

    \I__3889\ : Span4Mux_v
    port map (
            O => \N__18490\,
            I => \N__18479\
        );

    \I__3888\ : LocalMux
    port map (
            O => \N__18487\,
            I => \N__18479\
        );

    \I__3887\ : InMux
    port map (
            O => \N__18484\,
            I => \N__18476\
        );

    \I__3886\ : Span4Mux_h
    port map (
            O => \N__18479\,
            I => \N__18473\
        );

    \I__3885\ : LocalMux
    port map (
            O => \N__18476\,
            I => \ppm_encoder_1.rudderZ0Z_12\
        );

    \I__3884\ : Odrv4
    port map (
            O => \N__18473\,
            I => \ppm_encoder_1.rudderZ0Z_12\
        );

    \I__3883\ : InMux
    port map (
            O => \N__18468\,
            I => \N__18465\
        );

    \I__3882\ : LocalMux
    port map (
            O => \N__18465\,
            I => \N__18462\
        );

    \I__3881\ : Span4Mux_h
    port map (
            O => \N__18462\,
            I => \N__18459\
        );

    \I__3880\ : Span4Mux_v
    port map (
            O => \N__18459\,
            I => \N__18454\
        );

    \I__3879\ : InMux
    port map (
            O => \N__18458\,
            I => \N__18449\
        );

    \I__3878\ : InMux
    port map (
            O => \N__18457\,
            I => \N__18449\
        );

    \I__3877\ : Odrv4
    port map (
            O => \N__18454\,
            I => \ppm_encoder_1.elevatorZ0Z_11\
        );

    \I__3876\ : LocalMux
    port map (
            O => \N__18449\,
            I => \ppm_encoder_1.elevatorZ0Z_11\
        );

    \I__3875\ : CascadeMux
    port map (
            O => \N__18444\,
            I => \N__18441\
        );

    \I__3874\ : InMux
    port map (
            O => \N__18441\,
            I => \N__18438\
        );

    \I__3873\ : LocalMux
    port map (
            O => \N__18438\,
            I => \ppm_encoder_1.pulses2count_9_i_0_8\
        );

    \I__3872\ : InMux
    port map (
            O => \N__18435\,
            I => \N__18432\
        );

    \I__3871\ : LocalMux
    port map (
            O => \N__18432\,
            I => \N__18429\
        );

    \I__3870\ : Span4Mux_h
    port map (
            O => \N__18429\,
            I => \N__18424\
        );

    \I__3869\ : InMux
    port map (
            O => \N__18428\,
            I => \N__18419\
        );

    \I__3868\ : InMux
    port map (
            O => \N__18427\,
            I => \N__18419\
        );

    \I__3867\ : Odrv4
    port map (
            O => \N__18424\,
            I => \ppm_encoder_1.throttleZ0Z_8\
        );

    \I__3866\ : LocalMux
    port map (
            O => \N__18419\,
            I => \ppm_encoder_1.throttleZ0Z_8\
        );

    \I__3865\ : InMux
    port map (
            O => \N__18414\,
            I => \N__18410\
        );

    \I__3864\ : CascadeMux
    port map (
            O => \N__18413\,
            I => \N__18407\
        );

    \I__3863\ : LocalMux
    port map (
            O => \N__18410\,
            I => \N__18403\
        );

    \I__3862\ : InMux
    port map (
            O => \N__18407\,
            I => \N__18400\
        );

    \I__3861\ : InMux
    port map (
            O => \N__18406\,
            I => \N__18397\
        );

    \I__3860\ : Span4Mux_h
    port map (
            O => \N__18403\,
            I => \N__18392\
        );

    \I__3859\ : LocalMux
    port map (
            O => \N__18400\,
            I => \N__18392\
        );

    \I__3858\ : LocalMux
    port map (
            O => \N__18397\,
            I => \ppm_encoder_1.rudderZ0Z_11\
        );

    \I__3857\ : Odrv4
    port map (
            O => \N__18392\,
            I => \ppm_encoder_1.rudderZ0Z_11\
        );

    \I__3856\ : CascadeMux
    port map (
            O => \N__18387\,
            I => \N__18384\
        );

    \I__3855\ : InMux
    port map (
            O => \N__18384\,
            I => \N__18381\
        );

    \I__3854\ : LocalMux
    port map (
            O => \N__18381\,
            I => \ppm_encoder_1.N_391\
        );

    \I__3853\ : InMux
    port map (
            O => \N__18378\,
            I => \N__18375\
        );

    \I__3852\ : LocalMux
    port map (
            O => \N__18375\,
            I => \ppm_encoder_1.un1_init_pulses_11_15\
        );

    \I__3851\ : InMux
    port map (
            O => \N__18372\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_14\
        );

    \I__3850\ : InMux
    port map (
            O => \N__18369\,
            I => \N__18366\
        );

    \I__3849\ : LocalMux
    port map (
            O => \N__18366\,
            I => \N__18363\
        );

    \I__3848\ : Span4Mux_v
    port map (
            O => \N__18363\,
            I => \N__18360\
        );

    \I__3847\ : Odrv4
    port map (
            O => \N__18360\,
            I => \ppm_encoder_1.un1_init_pulses_11_16\
        );

    \I__3846\ : InMux
    port map (
            O => \N__18357\,
            I => \bfn_9_28_0_\
        );

    \I__3845\ : CascadeMux
    port map (
            O => \N__18354\,
            I => \N__18351\
        );

    \I__3844\ : InMux
    port map (
            O => \N__18351\,
            I => \N__18348\
        );

    \I__3843\ : LocalMux
    port map (
            O => \N__18348\,
            I => \N__18345\
        );

    \I__3842\ : Odrv4
    port map (
            O => \N__18345\,
            I => \ppm_encoder_1.un1_init_pulses_11_17\
        );

    \I__3841\ : InMux
    port map (
            O => \N__18342\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_16\
        );

    \I__3840\ : InMux
    port map (
            O => \N__18339\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_17\
        );

    \I__3839\ : InMux
    port map (
            O => \N__18336\,
            I => \N__18333\
        );

    \I__3838\ : LocalMux
    port map (
            O => \N__18333\,
            I => \N__18330\
        );

    \I__3837\ : Odrv4
    port map (
            O => \N__18330\,
            I => \ppm_encoder_1.un1_init_pulses_11_18\
        );

    \I__3836\ : InMux
    port map (
            O => \N__18327\,
            I => \N__18324\
        );

    \I__3835\ : LocalMux
    port map (
            O => \N__18324\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_16\
        );

    \I__3834\ : InMux
    port map (
            O => \N__18321\,
            I => \N__18318\
        );

    \I__3833\ : LocalMux
    port map (
            O => \N__18318\,
            I => \N__18314\
        );

    \I__3832\ : CascadeMux
    port map (
            O => \N__18317\,
            I => \N__18311\
        );

    \I__3831\ : Span4Mux_h
    port map (
            O => \N__18314\,
            I => \N__18308\
        );

    \I__3830\ : InMux
    port map (
            O => \N__18311\,
            I => \N__18305\
        );

    \I__3829\ : Odrv4
    port map (
            O => \N__18308\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_14\
        );

    \I__3828\ : LocalMux
    port map (
            O => \N__18305\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_14\
        );

    \I__3827\ : InMux
    port map (
            O => \N__18300\,
            I => \N__18297\
        );

    \I__3826\ : LocalMux
    port map (
            O => \N__18297\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_17\
        );

    \I__3825\ : CascadeMux
    port map (
            O => \N__18294\,
            I => \N__18291\
        );

    \I__3824\ : InMux
    port map (
            O => \N__18291\,
            I => \N__18286\
        );

    \I__3823\ : CascadeMux
    port map (
            O => \N__18290\,
            I => \N__18283\
        );

    \I__3822\ : InMux
    port map (
            O => \N__18289\,
            I => \N__18280\
        );

    \I__3821\ : LocalMux
    port map (
            O => \N__18286\,
            I => \N__18277\
        );

    \I__3820\ : InMux
    port map (
            O => \N__18283\,
            I => \N__18274\
        );

    \I__3819\ : LocalMux
    port map (
            O => \N__18280\,
            I => \N__18270\
        );

    \I__3818\ : Span4Mux_v
    port map (
            O => \N__18277\,
            I => \N__18267\
        );

    \I__3817\ : LocalMux
    port map (
            O => \N__18274\,
            I => \N__18264\
        );

    \I__3816\ : CascadeMux
    port map (
            O => \N__18273\,
            I => \N__18261\
        );

    \I__3815\ : Span4Mux_h
    port map (
            O => \N__18270\,
            I => \N__18258\
        );

    \I__3814\ : Span4Mux_h
    port map (
            O => \N__18267\,
            I => \N__18253\
        );

    \I__3813\ : Span4Mux_v
    port map (
            O => \N__18264\,
            I => \N__18253\
        );

    \I__3812\ : InMux
    port map (
            O => \N__18261\,
            I => \N__18250\
        );

    \I__3811\ : Odrv4
    port map (
            O => \N__18258\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_ns_2\
        );

    \I__3810\ : Odrv4
    port map (
            O => \N__18253\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_ns_2\
        );

    \I__3809\ : LocalMux
    port map (
            O => \N__18250\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_ns_2\
        );

    \I__3808\ : InMux
    port map (
            O => \N__18243\,
            I => \N__18240\
        );

    \I__3807\ : LocalMux
    port map (
            O => \N__18240\,
            I => \N__18237\
        );

    \I__3806\ : Odrv4
    port map (
            O => \N__18237\,
            I => \ppm_encoder_1.un1_init_pulses_11_7\
        );

    \I__3805\ : InMux
    port map (
            O => \N__18234\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_6\
        );

    \I__3804\ : CascadeMux
    port map (
            O => \N__18231\,
            I => \N__18228\
        );

    \I__3803\ : InMux
    port map (
            O => \N__18228\,
            I => \N__18225\
        );

    \I__3802\ : LocalMux
    port map (
            O => \N__18225\,
            I => \ppm_encoder_1.un1_init_pulses_11_8\
        );

    \I__3801\ : InMux
    port map (
            O => \N__18222\,
            I => \bfn_9_27_0_\
        );

    \I__3800\ : InMux
    port map (
            O => \N__18219\,
            I => \N__18216\
        );

    \I__3799\ : LocalMux
    port map (
            O => \N__18216\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_9\
        );

    \I__3798\ : InMux
    port map (
            O => \N__18213\,
            I => \N__18210\
        );

    \I__3797\ : LocalMux
    port map (
            O => \N__18210\,
            I => \ppm_encoder_1.un1_init_pulses_11_9\
        );

    \I__3796\ : InMux
    port map (
            O => \N__18207\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_8\
        );

    \I__3795\ : InMux
    port map (
            O => \N__18204\,
            I => \N__18201\
        );

    \I__3794\ : LocalMux
    port map (
            O => \N__18201\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_10\
        );

    \I__3793\ : InMux
    port map (
            O => \N__18198\,
            I => \N__18195\
        );

    \I__3792\ : LocalMux
    port map (
            O => \N__18195\,
            I => \ppm_encoder_1.un1_init_pulses_11_10\
        );

    \I__3791\ : InMux
    port map (
            O => \N__18192\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_9\
        );

    \I__3790\ : CascadeMux
    port map (
            O => \N__18189\,
            I => \N__18186\
        );

    \I__3789\ : InMux
    port map (
            O => \N__18186\,
            I => \N__18183\
        );

    \I__3788\ : LocalMux
    port map (
            O => \N__18183\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_11\
        );

    \I__3787\ : InMux
    port map (
            O => \N__18180\,
            I => \N__18177\
        );

    \I__3786\ : LocalMux
    port map (
            O => \N__18177\,
            I => \ppm_encoder_1.un1_init_pulses_11_11\
        );

    \I__3785\ : InMux
    port map (
            O => \N__18174\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_10\
        );

    \I__3784\ : InMux
    port map (
            O => \N__18171\,
            I => \N__18168\
        );

    \I__3783\ : LocalMux
    port map (
            O => \N__18168\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_12\
        );

    \I__3782\ : InMux
    port map (
            O => \N__18165\,
            I => \N__18162\
        );

    \I__3781\ : LocalMux
    port map (
            O => \N__18162\,
            I => \ppm_encoder_1.un1_init_pulses_11_12\
        );

    \I__3780\ : InMux
    port map (
            O => \N__18159\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_11\
        );

    \I__3779\ : InMux
    port map (
            O => \N__18156\,
            I => \N__18153\
        );

    \I__3778\ : LocalMux
    port map (
            O => \N__18153\,
            I => \N__18149\
        );

    \I__3777\ : InMux
    port map (
            O => \N__18152\,
            I => \N__18146\
        );

    \I__3776\ : Span4Mux_v
    port map (
            O => \N__18149\,
            I => \N__18140\
        );

    \I__3775\ : LocalMux
    port map (
            O => \N__18146\,
            I => \N__18140\
        );

    \I__3774\ : InMux
    port map (
            O => \N__18145\,
            I => \N__18137\
        );

    \I__3773\ : Span4Mux_h
    port map (
            O => \N__18140\,
            I => \N__18132\
        );

    \I__3772\ : LocalMux
    port map (
            O => \N__18137\,
            I => \N__18132\
        );

    \I__3771\ : Span4Mux_s3_v
    port map (
            O => \N__18132\,
            I => \N__18128\
        );

    \I__3770\ : InMux
    port map (
            O => \N__18131\,
            I => \N__18125\
        );

    \I__3769\ : Odrv4
    port map (
            O => \N__18128\,
            I => \ppm_encoder_1.N_259_i_i\
        );

    \I__3768\ : LocalMux
    port map (
            O => \N__18125\,
            I => \ppm_encoder_1.N_259_i_i\
        );

    \I__3767\ : CascadeMux
    port map (
            O => \N__18120\,
            I => \N__18117\
        );

    \I__3766\ : InMux
    port map (
            O => \N__18117\,
            I => \N__18114\
        );

    \I__3765\ : LocalMux
    port map (
            O => \N__18114\,
            I => \ppm_encoder_1.init_pulses_RNIKON03Z0Z_13\
        );

    \I__3764\ : InMux
    port map (
            O => \N__18111\,
            I => \N__18108\
        );

    \I__3763\ : LocalMux
    port map (
            O => \N__18108\,
            I => \ppm_encoder_1.un1_init_pulses_11_13\
        );

    \I__3762\ : InMux
    port map (
            O => \N__18105\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_12\
        );

    \I__3761\ : InMux
    port map (
            O => \N__18102\,
            I => \N__18099\
        );

    \I__3760\ : LocalMux
    port map (
            O => \N__18099\,
            I => \N__18096\
        );

    \I__3759\ : Odrv4
    port map (
            O => \N__18096\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_13_THRU_CO\
        );

    \I__3758\ : InMux
    port map (
            O => \N__18093\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_13\
        );

    \I__3757\ : CascadeMux
    port map (
            O => \N__18090\,
            I => \ppm_encoder_1.PPM_STATE_fast_RNI4RFRZ0Z_0_cascade_\
        );

    \I__3756\ : InMux
    port map (
            O => \N__18087\,
            I => \N__18084\
        );

    \I__3755\ : LocalMux
    port map (
            O => \N__18084\,
            I => \N__18081\
        );

    \I__3754\ : Span4Mux_v
    port map (
            O => \N__18081\,
            I => \N__18078\
        );

    \I__3753\ : Odrv4
    port map (
            O => \N__18078\,
            I => \ppm_encoder_1.init_pulses_RNI83R42Z0Z_0\
        );

    \I__3752\ : InMux
    port map (
            O => \N__18075\,
            I => \N__18072\
        );

    \I__3751\ : LocalMux
    port map (
            O => \N__18072\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_1\
        );

    \I__3750\ : InMux
    port map (
            O => \N__18069\,
            I => \N__18066\
        );

    \I__3749\ : LocalMux
    port map (
            O => \N__18066\,
            I => \ppm_encoder_1.un1_init_pulses_11_1\
        );

    \I__3748\ : InMux
    port map (
            O => \N__18063\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_0\
        );

    \I__3747\ : InMux
    port map (
            O => \N__18060\,
            I => \N__18057\
        );

    \I__3746\ : LocalMux
    port map (
            O => \N__18057\,
            I => \ppm_encoder_1.init_pulses_RNIGLA33Z0Z_2\
        );

    \I__3745\ : CascadeMux
    port map (
            O => \N__18054\,
            I => \N__18051\
        );

    \I__3744\ : InMux
    port map (
            O => \N__18051\,
            I => \N__18048\
        );

    \I__3743\ : LocalMux
    port map (
            O => \N__18048\,
            I => \N__18044\
        );

    \I__3742\ : CascadeMux
    port map (
            O => \N__18047\,
            I => \N__18041\
        );

    \I__3741\ : Span4Mux_h
    port map (
            O => \N__18044\,
            I => \N__18036\
        );

    \I__3740\ : InMux
    port map (
            O => \N__18041\,
            I => \N__18033\
        );

    \I__3739\ : InMux
    port map (
            O => \N__18040\,
            I => \N__18030\
        );

    \I__3738\ : InMux
    port map (
            O => \N__18039\,
            I => \N__18027\
        );

    \I__3737\ : Odrv4
    port map (
            O => \N__18036\,
            I => \ppm_encoder_1.N_249_i_i\
        );

    \I__3736\ : LocalMux
    port map (
            O => \N__18033\,
            I => \ppm_encoder_1.N_249_i_i\
        );

    \I__3735\ : LocalMux
    port map (
            O => \N__18030\,
            I => \ppm_encoder_1.N_249_i_i\
        );

    \I__3734\ : LocalMux
    port map (
            O => \N__18027\,
            I => \ppm_encoder_1.N_249_i_i\
        );

    \I__3733\ : InMux
    port map (
            O => \N__18018\,
            I => \N__18015\
        );

    \I__3732\ : LocalMux
    port map (
            O => \N__18015\,
            I => \N__18012\
        );

    \I__3731\ : Span4Mux_v
    port map (
            O => \N__18012\,
            I => \N__18009\
        );

    \I__3730\ : Odrv4
    port map (
            O => \N__18009\,
            I => \ppm_encoder_1.un1_init_pulses_11_2\
        );

    \I__3729\ : InMux
    port map (
            O => \N__18006\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_1\
        );

    \I__3728\ : InMux
    port map (
            O => \N__18003\,
            I => \N__18000\
        );

    \I__3727\ : LocalMux
    port map (
            O => \N__18000\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_3\
        );

    \I__3726\ : InMux
    port map (
            O => \N__17997\,
            I => \N__17994\
        );

    \I__3725\ : LocalMux
    port map (
            O => \N__17994\,
            I => \N__17991\
        );

    \I__3724\ : Odrv4
    port map (
            O => \N__17991\,
            I => \ppm_encoder_1.un1_init_pulses_11_3\
        );

    \I__3723\ : InMux
    port map (
            O => \N__17988\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_2\
        );

    \I__3722\ : InMux
    port map (
            O => \N__17985\,
            I => \N__17982\
        );

    \I__3721\ : LocalMux
    port map (
            O => \N__17982\,
            I => \N__17979\
        );

    \I__3720\ : Span4Mux_v
    port map (
            O => \N__17979\,
            I => \N__17976\
        );

    \I__3719\ : Odrv4
    port map (
            O => \N__17976\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_4\
        );

    \I__3718\ : InMux
    port map (
            O => \N__17973\,
            I => \N__17970\
        );

    \I__3717\ : LocalMux
    port map (
            O => \N__17970\,
            I => \N__17967\
        );

    \I__3716\ : Span4Mux_h
    port map (
            O => \N__17967\,
            I => \N__17964\
        );

    \I__3715\ : Odrv4
    port map (
            O => \N__17964\,
            I => \ppm_encoder_1.un1_init_pulses_11_4\
        );

    \I__3714\ : InMux
    port map (
            O => \N__17961\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_3\
        );

    \I__3713\ : InMux
    port map (
            O => \N__17958\,
            I => \N__17955\
        );

    \I__3712\ : LocalMux
    port map (
            O => \N__17955\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_5\
        );

    \I__3711\ : InMux
    port map (
            O => \N__17952\,
            I => \N__17949\
        );

    \I__3710\ : LocalMux
    port map (
            O => \N__17949\,
            I => \N__17946\
        );

    \I__3709\ : Odrv4
    port map (
            O => \N__17946\,
            I => \ppm_encoder_1.un1_init_pulses_11_5\
        );

    \I__3708\ : InMux
    port map (
            O => \N__17943\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_4\
        );

    \I__3707\ : InMux
    port map (
            O => \N__17940\,
            I => \N__17937\
        );

    \I__3706\ : LocalMux
    port map (
            O => \N__17937\,
            I => \ppm_encoder_1.init_pulses_RNI69BV2Z0Z_6\
        );

    \I__3705\ : CascadeMux
    port map (
            O => \N__17934\,
            I => \N__17930\
        );

    \I__3704\ : InMux
    port map (
            O => \N__17933\,
            I => \N__17926\
        );

    \I__3703\ : InMux
    port map (
            O => \N__17930\,
            I => \N__17923\
        );

    \I__3702\ : CascadeMux
    port map (
            O => \N__17929\,
            I => \N__17920\
        );

    \I__3701\ : LocalMux
    port map (
            O => \N__17926\,
            I => \N__17917\
        );

    \I__3700\ : LocalMux
    port map (
            O => \N__17923\,
            I => \N__17913\
        );

    \I__3699\ : InMux
    port map (
            O => \N__17920\,
            I => \N__17910\
        );

    \I__3698\ : Span4Mux_v
    port map (
            O => \N__17917\,
            I => \N__17907\
        );

    \I__3697\ : InMux
    port map (
            O => \N__17916\,
            I => \N__17904\
        );

    \I__3696\ : Odrv4
    port map (
            O => \N__17913\,
            I => \ppm_encoder_1.N_253_i_i\
        );

    \I__3695\ : LocalMux
    port map (
            O => \N__17910\,
            I => \ppm_encoder_1.N_253_i_i\
        );

    \I__3694\ : Odrv4
    port map (
            O => \N__17907\,
            I => \ppm_encoder_1.N_253_i_i\
        );

    \I__3693\ : LocalMux
    port map (
            O => \N__17904\,
            I => \ppm_encoder_1.N_253_i_i\
        );

    \I__3692\ : InMux
    port map (
            O => \N__17895\,
            I => \N__17892\
        );

    \I__3691\ : LocalMux
    port map (
            O => \N__17892\,
            I => \N__17889\
        );

    \I__3690\ : Odrv4
    port map (
            O => \N__17889\,
            I => \ppm_encoder_1.un1_init_pulses_11_6\
        );

    \I__3689\ : InMux
    port map (
            O => \N__17886\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_5\
        );

    \I__3688\ : InMux
    port map (
            O => \N__17883\,
            I => \N__17880\
        );

    \I__3687\ : LocalMux
    port map (
            O => \N__17880\,
            I => \N__17876\
        );

    \I__3686\ : InMux
    port map (
            O => \N__17879\,
            I => \N__17873\
        );

    \I__3685\ : Span4Mux_v
    port map (
            O => \N__17876\,
            I => \N__17866\
        );

    \I__3684\ : LocalMux
    port map (
            O => \N__17873\,
            I => \N__17866\
        );

    \I__3683\ : InMux
    port map (
            O => \N__17872\,
            I => \N__17861\
        );

    \I__3682\ : InMux
    port map (
            O => \N__17871\,
            I => \N__17858\
        );

    \I__3681\ : Span4Mux_h
    port map (
            O => \N__17866\,
            I => \N__17855\
        );

    \I__3680\ : InMux
    port map (
            O => \N__17865\,
            I => \N__17850\
        );

    \I__3679\ : InMux
    port map (
            O => \N__17864\,
            I => \N__17850\
        );

    \I__3678\ : LocalMux
    port map (
            O => \N__17861\,
            I => \N__17847\
        );

    \I__3677\ : LocalMux
    port map (
            O => \N__17858\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_1\
        );

    \I__3676\ : Odrv4
    port map (
            O => \N__17855\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_1\
        );

    \I__3675\ : LocalMux
    port map (
            O => \N__17850\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_1\
        );

    \I__3674\ : Odrv4
    port map (
            O => \N__17847\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_1\
        );

    \I__3673\ : CascadeMux
    port map (
            O => \N__17838\,
            I => \N__17835\
        );

    \I__3672\ : InMux
    port map (
            O => \N__17835\,
            I => \N__17831\
        );

    \I__3671\ : InMux
    port map (
            O => \N__17834\,
            I => \N__17828\
        );

    \I__3670\ : LocalMux
    port map (
            O => \N__17831\,
            I => \N__17825\
        );

    \I__3669\ : LocalMux
    port map (
            O => \N__17828\,
            I => \N__17822\
        );

    \I__3668\ : Odrv4
    port map (
            O => \N__17825\,
            I => \ppm_encoder_1.N_256_i_i\
        );

    \I__3667\ : Odrv12
    port map (
            O => \N__17822\,
            I => \ppm_encoder_1.N_256_i_i\
        );

    \I__3666\ : CascadeMux
    port map (
            O => \N__17817\,
            I => \N__17814\
        );

    \I__3665\ : InMux
    port map (
            O => \N__17814\,
            I => \N__17808\
        );

    \I__3664\ : CascadeMux
    port map (
            O => \N__17813\,
            I => \N__17799\
        );

    \I__3663\ : InMux
    port map (
            O => \N__17812\,
            I => \N__17796\
        );

    \I__3662\ : InMux
    port map (
            O => \N__17811\,
            I => \N__17793\
        );

    \I__3661\ : LocalMux
    port map (
            O => \N__17808\,
            I => \N__17790\
        );

    \I__3660\ : InMux
    port map (
            O => \N__17807\,
            I => \N__17787\
        );

    \I__3659\ : InMux
    port map (
            O => \N__17806\,
            I => \N__17782\
        );

    \I__3658\ : InMux
    port map (
            O => \N__17805\,
            I => \N__17782\
        );

    \I__3657\ : InMux
    port map (
            O => \N__17804\,
            I => \N__17777\
        );

    \I__3656\ : InMux
    port map (
            O => \N__17803\,
            I => \N__17777\
        );

    \I__3655\ : InMux
    port map (
            O => \N__17802\,
            I => \N__17772\
        );

    \I__3654\ : InMux
    port map (
            O => \N__17799\,
            I => \N__17772\
        );

    \I__3653\ : LocalMux
    port map (
            O => \N__17796\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_3_repZ0Z1\
        );

    \I__3652\ : LocalMux
    port map (
            O => \N__17793\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_3_repZ0Z1\
        );

    \I__3651\ : Odrv4
    port map (
            O => \N__17790\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_3_repZ0Z1\
        );

    \I__3650\ : LocalMux
    port map (
            O => \N__17787\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_3_repZ0Z1\
        );

    \I__3649\ : LocalMux
    port map (
            O => \N__17782\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_3_repZ0Z1\
        );

    \I__3648\ : LocalMux
    port map (
            O => \N__17777\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_3_repZ0Z1\
        );

    \I__3647\ : LocalMux
    port map (
            O => \N__17772\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_3_repZ0Z1\
        );

    \I__3646\ : InMux
    port map (
            O => \N__17757\,
            I => \N__17754\
        );

    \I__3645\ : LocalMux
    port map (
            O => \N__17754\,
            I => \N__17751\
        );

    \I__3644\ : Odrv4
    port map (
            O => \N__17751\,
            I => \ppm_encoder_1.un1_init_pulses_0_axb_16\
        );

    \I__3643\ : InMux
    port map (
            O => \N__17748\,
            I => \N__17745\
        );

    \I__3642\ : LocalMux
    port map (
            O => \N__17745\,
            I => \N__17741\
        );

    \I__3641\ : InMux
    port map (
            O => \N__17744\,
            I => \N__17738\
        );

    \I__3640\ : Span4Mux_h
    port map (
            O => \N__17741\,
            I => \N__17730\
        );

    \I__3639\ : LocalMux
    port map (
            O => \N__17738\,
            I => \N__17730\
        );

    \I__3638\ : InMux
    port map (
            O => \N__17737\,
            I => \N__17723\
        );

    \I__3637\ : InMux
    port map (
            O => \N__17736\,
            I => \N__17723\
        );

    \I__3636\ : InMux
    port map (
            O => \N__17735\,
            I => \N__17723\
        );

    \I__3635\ : Odrv4
    port map (
            O => \N__17730\,
            I => \ppm_encoder_1.N_305\
        );

    \I__3634\ : LocalMux
    port map (
            O => \N__17723\,
            I => \ppm_encoder_1.N_305\
        );

    \I__3633\ : InMux
    port map (
            O => \N__17718\,
            I => \N__17706\
        );

    \I__3632\ : InMux
    port map (
            O => \N__17717\,
            I => \N__17700\
        );

    \I__3631\ : InMux
    port map (
            O => \N__17716\,
            I => \N__17697\
        );

    \I__3630\ : InMux
    port map (
            O => \N__17715\,
            I => \N__17694\
        );

    \I__3629\ : InMux
    port map (
            O => \N__17714\,
            I => \N__17691\
        );

    \I__3628\ : InMux
    port map (
            O => \N__17713\,
            I => \N__17688\
        );

    \I__3627\ : InMux
    port map (
            O => \N__17712\,
            I => \N__17684\
        );

    \I__3626\ : InMux
    port map (
            O => \N__17711\,
            I => \N__17681\
        );

    \I__3625\ : InMux
    port map (
            O => \N__17710\,
            I => \N__17676\
        );

    \I__3624\ : InMux
    port map (
            O => \N__17709\,
            I => \N__17676\
        );

    \I__3623\ : LocalMux
    port map (
            O => \N__17706\,
            I => \N__17673\
        );

    \I__3622\ : InMux
    port map (
            O => \N__17705\,
            I => \N__17670\
        );

    \I__3621\ : CascadeMux
    port map (
            O => \N__17704\,
            I => \N__17663\
        );

    \I__3620\ : InMux
    port map (
            O => \N__17703\,
            I => \N__17660\
        );

    \I__3619\ : LocalMux
    port map (
            O => \N__17700\,
            I => \N__17657\
        );

    \I__3618\ : LocalMux
    port map (
            O => \N__17697\,
            I => \N__17650\
        );

    \I__3617\ : LocalMux
    port map (
            O => \N__17694\,
            I => \N__17650\
        );

    \I__3616\ : LocalMux
    port map (
            O => \N__17691\,
            I => \N__17650\
        );

    \I__3615\ : LocalMux
    port map (
            O => \N__17688\,
            I => \N__17647\
        );

    \I__3614\ : InMux
    port map (
            O => \N__17687\,
            I => \N__17644\
        );

    \I__3613\ : LocalMux
    port map (
            O => \N__17684\,
            I => \N__17637\
        );

    \I__3612\ : LocalMux
    port map (
            O => \N__17681\,
            I => \N__17637\
        );

    \I__3611\ : LocalMux
    port map (
            O => \N__17676\,
            I => \N__17637\
        );

    \I__3610\ : Span4Mux_v
    port map (
            O => \N__17673\,
            I => \N__17632\
        );

    \I__3609\ : LocalMux
    port map (
            O => \N__17670\,
            I => \N__17632\
        );

    \I__3608\ : InMux
    port map (
            O => \N__17669\,
            I => \N__17629\
        );

    \I__3607\ : InMux
    port map (
            O => \N__17668\,
            I => \N__17626\
        );

    \I__3606\ : InMux
    port map (
            O => \N__17667\,
            I => \N__17623\
        );

    \I__3605\ : InMux
    port map (
            O => \N__17666\,
            I => \N__17618\
        );

    \I__3604\ : InMux
    port map (
            O => \N__17663\,
            I => \N__17618\
        );

    \I__3603\ : LocalMux
    port map (
            O => \N__17660\,
            I => \N__17613\
        );

    \I__3602\ : Span4Mux_h
    port map (
            O => \N__17657\,
            I => \N__17613\
        );

    \I__3601\ : Span4Mux_v
    port map (
            O => \N__17650\,
            I => \N__17604\
        );

    \I__3600\ : Span4Mux_h
    port map (
            O => \N__17647\,
            I => \N__17604\
        );

    \I__3599\ : LocalMux
    port map (
            O => \N__17644\,
            I => \N__17604\
        );

    \I__3598\ : Span4Mux_v
    port map (
            O => \N__17637\,
            I => \N__17604\
        );

    \I__3597\ : Span4Mux_h
    port map (
            O => \N__17632\,
            I => \N__17601\
        );

    \I__3596\ : LocalMux
    port map (
            O => \N__17629\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIK17JZ0Z_3\
        );

    \I__3595\ : LocalMux
    port map (
            O => \N__17626\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIK17JZ0Z_3\
        );

    \I__3594\ : LocalMux
    port map (
            O => \N__17623\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIK17JZ0Z_3\
        );

    \I__3593\ : LocalMux
    port map (
            O => \N__17618\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIK17JZ0Z_3\
        );

    \I__3592\ : Odrv4
    port map (
            O => \N__17613\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIK17JZ0Z_3\
        );

    \I__3591\ : Odrv4
    port map (
            O => \N__17604\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIK17JZ0Z_3\
        );

    \I__3590\ : Odrv4
    port map (
            O => \N__17601\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIK17JZ0Z_3\
        );

    \I__3589\ : CascadeMux
    port map (
            O => \N__17586\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_2_cascade_\
        );

    \I__3588\ : InMux
    port map (
            O => \N__17583\,
            I => \N__17580\
        );

    \I__3587\ : LocalMux
    port map (
            O => \N__17580\,
            I => \N__17576\
        );

    \I__3586\ : InMux
    port map (
            O => \N__17579\,
            I => \N__17573\
        );

    \I__3585\ : Span4Mux_v
    port map (
            O => \N__17576\,
            I => \N__17568\
        );

    \I__3584\ : LocalMux
    port map (
            O => \N__17573\,
            I => \N__17568\
        );

    \I__3583\ : Odrv4
    port map (
            O => \N__17568\,
            I => \ppm_encoder_1.N_260_i_i\
        );

    \I__3582\ : CascadeMux
    port map (
            O => \N__17565\,
            I => \N__17556\
        );

    \I__3581\ : CascadeMux
    port map (
            O => \N__17564\,
            I => \N__17553\
        );

    \I__3580\ : InMux
    port map (
            O => \N__17563\,
            I => \N__17549\
        );

    \I__3579\ : CascadeMux
    port map (
            O => \N__17562\,
            I => \N__17545\
        );

    \I__3578\ : CascadeMux
    port map (
            O => \N__17561\,
            I => \N__17542\
        );

    \I__3577\ : CascadeMux
    port map (
            O => \N__17560\,
            I => \N__17536\
        );

    \I__3576\ : CascadeMux
    port map (
            O => \N__17559\,
            I => \N__17531\
        );

    \I__3575\ : InMux
    port map (
            O => \N__17556\,
            I => \N__17524\
        );

    \I__3574\ : InMux
    port map (
            O => \N__17553\,
            I => \N__17524\
        );

    \I__3573\ : CascadeMux
    port map (
            O => \N__17552\,
            I => \N__17521\
        );

    \I__3572\ : LocalMux
    port map (
            O => \N__17549\,
            I => \N__17517\
        );

    \I__3571\ : InMux
    port map (
            O => \N__17548\,
            I => \N__17510\
        );

    \I__3570\ : InMux
    port map (
            O => \N__17545\,
            I => \N__17510\
        );

    \I__3569\ : InMux
    port map (
            O => \N__17542\,
            I => \N__17510\
        );

    \I__3568\ : CascadeMux
    port map (
            O => \N__17541\,
            I => \N__17504\
        );

    \I__3567\ : CascadeMux
    port map (
            O => \N__17540\,
            I => \N__17501\
        );

    \I__3566\ : InMux
    port map (
            O => \N__17539\,
            I => \N__17496\
        );

    \I__3565\ : InMux
    port map (
            O => \N__17536\,
            I => \N__17496\
        );

    \I__3564\ : CascadeMux
    port map (
            O => \N__17535\,
            I => \N__17493\
        );

    \I__3563\ : InMux
    port map (
            O => \N__17534\,
            I => \N__17488\
        );

    \I__3562\ : InMux
    port map (
            O => \N__17531\,
            I => \N__17488\
        );

    \I__3561\ : CascadeMux
    port map (
            O => \N__17530\,
            I => \N__17480\
        );

    \I__3560\ : CascadeMux
    port map (
            O => \N__17529\,
            I => \N__17477\
        );

    \I__3559\ : LocalMux
    port map (
            O => \N__17524\,
            I => \N__17473\
        );

    \I__3558\ : InMux
    port map (
            O => \N__17521\,
            I => \N__17468\
        );

    \I__3557\ : InMux
    port map (
            O => \N__17520\,
            I => \N__17468\
        );

    \I__3556\ : Span4Mux_h
    port map (
            O => \N__17517\,
            I => \N__17463\
        );

    \I__3555\ : LocalMux
    port map (
            O => \N__17510\,
            I => \N__17463\
        );

    \I__3554\ : CascadeMux
    port map (
            O => \N__17509\,
            I => \N__17455\
        );

    \I__3553\ : InMux
    port map (
            O => \N__17508\,
            I => \N__17448\
        );

    \I__3552\ : InMux
    port map (
            O => \N__17507\,
            I => \N__17448\
        );

    \I__3551\ : InMux
    port map (
            O => \N__17504\,
            I => \N__17448\
        );

    \I__3550\ : InMux
    port map (
            O => \N__17501\,
            I => \N__17445\
        );

    \I__3549\ : LocalMux
    port map (
            O => \N__17496\,
            I => \N__17442\
        );

    \I__3548\ : InMux
    port map (
            O => \N__17493\,
            I => \N__17439\
        );

    \I__3547\ : LocalMux
    port map (
            O => \N__17488\,
            I => \N__17436\
        );

    \I__3546\ : InMux
    port map (
            O => \N__17487\,
            I => \N__17429\
        );

    \I__3545\ : InMux
    port map (
            O => \N__17486\,
            I => \N__17414\
        );

    \I__3544\ : InMux
    port map (
            O => \N__17485\,
            I => \N__17414\
        );

    \I__3543\ : InMux
    port map (
            O => \N__17484\,
            I => \N__17414\
        );

    \I__3542\ : InMux
    port map (
            O => \N__17483\,
            I => \N__17414\
        );

    \I__3541\ : InMux
    port map (
            O => \N__17480\,
            I => \N__17414\
        );

    \I__3540\ : InMux
    port map (
            O => \N__17477\,
            I => \N__17414\
        );

    \I__3539\ : InMux
    port map (
            O => \N__17476\,
            I => \N__17414\
        );

    \I__3538\ : Span4Mux_s3_v
    port map (
            O => \N__17473\,
            I => \N__17411\
        );

    \I__3537\ : LocalMux
    port map (
            O => \N__17468\,
            I => \N__17406\
        );

    \I__3536\ : Span4Mux_v
    port map (
            O => \N__17463\,
            I => \N__17406\
        );

    \I__3535\ : InMux
    port map (
            O => \N__17462\,
            I => \N__17403\
        );

    \I__3534\ : CascadeMux
    port map (
            O => \N__17461\,
            I => \N__17400\
        );

    \I__3533\ : CascadeMux
    port map (
            O => \N__17460\,
            I => \N__17397\
        );

    \I__3532\ : InMux
    port map (
            O => \N__17459\,
            I => \N__17390\
        );

    \I__3531\ : InMux
    port map (
            O => \N__17458\,
            I => \N__17390\
        );

    \I__3530\ : InMux
    port map (
            O => \N__17455\,
            I => \N__17390\
        );

    \I__3529\ : LocalMux
    port map (
            O => \N__17448\,
            I => \N__17383\
        );

    \I__3528\ : LocalMux
    port map (
            O => \N__17445\,
            I => \N__17383\
        );

    \I__3527\ : Span4Mux_s3_v
    port map (
            O => \N__17442\,
            I => \N__17383\
        );

    \I__3526\ : LocalMux
    port map (
            O => \N__17439\,
            I => \N__17380\
        );

    \I__3525\ : Span4Mux_h
    port map (
            O => \N__17436\,
            I => \N__17377\
        );

    \I__3524\ : InMux
    port map (
            O => \N__17435\,
            I => \N__17374\
        );

    \I__3523\ : InMux
    port map (
            O => \N__17434\,
            I => \N__17367\
        );

    \I__3522\ : InMux
    port map (
            O => \N__17433\,
            I => \N__17367\
        );

    \I__3521\ : InMux
    port map (
            O => \N__17432\,
            I => \N__17367\
        );

    \I__3520\ : LocalMux
    port map (
            O => \N__17429\,
            I => \N__17364\
        );

    \I__3519\ : LocalMux
    port map (
            O => \N__17414\,
            I => \N__17359\
        );

    \I__3518\ : Span4Mux_h
    port map (
            O => \N__17411\,
            I => \N__17359\
        );

    \I__3517\ : Span4Mux_h
    port map (
            O => \N__17406\,
            I => \N__17354\
        );

    \I__3516\ : LocalMux
    port map (
            O => \N__17403\,
            I => \N__17354\
        );

    \I__3515\ : InMux
    port map (
            O => \N__17400\,
            I => \N__17351\
        );

    \I__3514\ : InMux
    port map (
            O => \N__17397\,
            I => \N__17348\
        );

    \I__3513\ : LocalMux
    port map (
            O => \N__17390\,
            I => \N__17345\
        );

    \I__3512\ : Span4Mux_v
    port map (
            O => \N__17383\,
            I => \N__17342\
        );

    \I__3511\ : Span12Mux_h
    port map (
            O => \N__17380\,
            I => \N__17339\
        );

    \I__3510\ : Sp12to4
    port map (
            O => \N__17377\,
            I => \N__17336\
        );

    \I__3509\ : LocalMux
    port map (
            O => \N__17374\,
            I => \N__17325\
        );

    \I__3508\ : LocalMux
    port map (
            O => \N__17367\,
            I => \N__17325\
        );

    \I__3507\ : Span4Mux_h
    port map (
            O => \N__17364\,
            I => \N__17325\
        );

    \I__3506\ : Span4Mux_v
    port map (
            O => \N__17359\,
            I => \N__17325\
        );

    \I__3505\ : Span4Mux_h
    port map (
            O => \N__17354\,
            I => \N__17325\
        );

    \I__3504\ : LocalMux
    port map (
            O => \N__17351\,
            I => scaler_1_dv
        );

    \I__3503\ : LocalMux
    port map (
            O => \N__17348\,
            I => scaler_1_dv
        );

    \I__3502\ : Odrv12
    port map (
            O => \N__17345\,
            I => scaler_1_dv
        );

    \I__3501\ : Odrv4
    port map (
            O => \N__17342\,
            I => scaler_1_dv
        );

    \I__3500\ : Odrv12
    port map (
            O => \N__17339\,
            I => scaler_1_dv
        );

    \I__3499\ : Odrv12
    port map (
            O => \N__17336\,
            I => scaler_1_dv
        );

    \I__3498\ : Odrv4
    port map (
            O => \N__17325\,
            I => scaler_1_dv
        );

    \I__3497\ : InMux
    port map (
            O => \N__17310\,
            I => \N__17307\
        );

    \I__3496\ : LocalMux
    port map (
            O => \N__17307\,
            I => \N__17301\
        );

    \I__3495\ : InMux
    port map (
            O => \N__17306\,
            I => \N__17296\
        );

    \I__3494\ : InMux
    port map (
            O => \N__17305\,
            I => \N__17296\
        );

    \I__3493\ : InMux
    port map (
            O => \N__17304\,
            I => \N__17293\
        );

    \I__3492\ : Span4Mux_h
    port map (
            O => \N__17301\,
            I => \N__17288\
        );

    \I__3491\ : LocalMux
    port map (
            O => \N__17296\,
            I => \N__17288\
        );

    \I__3490\ : LocalMux
    port map (
            O => \N__17293\,
            I => \ppm_encoder_1.init_pulsesZ0Z_1\
        );

    \I__3489\ : Odrv4
    port map (
            O => \N__17288\,
            I => \ppm_encoder_1.init_pulsesZ0Z_1\
        );

    \I__3488\ : CascadeMux
    port map (
            O => \N__17283\,
            I => \N__17280\
        );

    \I__3487\ : InMux
    port map (
            O => \N__17280\,
            I => \N__17277\
        );

    \I__3486\ : LocalMux
    port map (
            O => \N__17277\,
            I => \N__17273\
        );

    \I__3485\ : InMux
    port map (
            O => \N__17276\,
            I => \N__17270\
        );

    \I__3484\ : Odrv4
    port map (
            O => \N__17273\,
            I => \ppm_encoder_1.N_248_i_i\
        );

    \I__3483\ : LocalMux
    port map (
            O => \N__17270\,
            I => \ppm_encoder_1.N_248_i_i\
        );

    \I__3482\ : CascadeMux
    port map (
            O => \N__17265\,
            I => \N__17262\
        );

    \I__3481\ : InMux
    port map (
            O => \N__17262\,
            I => \N__17259\
        );

    \I__3480\ : LocalMux
    port map (
            O => \N__17259\,
            I => \N__17255\
        );

    \I__3479\ : InMux
    port map (
            O => \N__17258\,
            I => \N__17252\
        );

    \I__3478\ : Odrv4
    port map (
            O => \N__17255\,
            I => \ppm_encoder_1.N_250_i_i\
        );

    \I__3477\ : LocalMux
    port map (
            O => \N__17252\,
            I => \ppm_encoder_1.N_250_i_i\
        );

    \I__3476\ : CascadeMux
    port map (
            O => \N__17247\,
            I => \N__17244\
        );

    \I__3475\ : InMux
    port map (
            O => \N__17244\,
            I => \N__17241\
        );

    \I__3474\ : LocalMux
    port map (
            O => \N__17241\,
            I => \N__17238\
        );

    \I__3473\ : Span4Mux_v
    port map (
            O => \N__17238\,
            I => \N__17235\
        );

    \I__3472\ : Span4Mux_h
    port map (
            O => \N__17235\,
            I => \N__17231\
        );

    \I__3471\ : InMux
    port map (
            O => \N__17234\,
            I => \N__17228\
        );

    \I__3470\ : Odrv4
    port map (
            O => \N__17231\,
            I => \ppm_encoder_1.N_254_i_i\
        );

    \I__3469\ : LocalMux
    port map (
            O => \N__17228\,
            I => \ppm_encoder_1.N_254_i_i\
        );

    \I__3468\ : CascadeMux
    port map (
            O => \N__17223\,
            I => \ppm_encoder_1.PPM_STATE_fast_RNICIABZ0Z_0_cascade_\
        );

    \I__3467\ : CascadeMux
    port map (
            O => \N__17220\,
            I => \N__17217\
        );

    \I__3466\ : InMux
    port map (
            O => \N__17217\,
            I => \N__17213\
        );

    \I__3465\ : InMux
    port map (
            O => \N__17216\,
            I => \N__17210\
        );

    \I__3464\ : LocalMux
    port map (
            O => \N__17213\,
            I => \N__17205\
        );

    \I__3463\ : LocalMux
    port map (
            O => \N__17210\,
            I => \N__17205\
        );

    \I__3462\ : Odrv12
    port map (
            O => \N__17205\,
            I => \ppm_encoder_1.N_246_i_i\
        );

    \I__3461\ : CascadeMux
    port map (
            O => \N__17202\,
            I => \ppm_encoder_1.un2_throttle_0_0_7_cascade_\
        );

    \I__3460\ : InMux
    port map (
            O => \N__17199\,
            I => \N__17196\
        );

    \I__3459\ : LocalMux
    port map (
            O => \N__17196\,
            I => \ppm_encoder_1.un1_init_pulses_0_axb_7\
        );

    \I__3458\ : InMux
    port map (
            O => \N__17193\,
            I => \N__17189\
        );

    \I__3457\ : InMux
    port map (
            O => \N__17192\,
            I => \N__17185\
        );

    \I__3456\ : LocalMux
    port map (
            O => \N__17189\,
            I => \N__17178\
        );

    \I__3455\ : InMux
    port map (
            O => \N__17188\,
            I => \N__17175\
        );

    \I__3454\ : LocalMux
    port map (
            O => \N__17185\,
            I => \N__17172\
        );

    \I__3453\ : InMux
    port map (
            O => \N__17184\,
            I => \N__17169\
        );

    \I__3452\ : InMux
    port map (
            O => \N__17183\,
            I => \N__17162\
        );

    \I__3451\ : InMux
    port map (
            O => \N__17182\,
            I => \N__17162\
        );

    \I__3450\ : InMux
    port map (
            O => \N__17181\,
            I => \N__17162\
        );

    \I__3449\ : Odrv4
    port map (
            O => \N__17178\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0\
        );

    \I__3448\ : LocalMux
    port map (
            O => \N__17175\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0\
        );

    \I__3447\ : Odrv4
    port map (
            O => \N__17172\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0\
        );

    \I__3446\ : LocalMux
    port map (
            O => \N__17169\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0\
        );

    \I__3445\ : LocalMux
    port map (
            O => \N__17162\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0\
        );

    \I__3444\ : CascadeMux
    port map (
            O => \N__17151\,
            I => \N__17148\
        );

    \I__3443\ : InMux
    port map (
            O => \N__17148\,
            I => \N__17144\
        );

    \I__3442\ : InMux
    port map (
            O => \N__17147\,
            I => \N__17141\
        );

    \I__3441\ : LocalMux
    port map (
            O => \N__17144\,
            I => \N__17138\
        );

    \I__3440\ : LocalMux
    port map (
            O => \N__17141\,
            I => \ppm_encoder_1.elevatorZ0Z_7\
        );

    \I__3439\ : Odrv12
    port map (
            O => \N__17138\,
            I => \ppm_encoder_1.elevatorZ0Z_7\
        );

    \I__3438\ : InMux
    port map (
            O => \N__17133\,
            I => \N__17130\
        );

    \I__3437\ : LocalMux
    port map (
            O => \N__17130\,
            I => \ppm_encoder_1.un2_throttle_iv_0_rn_0_7\
        );

    \I__3436\ : InMux
    port map (
            O => \N__17127\,
            I => \N__17124\
        );

    \I__3435\ : LocalMux
    port map (
            O => \N__17124\,
            I => \N__17121\
        );

    \I__3434\ : Span4Mux_v
    port map (
            O => \N__17121\,
            I => \N__17118\
        );

    \I__3433\ : Span4Mux_h
    port map (
            O => \N__17118\,
            I => \N__17115\
        );

    \I__3432\ : Odrv4
    port map (
            O => \N__17115\,
            I => \ppm_encoder_1.un1_aileron_cry_6_THRU_CO\
        );

    \I__3431\ : InMux
    port map (
            O => \N__17112\,
            I => \N__17109\
        );

    \I__3430\ : LocalMux
    port map (
            O => \N__17109\,
            I => \N__17106\
        );

    \I__3429\ : Span4Mux_h
    port map (
            O => \N__17106\,
            I => \N__17102\
        );

    \I__3428\ : InMux
    port map (
            O => \N__17105\,
            I => \N__17099\
        );

    \I__3427\ : Span4Mux_h
    port map (
            O => \N__17102\,
            I => \N__17096\
        );

    \I__3426\ : LocalMux
    port map (
            O => \N__17099\,
            I => \N__17093\
        );

    \I__3425\ : Odrv4
    port map (
            O => \N__17096\,
            I => scaler_2_data_7
        );

    \I__3424\ : Odrv4
    port map (
            O => \N__17093\,
            I => scaler_2_data_7
        );

    \I__3423\ : InMux
    port map (
            O => \N__17088\,
            I => \N__17082\
        );

    \I__3422\ : InMux
    port map (
            O => \N__17087\,
            I => \N__17082\
        );

    \I__3421\ : LocalMux
    port map (
            O => \N__17082\,
            I => \ppm_encoder_1.aileronZ0Z_7\
        );

    \I__3420\ : CascadeMux
    port map (
            O => \N__17079\,
            I => \ppm_encoder_1.un1_init_pulses_0_axb_1_cascade_\
        );

    \I__3419\ : InMux
    port map (
            O => \N__17076\,
            I => \N__17073\
        );

    \I__3418\ : LocalMux
    port map (
            O => \N__17073\,
            I => \N__17070\
        );

    \I__3417\ : Odrv4
    port map (
            O => \N__17070\,
            I => \ppm_encoder_1.init_pulses_RNIOC8K3Z0Z_1\
        );

    \I__3416\ : InMux
    port map (
            O => \N__17067\,
            I => \N__17064\
        );

    \I__3415\ : LocalMux
    port map (
            O => \N__17064\,
            I => \ppm_encoder_1.N_426\
        );

    \I__3414\ : InMux
    port map (
            O => \N__17061\,
            I => \N__17055\
        );

    \I__3413\ : InMux
    port map (
            O => \N__17060\,
            I => \N__17052\
        );

    \I__3412\ : InMux
    port map (
            O => \N__17059\,
            I => \N__17046\
        );

    \I__3411\ : InMux
    port map (
            O => \N__17058\,
            I => \N__17041\
        );

    \I__3410\ : LocalMux
    port map (
            O => \N__17055\,
            I => \N__17038\
        );

    \I__3409\ : LocalMux
    port map (
            O => \N__17052\,
            I => \N__17033\
        );

    \I__3408\ : InMux
    port map (
            O => \N__17051\,
            I => \N__17030\
        );

    \I__3407\ : InMux
    port map (
            O => \N__17050\,
            I => \N__17024\
        );

    \I__3406\ : InMux
    port map (
            O => \N__17049\,
            I => \N__17021\
        );

    \I__3405\ : LocalMux
    port map (
            O => \N__17046\,
            I => \N__17018\
        );

    \I__3404\ : InMux
    port map (
            O => \N__17045\,
            I => \N__17015\
        );

    \I__3403\ : InMux
    port map (
            O => \N__17044\,
            I => \N__17012\
        );

    \I__3402\ : LocalMux
    port map (
            O => \N__17041\,
            I => \N__17007\
        );

    \I__3401\ : Span4Mux_v
    port map (
            O => \N__17038\,
            I => \N__17007\
        );

    \I__3400\ : InMux
    port map (
            O => \N__17037\,
            I => \N__17002\
        );

    \I__3399\ : InMux
    port map (
            O => \N__17036\,
            I => \N__17002\
        );

    \I__3398\ : Span4Mux_v
    port map (
            O => \N__17033\,
            I => \N__16997\
        );

    \I__3397\ : LocalMux
    port map (
            O => \N__17030\,
            I => \N__16997\
        );

    \I__3396\ : InMux
    port map (
            O => \N__17029\,
            I => \N__16994\
        );

    \I__3395\ : InMux
    port map (
            O => \N__17028\,
            I => \N__16989\
        );

    \I__3394\ : InMux
    port map (
            O => \N__17027\,
            I => \N__16989\
        );

    \I__3393\ : LocalMux
    port map (
            O => \N__17024\,
            I => \N__16984\
        );

    \I__3392\ : LocalMux
    port map (
            O => \N__17021\,
            I => \N__16984\
        );

    \I__3391\ : Span4Mux_h
    port map (
            O => \N__17018\,
            I => \N__16981\
        );

    \I__3390\ : LocalMux
    port map (
            O => \N__17015\,
            I => \ppm_encoder_1.N_246\
        );

    \I__3389\ : LocalMux
    port map (
            O => \N__17012\,
            I => \ppm_encoder_1.N_246\
        );

    \I__3388\ : Odrv4
    port map (
            O => \N__17007\,
            I => \ppm_encoder_1.N_246\
        );

    \I__3387\ : LocalMux
    port map (
            O => \N__17002\,
            I => \ppm_encoder_1.N_246\
        );

    \I__3386\ : Odrv4
    port map (
            O => \N__16997\,
            I => \ppm_encoder_1.N_246\
        );

    \I__3385\ : LocalMux
    port map (
            O => \N__16994\,
            I => \ppm_encoder_1.N_246\
        );

    \I__3384\ : LocalMux
    port map (
            O => \N__16989\,
            I => \ppm_encoder_1.N_246\
        );

    \I__3383\ : Odrv4
    port map (
            O => \N__16984\,
            I => \ppm_encoder_1.N_246\
        );

    \I__3382\ : Odrv4
    port map (
            O => \N__16981\,
            I => \ppm_encoder_1.N_246\
        );

    \I__3381\ : CascadeMux
    port map (
            O => \N__16962\,
            I => \ppm_encoder_1.N_426_cascade_\
        );

    \I__3380\ : CascadeMux
    port map (
            O => \N__16959\,
            I => \ppm_encoder_1.un1_init_pulses_0_axb_3_cascade_\
        );

    \I__3379\ : InMux
    port map (
            O => \N__16956\,
            I => \N__16953\
        );

    \I__3378\ : LocalMux
    port map (
            O => \N__16953\,
            I => \N__16950\
        );

    \I__3377\ : Odrv4
    port map (
            O => \N__16950\,
            I => \ppm_encoder_1.init_pulses_RNISG8K3Z0Z_3\
        );

    \I__3376\ : InMux
    port map (
            O => \N__16947\,
            I => \N__16944\
        );

    \I__3375\ : LocalMux
    port map (
            O => \N__16944\,
            I => \N__16941\
        );

    \I__3374\ : Span4Mux_v
    port map (
            O => \N__16941\,
            I => \N__16938\
        );

    \I__3373\ : Odrv4
    port map (
            O => \N__16938\,
            I => \ppm_encoder_1.un1_init_pulses_10_6\
        );

    \I__3372\ : InMux
    port map (
            O => \N__16935\,
            I => \N__16932\
        );

    \I__3371\ : LocalMux
    port map (
            O => \N__16932\,
            I => \N__16929\
        );

    \I__3370\ : Span4Mux_v
    port map (
            O => \N__16929\,
            I => \N__16926\
        );

    \I__3369\ : Odrv4
    port map (
            O => \N__16926\,
            I => \ppm_encoder_1.un1_init_pulses_10_7\
        );

    \I__3368\ : CascadeMux
    port map (
            O => \N__16923\,
            I => \N__16915\
        );

    \I__3367\ : CascadeMux
    port map (
            O => \N__16922\,
            I => \N__16911\
        );

    \I__3366\ : CascadeMux
    port map (
            O => \N__16921\,
            I => \N__16907\
        );

    \I__3365\ : CascadeMux
    port map (
            O => \N__16920\,
            I => \N__16904\
        );

    \I__3364\ : CascadeMux
    port map (
            O => \N__16919\,
            I => \N__16901\
        );

    \I__3363\ : InMux
    port map (
            O => \N__16918\,
            I => \N__16896\
        );

    \I__3362\ : InMux
    port map (
            O => \N__16915\,
            I => \N__16896\
        );

    \I__3361\ : InMux
    port map (
            O => \N__16914\,
            I => \N__16889\
        );

    \I__3360\ : InMux
    port map (
            O => \N__16911\,
            I => \N__16889\
        );

    \I__3359\ : InMux
    port map (
            O => \N__16910\,
            I => \N__16889\
        );

    \I__3358\ : InMux
    port map (
            O => \N__16907\,
            I => \N__16882\
        );

    \I__3357\ : InMux
    port map (
            O => \N__16904\,
            I => \N__16882\
        );

    \I__3356\ : InMux
    port map (
            O => \N__16901\,
            I => \N__16882\
        );

    \I__3355\ : LocalMux
    port map (
            O => \N__16896\,
            I => \N__16872\
        );

    \I__3354\ : LocalMux
    port map (
            O => \N__16889\,
            I => \N__16867\
        );

    \I__3353\ : LocalMux
    port map (
            O => \N__16882\,
            I => \N__16867\
        );

    \I__3352\ : CascadeMux
    port map (
            O => \N__16881\,
            I => \N__16864\
        );

    \I__3351\ : CascadeMux
    port map (
            O => \N__16880\,
            I => \N__16860\
        );

    \I__3350\ : CascadeMux
    port map (
            O => \N__16879\,
            I => \N__16857\
        );

    \I__3349\ : CascadeMux
    port map (
            O => \N__16878\,
            I => \N__16854\
        );

    \I__3348\ : CascadeMux
    port map (
            O => \N__16877\,
            I => \N__16850\
        );

    \I__3347\ : CascadeMux
    port map (
            O => \N__16876\,
            I => \N__16847\
        );

    \I__3346\ : CascadeMux
    port map (
            O => \N__16875\,
            I => \N__16844\
        );

    \I__3345\ : Span4Mux_v
    port map (
            O => \N__16872\,
            I => \N__16838\
        );

    \I__3344\ : Span4Mux_h
    port map (
            O => \N__16867\,
            I => \N__16838\
        );

    \I__3343\ : InMux
    port map (
            O => \N__16864\,
            I => \N__16833\
        );

    \I__3342\ : InMux
    port map (
            O => \N__16863\,
            I => \N__16833\
        );

    \I__3341\ : InMux
    port map (
            O => \N__16860\,
            I => \N__16826\
        );

    \I__3340\ : InMux
    port map (
            O => \N__16857\,
            I => \N__16826\
        );

    \I__3339\ : InMux
    port map (
            O => \N__16854\,
            I => \N__16826\
        );

    \I__3338\ : InMux
    port map (
            O => \N__16853\,
            I => \N__16823\
        );

    \I__3337\ : InMux
    port map (
            O => \N__16850\,
            I => \N__16816\
        );

    \I__3336\ : InMux
    port map (
            O => \N__16847\,
            I => \N__16816\
        );

    \I__3335\ : InMux
    port map (
            O => \N__16844\,
            I => \N__16816\
        );

    \I__3334\ : InMux
    port map (
            O => \N__16843\,
            I => \N__16813\
        );

    \I__3333\ : Odrv4
    port map (
            O => \N__16838\,
            I => \ppm_encoder_1.N_241\
        );

    \I__3332\ : LocalMux
    port map (
            O => \N__16833\,
            I => \ppm_encoder_1.N_241\
        );

    \I__3331\ : LocalMux
    port map (
            O => \N__16826\,
            I => \ppm_encoder_1.N_241\
        );

    \I__3330\ : LocalMux
    port map (
            O => \N__16823\,
            I => \ppm_encoder_1.N_241\
        );

    \I__3329\ : LocalMux
    port map (
            O => \N__16816\,
            I => \ppm_encoder_1.N_241\
        );

    \I__3328\ : LocalMux
    port map (
            O => \N__16813\,
            I => \ppm_encoder_1.N_241\
        );

    \I__3327\ : CascadeMux
    port map (
            O => \N__16800\,
            I => \N__16783\
        );

    \I__3326\ : InMux
    port map (
            O => \N__16799\,
            I => \N__16767\
        );

    \I__3325\ : InMux
    port map (
            O => \N__16798\,
            I => \N__16767\
        );

    \I__3324\ : InMux
    port map (
            O => \N__16797\,
            I => \N__16767\
        );

    \I__3323\ : InMux
    port map (
            O => \N__16796\,
            I => \N__16767\
        );

    \I__3322\ : InMux
    port map (
            O => \N__16795\,
            I => \N__16767\
        );

    \I__3321\ : InMux
    port map (
            O => \N__16794\,
            I => \N__16767\
        );

    \I__3320\ : InMux
    port map (
            O => \N__16793\,
            I => \N__16762\
        );

    \I__3319\ : InMux
    port map (
            O => \N__16792\,
            I => \N__16762\
        );

    \I__3318\ : InMux
    port map (
            O => \N__16791\,
            I => \N__16759\
        );

    \I__3317\ : InMux
    port map (
            O => \N__16790\,
            I => \N__16748\
        );

    \I__3316\ : InMux
    port map (
            O => \N__16789\,
            I => \N__16748\
        );

    \I__3315\ : InMux
    port map (
            O => \N__16788\,
            I => \N__16748\
        );

    \I__3314\ : InMux
    port map (
            O => \N__16787\,
            I => \N__16748\
        );

    \I__3313\ : InMux
    port map (
            O => \N__16786\,
            I => \N__16748\
        );

    \I__3312\ : InMux
    port map (
            O => \N__16783\,
            I => \N__16739\
        );

    \I__3311\ : InMux
    port map (
            O => \N__16782\,
            I => \N__16739\
        );

    \I__3310\ : InMux
    port map (
            O => \N__16781\,
            I => \N__16739\
        );

    \I__3309\ : InMux
    port map (
            O => \N__16780\,
            I => \N__16739\
        );

    \I__3308\ : LocalMux
    port map (
            O => \N__16767\,
            I => \N__16736\
        );

    \I__3307\ : LocalMux
    port map (
            O => \N__16762\,
            I => \N__16733\
        );

    \I__3306\ : LocalMux
    port map (
            O => \N__16759\,
            I => \ppm_encoder_1.N_348\
        );

    \I__3305\ : LocalMux
    port map (
            O => \N__16748\,
            I => \ppm_encoder_1.N_348\
        );

    \I__3304\ : LocalMux
    port map (
            O => \N__16739\,
            I => \ppm_encoder_1.N_348\
        );

    \I__3303\ : Odrv4
    port map (
            O => \N__16736\,
            I => \ppm_encoder_1.N_348\
        );

    \I__3302\ : Odrv12
    port map (
            O => \N__16733\,
            I => \ppm_encoder_1.N_348\
        );

    \I__3301\ : InMux
    port map (
            O => \N__16722\,
            I => \N__16719\
        );

    \I__3300\ : LocalMux
    port map (
            O => \N__16719\,
            I => \N__16716\
        );

    \I__3299\ : Span4Mux_v
    port map (
            O => \N__16716\,
            I => \N__16713\
        );

    \I__3298\ : Odrv4
    port map (
            O => \N__16713\,
            I => \ppm_encoder_1.un1_init_pulses_10_8\
        );

    \I__3297\ : InMux
    port map (
            O => \N__16710\,
            I => \N__16707\
        );

    \I__3296\ : LocalMux
    port map (
            O => \N__16707\,
            I => \N__16704\
        );

    \I__3295\ : Span12Mux_v
    port map (
            O => \N__16704\,
            I => \N__16701\
        );

    \I__3294\ : Odrv12
    port map (
            O => \N__16701\,
            I => \ppm_encoder_1.un1_rudder_cry_7_THRU_CO\
        );

    \I__3293\ : InMux
    port map (
            O => \N__16698\,
            I => \N__16695\
        );

    \I__3292\ : LocalMux
    port map (
            O => \N__16695\,
            I => \N__16692\
        );

    \I__3291\ : Span4Mux_h
    port map (
            O => \N__16692\,
            I => \N__16689\
        );

    \I__3290\ : Span4Mux_v
    port map (
            O => \N__16689\,
            I => \N__16685\
        );

    \I__3289\ : InMux
    port map (
            O => \N__16688\,
            I => \N__16682\
        );

    \I__3288\ : Span4Mux_h
    port map (
            O => \N__16685\,
            I => \N__16677\
        );

    \I__3287\ : LocalMux
    port map (
            O => \N__16682\,
            I => \N__16677\
        );

    \I__3286\ : Odrv4
    port map (
            O => \N__16677\,
            I => scaler_4_data_8
        );

    \I__3285\ : InMux
    port map (
            O => \N__16674\,
            I => \N__16671\
        );

    \I__3284\ : LocalMux
    port map (
            O => \N__16671\,
            I => \N__16668\
        );

    \I__3283\ : Span4Mux_h
    port map (
            O => \N__16668\,
            I => \N__16665\
        );

    \I__3282\ : Span4Mux_v
    port map (
            O => \N__16665\,
            I => \N__16662\
        );

    \I__3281\ : Span4Mux_v
    port map (
            O => \N__16662\,
            I => \N__16659\
        );

    \I__3280\ : Odrv4
    port map (
            O => \N__16659\,
            I => \ppm_encoder_1.un1_throttle_cry_6_THRU_CO\
        );

    \I__3279\ : InMux
    port map (
            O => \N__16656\,
            I => \N__16653\
        );

    \I__3278\ : LocalMux
    port map (
            O => \N__16653\,
            I => \N__16650\
        );

    \I__3277\ : Span12Mux_v
    port map (
            O => \N__16650\,
            I => \N__16646\
        );

    \I__3276\ : InMux
    port map (
            O => \N__16649\,
            I => \N__16643\
        );

    \I__3275\ : Odrv12
    port map (
            O => \N__16646\,
            I => scaler_1_data_7
        );

    \I__3274\ : LocalMux
    port map (
            O => \N__16643\,
            I => scaler_1_data_7
        );

    \I__3273\ : InMux
    port map (
            O => \N__16638\,
            I => \N__16635\
        );

    \I__3272\ : LocalMux
    port map (
            O => \N__16635\,
            I => \N__16632\
        );

    \I__3271\ : Sp12to4
    port map (
            O => \N__16632\,
            I => \N__16629\
        );

    \I__3270\ : Span12Mux_v
    port map (
            O => \N__16629\,
            I => \N__16626\
        );

    \I__3269\ : Odrv12
    port map (
            O => \N__16626\,
            I => \ppm_encoder_1.un1_rudder_cry_6_THRU_CO\
        );

    \I__3268\ : InMux
    port map (
            O => \N__16623\,
            I => \N__16620\
        );

    \I__3267\ : LocalMux
    port map (
            O => \N__16620\,
            I => \N__16617\
        );

    \I__3266\ : Span4Mux_h
    port map (
            O => \N__16617\,
            I => \N__16614\
        );

    \I__3265\ : Span4Mux_v
    port map (
            O => \N__16614\,
            I => \N__16610\
        );

    \I__3264\ : InMux
    port map (
            O => \N__16613\,
            I => \N__16607\
        );

    \I__3263\ : Span4Mux_h
    port map (
            O => \N__16610\,
            I => \N__16602\
        );

    \I__3262\ : LocalMux
    port map (
            O => \N__16607\,
            I => \N__16602\
        );

    \I__3261\ : Odrv4
    port map (
            O => \N__16602\,
            I => scaler_4_data_7
        );

    \I__3260\ : CascadeMux
    port map (
            O => \N__16599\,
            I => \ppm_encoder_1.un2_throttle_iv_0_sn_7_cascade_\
        );

    \I__3259\ : InMux
    port map (
            O => \N__16596\,
            I => \N__16593\
        );

    \I__3258\ : LocalMux
    port map (
            O => \N__16593\,
            I => \N__16590\
        );

    \I__3257\ : Odrv4
    port map (
            O => \N__16590\,
            I => \ppm_encoder_1.un1_init_pulses_10_10\
        );

    \I__3256\ : InMux
    port map (
            O => \N__16587\,
            I => \N__16584\
        );

    \I__3255\ : LocalMux
    port map (
            O => \N__16584\,
            I => \N__16581\
        );

    \I__3254\ : Odrv4
    port map (
            O => \N__16581\,
            I => \ppm_encoder_1.un1_init_pulses_10_11\
        );

    \I__3253\ : InMux
    port map (
            O => \N__16578\,
            I => \N__16575\
        );

    \I__3252\ : LocalMux
    port map (
            O => \N__16575\,
            I => \N__16572\
        );

    \I__3251\ : Odrv4
    port map (
            O => \N__16572\,
            I => \ppm_encoder_1.un1_init_pulses_10_12\
        );

    \I__3250\ : InMux
    port map (
            O => \N__16569\,
            I => \N__16566\
        );

    \I__3249\ : LocalMux
    port map (
            O => \N__16566\,
            I => \N__16563\
        );

    \I__3248\ : Span4Mux_v
    port map (
            O => \N__16563\,
            I => \N__16560\
        );

    \I__3247\ : Odrv4
    port map (
            O => \N__16560\,
            I => \ppm_encoder_1.un1_init_pulses_10_2\
        );

    \I__3246\ : CascadeMux
    port map (
            O => \N__16557\,
            I => \N__16554\
        );

    \I__3245\ : InMux
    port map (
            O => \N__16554\,
            I => \N__16551\
        );

    \I__3244\ : LocalMux
    port map (
            O => \N__16551\,
            I => \N__16548\
        );

    \I__3243\ : Span4Mux_v
    port map (
            O => \N__16548\,
            I => \N__16545\
        );

    \I__3242\ : Odrv4
    port map (
            O => \N__16545\,
            I => \ppm_encoder_1.un1_init_pulses_10_3\
        );

    \I__3241\ : InMux
    port map (
            O => \N__16542\,
            I => \N__16539\
        );

    \I__3240\ : LocalMux
    port map (
            O => \N__16539\,
            I => \N__16536\
        );

    \I__3239\ : Span4Mux_v
    port map (
            O => \N__16536\,
            I => \N__16533\
        );

    \I__3238\ : Odrv4
    port map (
            O => \N__16533\,
            I => \ppm_encoder_1.un1_init_pulses_10_5\
        );

    \I__3237\ : InMux
    port map (
            O => \N__16530\,
            I => \N__16527\
        );

    \I__3236\ : LocalMux
    port map (
            O => \N__16527\,
            I => \N__16524\
        );

    \I__3235\ : Span4Mux_v
    port map (
            O => \N__16524\,
            I => \N__16521\
        );

    \I__3234\ : Odrv4
    port map (
            O => \N__16521\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_13\
        );

    \I__3233\ : InMux
    port map (
            O => \N__16518\,
            I => \N__16515\
        );

    \I__3232\ : LocalMux
    port map (
            O => \N__16515\,
            I => \N__16512\
        );

    \I__3231\ : Odrv4
    port map (
            O => \N__16512\,
            I => \ppm_encoder_1.un1_init_pulses_10_13\
        );

    \I__3230\ : InMux
    port map (
            O => \N__16509\,
            I => \N__16506\
        );

    \I__3229\ : LocalMux
    port map (
            O => \N__16506\,
            I => \ppm_encoder_1.un1_init_pulses_10_17\
        );

    \I__3228\ : InMux
    port map (
            O => \N__16503\,
            I => \N__16500\
        );

    \I__3227\ : LocalMux
    port map (
            O => \N__16500\,
            I => \ppm_encoder_1.un1_init_pulses_10_18\
        );

    \I__3226\ : InMux
    port map (
            O => \N__16497\,
            I => \N__16494\
        );

    \I__3225\ : LocalMux
    port map (
            O => \N__16494\,
            I => \N__16491\
        );

    \I__3224\ : Span4Mux_v
    port map (
            O => \N__16491\,
            I => \N__16488\
        );

    \I__3223\ : Odrv4
    port map (
            O => \N__16488\,
            I => \ppm_encoder_1.un1_init_pulses_10_1\
        );

    \I__3222\ : InMux
    port map (
            O => \N__16485\,
            I => \N__16482\
        );

    \I__3221\ : LocalMux
    port map (
            O => \N__16482\,
            I => \N__16479\
        );

    \I__3220\ : Odrv4
    port map (
            O => \N__16479\,
            I => \ppm_encoder_1.un1_init_pulses_10_15\
        );

    \I__3219\ : InMux
    port map (
            O => \N__16476\,
            I => \N__16473\
        );

    \I__3218\ : LocalMux
    port map (
            O => \N__16473\,
            I => \N__16469\
        );

    \I__3217\ : InMux
    port map (
            O => \N__16472\,
            I => \N__16466\
        );

    \I__3216\ : Odrv4
    port map (
            O => \N__16469\,
            I => \ppm_encoder_1.N_245_i_i\
        );

    \I__3215\ : LocalMux
    port map (
            O => \N__16466\,
            I => \ppm_encoder_1.N_245_i_i\
        );

    \I__3214\ : InMux
    port map (
            O => \N__16461\,
            I => \N__16458\
        );

    \I__3213\ : LocalMux
    port map (
            O => \N__16458\,
            I => \N__16455\
        );

    \I__3212\ : Span4Mux_v
    port map (
            O => \N__16455\,
            I => \N__16452\
        );

    \I__3211\ : Odrv4
    port map (
            O => \N__16452\,
            I => \ppm_encoder_1.un1_init_pulses_10_9\
        );

    \I__3210\ : InMux
    port map (
            O => \N__16449\,
            I => \N__16445\
        );

    \I__3209\ : CascadeMux
    port map (
            O => \N__16448\,
            I => \N__16442\
        );

    \I__3208\ : LocalMux
    port map (
            O => \N__16445\,
            I => \N__16439\
        );

    \I__3207\ : InMux
    port map (
            O => \N__16442\,
            I => \N__16436\
        );

    \I__3206\ : Span4Mux_h
    port map (
            O => \N__16439\,
            I => \N__16433\
        );

    \I__3205\ : LocalMux
    port map (
            O => \N__16436\,
            I => \ppm_encoder_1.N_251_i_i\
        );

    \I__3204\ : Odrv4
    port map (
            O => \N__16433\,
            I => \ppm_encoder_1.N_251_i_i\
        );

    \I__3203\ : InMux
    port map (
            O => \N__16428\,
            I => \N__16425\
        );

    \I__3202\ : LocalMux
    port map (
            O => \N__16425\,
            I => \N__16422\
        );

    \I__3201\ : Odrv12
    port map (
            O => \N__16422\,
            I => \ppm_encoder_1.aileronZ0Z_14\
        );

    \I__3200\ : CascadeMux
    port map (
            O => \N__16419\,
            I => \N__16416\
        );

    \I__3199\ : InMux
    port map (
            O => \N__16416\,
            I => \N__16413\
        );

    \I__3198\ : LocalMux
    port map (
            O => \N__16413\,
            I => \N__16410\
        );

    \I__3197\ : Span4Mux_h
    port map (
            O => \N__16410\,
            I => \N__16407\
        );

    \I__3196\ : Odrv4
    port map (
            O => \N__16407\,
            I => \ppm_encoder_1.elevatorZ0Z_14\
        );

    \I__3195\ : InMux
    port map (
            O => \N__16404\,
            I => \N__16401\
        );

    \I__3194\ : LocalMux
    port map (
            O => \N__16401\,
            I => \ppm_encoder_1.pulses2count_9_i_o2_0_14\
        );

    \I__3193\ : InMux
    port map (
            O => \N__16398\,
            I => \N__16395\
        );

    \I__3192\ : LocalMux
    port map (
            O => \N__16395\,
            I => \ppm_encoder_1.un2_throttle_iv_0_2_12\
        );

    \I__3191\ : CascadeMux
    port map (
            O => \N__16392\,
            I => \ppm_encoder_1.un1_init_pulses_0_axb_12_cascade_\
        );

    \I__3190\ : InMux
    port map (
            O => \N__16389\,
            I => \N__16386\
        );

    \I__3189\ : LocalMux
    port map (
            O => \N__16386\,
            I => \ppm_encoder_1.init_pulses_RNI5FJB5Z0Z_12\
        );

    \I__3188\ : CascadeMux
    port map (
            O => \N__16383\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_6_cascade_\
        );

    \I__3187\ : InMux
    port map (
            O => \N__16380\,
            I => \N__16377\
        );

    \I__3186\ : LocalMux
    port map (
            O => \N__16377\,
            I => \ppm_encoder_1.init_pulses_RNIUBDK6Z0Z_7\
        );

    \I__3185\ : CascadeMux
    port map (
            O => \N__16374\,
            I => \N__16371\
        );

    \I__3184\ : InMux
    port map (
            O => \N__16371\,
            I => \N__16367\
        );

    \I__3183\ : InMux
    port map (
            O => \N__16370\,
            I => \N__16364\
        );

    \I__3182\ : LocalMux
    port map (
            O => \N__16367\,
            I => \N__16360\
        );

    \I__3181\ : LocalMux
    port map (
            O => \N__16364\,
            I => \N__16357\
        );

    \I__3180\ : CascadeMux
    port map (
            O => \N__16363\,
            I => \N__16354\
        );

    \I__3179\ : Span4Mux_h
    port map (
            O => \N__16360\,
            I => \N__16351\
        );

    \I__3178\ : Span4Mux_v
    port map (
            O => \N__16357\,
            I => \N__16348\
        );

    \I__3177\ : InMux
    port map (
            O => \N__16354\,
            I => \N__16345\
        );

    \I__3176\ : Odrv4
    port map (
            O => \N__16351\,
            I => \ppm_encoder_1.N_114\
        );

    \I__3175\ : Odrv4
    port map (
            O => \N__16348\,
            I => \ppm_encoder_1.N_114\
        );

    \I__3174\ : LocalMux
    port map (
            O => \N__16345\,
            I => \ppm_encoder_1.N_114\
        );

    \I__3173\ : InMux
    port map (
            O => \N__16338\,
            I => \N__16335\
        );

    \I__3172\ : LocalMux
    port map (
            O => \N__16335\,
            I => \ppm_encoder_1.un2_throttle_iv_0_1_12\
        );

    \I__3171\ : CascadeMux
    port map (
            O => \N__16332\,
            I => \ppm_encoder_1.N_407_cascade_\
        );

    \I__3170\ : CascadeMux
    port map (
            O => \N__16329\,
            I => \ppm_encoder_1.un1_init_pulses_0_axb_2_1_cascade_\
        );

    \I__3169\ : CascadeMux
    port map (
            O => \N__16326\,
            I => \ppm_encoder_1.un1_init_pulses_0_axb_2_cascade_\
        );

    \I__3168\ : InMux
    port map (
            O => \N__16323\,
            I => \N__16320\
        );

    \I__3167\ : LocalMux
    port map (
            O => \N__16320\,
            I => \ppm_encoder_1.init_pulses_RNIE48O3Z0Z_2\
        );

    \I__3166\ : InMux
    port map (
            O => \N__16317\,
            I => \N__16314\
        );

    \I__3165\ : LocalMux
    port map (
            O => \N__16314\,
            I => \ppm_encoder_1.un2_throttle_iv_0_0_14\
        );

    \I__3164\ : CascadeMux
    port map (
            O => \N__16311\,
            I => \ppm_encoder_1.un1_init_pulses_0_axb_5_cascade_\
        );

    \I__3163\ : InMux
    port map (
            O => \N__16308\,
            I => \N__16305\
        );

    \I__3162\ : LocalMux
    port map (
            O => \N__16305\,
            I => \ppm_encoder_1.init_pulses_RNIT8FS5Z0Z_5\
        );

    \I__3161\ : InMux
    port map (
            O => \N__16302\,
            I => \N__16299\
        );

    \I__3160\ : LocalMux
    port map (
            O => \N__16299\,
            I => \ppm_encoder_1.un1_init_pulses_0_axb_5_1_rn_0\
        );

    \I__3159\ : InMux
    port map (
            O => \N__16296\,
            I => \N__16293\
        );

    \I__3158\ : LocalMux
    port map (
            O => \N__16293\,
            I => \N__16290\
        );

    \I__3157\ : Odrv12
    port map (
            O => \N__16290\,
            I => scaler_2_data_5
        );

    \I__3156\ : InMux
    port map (
            O => \N__16287\,
            I => \N__16284\
        );

    \I__3155\ : LocalMux
    port map (
            O => \N__16284\,
            I => \ppm_encoder_1.aileronZ0Z_5\
        );

    \I__3154\ : InMux
    port map (
            O => \N__16281\,
            I => \N__16278\
        );

    \I__3153\ : LocalMux
    port map (
            O => \N__16278\,
            I => \N__16275\
        );

    \I__3152\ : Span4Mux_h
    port map (
            O => \N__16275\,
            I => \N__16272\
        );

    \I__3151\ : Span4Mux_h
    port map (
            O => \N__16272\,
            I => \N__16269\
        );

    \I__3150\ : Odrv4
    port map (
            O => \N__16269\,
            I => scaler_4_data_5
        );

    \I__3149\ : CEMux
    port map (
            O => \N__16266\,
            I => \N__16263\
        );

    \I__3148\ : LocalMux
    port map (
            O => \N__16263\,
            I => \N__16258\
        );

    \I__3147\ : CEMux
    port map (
            O => \N__16262\,
            I => \N__16255\
        );

    \I__3146\ : CEMux
    port map (
            O => \N__16261\,
            I => \N__16250\
        );

    \I__3145\ : IoSpan4Mux
    port map (
            O => \N__16258\,
            I => \N__16245\
        );

    \I__3144\ : LocalMux
    port map (
            O => \N__16255\,
            I => \N__16245\
        );

    \I__3143\ : CEMux
    port map (
            O => \N__16254\,
            I => \N__16240\
        );

    \I__3142\ : CEMux
    port map (
            O => \N__16253\,
            I => \N__16237\
        );

    \I__3141\ : LocalMux
    port map (
            O => \N__16250\,
            I => \N__16234\
        );

    \I__3140\ : Span4Mux_s1_v
    port map (
            O => \N__16245\,
            I => \N__16231\
        );

    \I__3139\ : CEMux
    port map (
            O => \N__16244\,
            I => \N__16228\
        );

    \I__3138\ : CEMux
    port map (
            O => \N__16243\,
            I => \N__16225\
        );

    \I__3137\ : LocalMux
    port map (
            O => \N__16240\,
            I => \N__16222\
        );

    \I__3136\ : LocalMux
    port map (
            O => \N__16237\,
            I => \N__16215\
        );

    \I__3135\ : Span4Mux_v
    port map (
            O => \N__16234\,
            I => \N__16215\
        );

    \I__3134\ : Span4Mux_v
    port map (
            O => \N__16231\,
            I => \N__16215\
        );

    \I__3133\ : LocalMux
    port map (
            O => \N__16228\,
            I => \N__16212\
        );

    \I__3132\ : LocalMux
    port map (
            O => \N__16225\,
            I => \N__16209\
        );

    \I__3131\ : Span4Mux_v
    port map (
            O => \N__16222\,
            I => \N__16206\
        );

    \I__3130\ : Span4Mux_h
    port map (
            O => \N__16215\,
            I => \N__16203\
        );

    \I__3129\ : Span4Mux_v
    port map (
            O => \N__16212\,
            I => \N__16200\
        );

    \I__3128\ : Span4Mux_h
    port map (
            O => \N__16209\,
            I => \N__16193\
        );

    \I__3127\ : Span4Mux_h
    port map (
            O => \N__16206\,
            I => \N__16193\
        );

    \I__3126\ : Span4Mux_v
    port map (
            O => \N__16203\,
            I => \N__16193\
        );

    \I__3125\ : Odrv4
    port map (
            O => \N__16200\,
            I => \ppm_encoder_1.scaler_1_dv_0\
        );

    \I__3124\ : Odrv4
    port map (
            O => \N__16193\,
            I => \ppm_encoder_1.scaler_1_dv_0\
        );

    \I__3123\ : CascadeMux
    port map (
            O => \N__16188\,
            I => \N__16185\
        );

    \I__3122\ : InMux
    port map (
            O => \N__16185\,
            I => \N__16181\
        );

    \I__3121\ : InMux
    port map (
            O => \N__16184\,
            I => \N__16178\
        );

    \I__3120\ : LocalMux
    port map (
            O => \N__16181\,
            I => \ppm_encoder_1.N_252_i_i\
        );

    \I__3119\ : LocalMux
    port map (
            O => \N__16178\,
            I => \ppm_encoder_1.N_252_i_i\
        );

    \I__3118\ : InMux
    port map (
            O => \N__16173\,
            I => \N__16170\
        );

    \I__3117\ : LocalMux
    port map (
            O => \N__16170\,
            I => \N__16167\
        );

    \I__3116\ : Odrv4
    port map (
            O => \N__16167\,
            I => \ppm_encoder_1.un1_init_pulses_0_axb_8\
        );

    \I__3115\ : InMux
    port map (
            O => \N__16164\,
            I => \N__16161\
        );

    \I__3114\ : LocalMux
    port map (
            O => \N__16161\,
            I => \ppm_encoder_1.init_pulses_RNITQDQ5Z0Z_8\
        );

    \I__3113\ : CascadeMux
    port map (
            O => \N__16158\,
            I => \ppm_encoder_1.N_235_cascade_\
        );

    \I__3112\ : InMux
    port map (
            O => \N__16155\,
            I => \N__16152\
        );

    \I__3111\ : LocalMux
    port map (
            O => \N__16152\,
            I => \N__16149\
        );

    \I__3110\ : Span4Mux_h
    port map (
            O => \N__16149\,
            I => \N__16146\
        );

    \I__3109\ : Span4Mux_v
    port map (
            O => \N__16146\,
            I => \N__16143\
        );

    \I__3108\ : Odrv4
    port map (
            O => \N__16143\,
            I => \ppm_encoder_1.un1_elevator_cry_7_THRU_CO\
        );

    \I__3107\ : InMux
    port map (
            O => \N__16140\,
            I => \N__16137\
        );

    \I__3106\ : LocalMux
    port map (
            O => \N__16137\,
            I => \N__16134\
        );

    \I__3105\ : Span4Mux_v
    port map (
            O => \N__16134\,
            I => \N__16130\
        );

    \I__3104\ : InMux
    port map (
            O => \N__16133\,
            I => \N__16127\
        );

    \I__3103\ : Span4Mux_v
    port map (
            O => \N__16130\,
            I => \N__16124\
        );

    \I__3102\ : LocalMux
    port map (
            O => \N__16127\,
            I => \N__16121\
        );

    \I__3101\ : Span4Mux_h
    port map (
            O => \N__16124\,
            I => \N__16116\
        );

    \I__3100\ : Span4Mux_v
    port map (
            O => \N__16121\,
            I => \N__16116\
        );

    \I__3099\ : Odrv4
    port map (
            O => \N__16116\,
            I => scaler_3_data_8
        );

    \I__3098\ : InMux
    port map (
            O => \N__16113\,
            I => \N__16110\
        );

    \I__3097\ : LocalMux
    port map (
            O => \N__16110\,
            I => \N__16107\
        );

    \I__3096\ : Span4Mux_h
    port map (
            O => \N__16107\,
            I => \N__16104\
        );

    \I__3095\ : Span4Mux_h
    port map (
            O => \N__16104\,
            I => \N__16101\
        );

    \I__3094\ : Odrv4
    port map (
            O => \N__16101\,
            I => scaler_3_data_5
        );

    \I__3093\ : InMux
    port map (
            O => \N__16098\,
            I => \N__16095\
        );

    \I__3092\ : LocalMux
    port map (
            O => \N__16095\,
            I => \N__16092\
        );

    \I__3091\ : Span4Mux_h
    port map (
            O => \N__16092\,
            I => \N__16088\
        );

    \I__3090\ : CascadeMux
    port map (
            O => \N__16091\,
            I => \N__16085\
        );

    \I__3089\ : Span4Mux_h
    port map (
            O => \N__16088\,
            I => \N__16082\
        );

    \I__3088\ : InMux
    port map (
            O => \N__16085\,
            I => \N__16079\
        );

    \I__3087\ : Odrv4
    port map (
            O => \N__16082\,
            I => scaler_4_data_4
        );

    \I__3086\ : LocalMux
    port map (
            O => \N__16079\,
            I => scaler_4_data_4
        );

    \I__3085\ : InMux
    port map (
            O => \N__16074\,
            I => \N__16071\
        );

    \I__3084\ : LocalMux
    port map (
            O => \N__16071\,
            I => \N__16068\
        );

    \I__3083\ : Span4Mux_h
    port map (
            O => \N__16068\,
            I => \N__16064\
        );

    \I__3082\ : CascadeMux
    port map (
            O => \N__16067\,
            I => \N__16061\
        );

    \I__3081\ : Span4Mux_h
    port map (
            O => \N__16064\,
            I => \N__16058\
        );

    \I__3080\ : InMux
    port map (
            O => \N__16061\,
            I => \N__16055\
        );

    \I__3079\ : Odrv4
    port map (
            O => \N__16058\,
            I => scaler_1_data_4
        );

    \I__3078\ : LocalMux
    port map (
            O => \N__16055\,
            I => scaler_1_data_4
        );

    \I__3077\ : InMux
    port map (
            O => \N__16050\,
            I => \N__16047\
        );

    \I__3076\ : LocalMux
    port map (
            O => \N__16047\,
            I => \N__16044\
        );

    \I__3075\ : Span12Mux_h
    port map (
            O => \N__16044\,
            I => \N__16041\
        );

    \I__3074\ : Odrv12
    port map (
            O => \N__16041\,
            I => scaler_1_data_5
        );

    \I__3073\ : CascadeMux
    port map (
            O => \N__16038\,
            I => \N__16035\
        );

    \I__3072\ : InMux
    port map (
            O => \N__16035\,
            I => \N__16032\
        );

    \I__3071\ : LocalMux
    port map (
            O => \N__16032\,
            I => \ppm_encoder_1.elevatorZ0Z_5\
        );

    \I__3070\ : CascadeMux
    port map (
            O => \N__16029\,
            I => \ppm_encoder_1.un1_init_pulses_0_axb_5_1_sn_cascade_\
        );

    \I__3069\ : CascadeMux
    port map (
            O => \N__16026\,
            I => \ppm_encoder_1.un1_init_pulses_0_axb_5_1_cascade_\
        );

    \I__3068\ : InMux
    port map (
            O => \N__16023\,
            I => \N__16020\
        );

    \I__3067\ : LocalMux
    port map (
            O => \N__16020\,
            I => \N__16017\
        );

    \I__3066\ : Span4Mux_h
    port map (
            O => \N__16017\,
            I => \N__16013\
        );

    \I__3065\ : InMux
    port map (
            O => \N__16016\,
            I => \N__16010\
        );

    \I__3064\ : Odrv4
    port map (
            O => \N__16013\,
            I => scaler_1_data_11
        );

    \I__3063\ : LocalMux
    port map (
            O => \N__16010\,
            I => scaler_1_data_11
        );

    \I__3062\ : InMux
    port map (
            O => \N__16005\,
            I => \N__16002\
        );

    \I__3061\ : LocalMux
    port map (
            O => \N__16002\,
            I => \N__15999\
        );

    \I__3060\ : Odrv4
    port map (
            O => \N__15999\,
            I => \ppm_encoder_1.un1_throttle_cry_10_THRU_CO\
        );

    \I__3059\ : InMux
    port map (
            O => \N__15996\,
            I => \N__15993\
        );

    \I__3058\ : LocalMux
    port map (
            O => \N__15993\,
            I => \N__15989\
        );

    \I__3057\ : CascadeMux
    port map (
            O => \N__15992\,
            I => \N__15986\
        );

    \I__3056\ : Span4Mux_v
    port map (
            O => \N__15989\,
            I => \N__15983\
        );

    \I__3055\ : InMux
    port map (
            O => \N__15986\,
            I => \N__15980\
        );

    \I__3054\ : Span4Mux_h
    port map (
            O => \N__15983\,
            I => \N__15975\
        );

    \I__3053\ : LocalMux
    port map (
            O => \N__15980\,
            I => \N__15975\
        );

    \I__3052\ : Odrv4
    port map (
            O => \N__15975\,
            I => scaler_2_data_12
        );

    \I__3051\ : InMux
    port map (
            O => \N__15972\,
            I => \N__15969\
        );

    \I__3050\ : LocalMux
    port map (
            O => \N__15969\,
            I => \N__15966\
        );

    \I__3049\ : Span4Mux_v
    port map (
            O => \N__15966\,
            I => \N__15963\
        );

    \I__3048\ : Span4Mux_h
    port map (
            O => \N__15963\,
            I => \N__15960\
        );

    \I__3047\ : Odrv4
    port map (
            O => \N__15960\,
            I => \ppm_encoder_1.un1_aileron_cry_11_THRU_CO\
        );

    \I__3046\ : InMux
    port map (
            O => \N__15957\,
            I => \N__15954\
        );

    \I__3045\ : LocalMux
    port map (
            O => \N__15954\,
            I => \ppm_encoder_1.N_418\
        );

    \I__3044\ : CascadeMux
    port map (
            O => \N__15951\,
            I => \ppm_encoder_1.N_417_cascade_\
        );

    \I__3043\ : CascadeMux
    port map (
            O => \N__15948\,
            I => \ppm_encoder_1.un2_throttle_iv_0_1_8_cascade_\
        );

    \I__3042\ : InMux
    port map (
            O => \N__15945\,
            I => \N__15942\
        );

    \I__3041\ : LocalMux
    port map (
            O => \N__15942\,
            I => \N__15939\
        );

    \I__3040\ : Span4Mux_h
    port map (
            O => \N__15939\,
            I => \N__15936\
        );

    \I__3039\ : Odrv4
    port map (
            O => \N__15936\,
            I => \ppm_encoder_1.un1_aileron_cry_7_THRU_CO\
        );

    \I__3038\ : InMux
    port map (
            O => \N__15933\,
            I => \N__15930\
        );

    \I__3037\ : LocalMux
    port map (
            O => \N__15930\,
            I => \N__15926\
        );

    \I__3036\ : InMux
    port map (
            O => \N__15929\,
            I => \N__15923\
        );

    \I__3035\ : Span12Mux_h
    port map (
            O => \N__15926\,
            I => \N__15920\
        );

    \I__3034\ : LocalMux
    port map (
            O => \N__15923\,
            I => \N__15917\
        );

    \I__3033\ : Odrv12
    port map (
            O => \N__15920\,
            I => scaler_2_data_8
        );

    \I__3032\ : Odrv4
    port map (
            O => \N__15917\,
            I => scaler_2_data_8
        );

    \I__3031\ : InMux
    port map (
            O => \N__15912\,
            I => \N__15909\
        );

    \I__3030\ : LocalMux
    port map (
            O => \N__15909\,
            I => \N__15906\
        );

    \I__3029\ : Span4Mux_h
    port map (
            O => \N__15906\,
            I => \N__15903\
        );

    \I__3028\ : Span4Mux_v
    port map (
            O => \N__15903\,
            I => \N__15900\
        );

    \I__3027\ : Span4Mux_v
    port map (
            O => \N__15900\,
            I => \N__15897\
        );

    \I__3026\ : Odrv4
    port map (
            O => \N__15897\,
            I => \ppm_encoder_1.un1_throttle_cry_7_THRU_CO\
        );

    \I__3025\ : CascadeMux
    port map (
            O => \N__15894\,
            I => \N__15891\
        );

    \I__3024\ : InMux
    port map (
            O => \N__15891\,
            I => \N__15888\
        );

    \I__3023\ : LocalMux
    port map (
            O => \N__15888\,
            I => \N__15885\
        );

    \I__3022\ : Span4Mux_h
    port map (
            O => \N__15885\,
            I => \N__15882\
        );

    \I__3021\ : Span4Mux_v
    port map (
            O => \N__15882\,
            I => \N__15879\
        );

    \I__3020\ : Span4Mux_h
    port map (
            O => \N__15879\,
            I => \N__15875\
        );

    \I__3019\ : InMux
    port map (
            O => \N__15878\,
            I => \N__15872\
        );

    \I__3018\ : Odrv4
    port map (
            O => \N__15875\,
            I => scaler_1_data_8
        );

    \I__3017\ : LocalMux
    port map (
            O => \N__15872\,
            I => scaler_1_data_8
        );

    \I__3016\ : CascadeMux
    port map (
            O => \N__15867\,
            I => \N__15863\
        );

    \I__3015\ : InMux
    port map (
            O => \N__15866\,
            I => \N__15860\
        );

    \I__3014\ : InMux
    port map (
            O => \N__15863\,
            I => \N__15857\
        );

    \I__3013\ : LocalMux
    port map (
            O => \N__15860\,
            I => \N__15854\
        );

    \I__3012\ : LocalMux
    port map (
            O => \N__15857\,
            I => \ppm_encoder_1.throttleZ0Z_13\
        );

    \I__3011\ : Odrv4
    port map (
            O => \N__15854\,
            I => \ppm_encoder_1.throttleZ0Z_13\
        );

    \I__3010\ : CascadeMux
    port map (
            O => \N__15849\,
            I => \ppm_encoder_1.pulses2count_9_0_o2_0_13_cascade_\
        );

    \I__3009\ : InMux
    port map (
            O => \N__15846\,
            I => \N__15843\
        );

    \I__3008\ : LocalMux
    port map (
            O => \N__15843\,
            I => \N__15840\
        );

    \I__3007\ : Span4Mux_v
    port map (
            O => \N__15840\,
            I => \N__15836\
        );

    \I__3006\ : InMux
    port map (
            O => \N__15839\,
            I => \N__15833\
        );

    \I__3005\ : Span4Mux_h
    port map (
            O => \N__15836\,
            I => \N__15830\
        );

    \I__3004\ : LocalMux
    port map (
            O => \N__15833\,
            I => \N__15827\
        );

    \I__3003\ : Odrv4
    port map (
            O => \N__15830\,
            I => scaler_2_data_13
        );

    \I__3002\ : Odrv4
    port map (
            O => \N__15827\,
            I => scaler_2_data_13
        );

    \I__3001\ : InMux
    port map (
            O => \N__15822\,
            I => \N__15819\
        );

    \I__3000\ : LocalMux
    port map (
            O => \N__15819\,
            I => \N__15816\
        );

    \I__2999\ : Span4Mux_s3_v
    port map (
            O => \N__15816\,
            I => \N__15813\
        );

    \I__2998\ : Span4Mux_h
    port map (
            O => \N__15813\,
            I => \N__15810\
        );

    \I__2997\ : Odrv4
    port map (
            O => \N__15810\,
            I => \ppm_encoder_1.un1_aileron_cry_12_THRU_CO\
        );

    \I__2996\ : InMux
    port map (
            O => \N__15807\,
            I => \N__15801\
        );

    \I__2995\ : InMux
    port map (
            O => \N__15806\,
            I => \N__15801\
        );

    \I__2994\ : LocalMux
    port map (
            O => \N__15801\,
            I => \ppm_encoder_1.aileronZ0Z_13\
        );

    \I__2993\ : CascadeMux
    port map (
            O => \N__15798\,
            I => \ppm_encoder_1.un2_throttle_iv_0_0_13_cascade_\
        );

    \I__2992\ : CascadeMux
    port map (
            O => \N__15795\,
            I => \ppm_encoder_1.un1_init_pulses_0_axb_13_cascade_\
        );

    \I__2991\ : CascadeMux
    port map (
            O => \N__15792\,
            I => \N__15789\
        );

    \I__2990\ : InMux
    port map (
            O => \N__15789\,
            I => \N__15786\
        );

    \I__2989\ : LocalMux
    port map (
            O => \N__15786\,
            I => \N__15783\
        );

    \I__2988\ : Odrv12
    port map (
            O => \N__15783\,
            I => \ppm_encoder_1.init_pulses_RNIC11J5Z0Z_13\
        );

    \I__2987\ : InMux
    port map (
            O => \N__15780\,
            I => \N__15777\
        );

    \I__2986\ : LocalMux
    port map (
            O => \N__15777\,
            I => \N__15773\
        );

    \I__2985\ : InMux
    port map (
            O => \N__15776\,
            I => \N__15770\
        );

    \I__2984\ : Span4Mux_h
    port map (
            O => \N__15773\,
            I => \N__15767\
        );

    \I__2983\ : LocalMux
    port map (
            O => \N__15770\,
            I => \N__15764\
        );

    \I__2982\ : Span4Mux_h
    port map (
            O => \N__15767\,
            I => \N__15761\
        );

    \I__2981\ : Span4Mux_h
    port map (
            O => \N__15764\,
            I => \N__15758\
        );

    \I__2980\ : Odrv4
    port map (
            O => \N__15761\,
            I => scaler_3_data_13
        );

    \I__2979\ : Odrv4
    port map (
            O => \N__15758\,
            I => scaler_3_data_13
        );

    \I__2978\ : InMux
    port map (
            O => \N__15753\,
            I => \N__15750\
        );

    \I__2977\ : LocalMux
    port map (
            O => \N__15750\,
            I => \N__15747\
        );

    \I__2976\ : Span4Mux_h
    port map (
            O => \N__15747\,
            I => \N__15744\
        );

    \I__2975\ : Odrv4
    port map (
            O => \N__15744\,
            I => \ppm_encoder_1.un1_elevator_cry_12_THRU_CO\
        );

    \I__2974\ : CascadeMux
    port map (
            O => \N__15741\,
            I => \N__15737\
        );

    \I__2973\ : InMux
    port map (
            O => \N__15740\,
            I => \N__15732\
        );

    \I__2972\ : InMux
    port map (
            O => \N__15737\,
            I => \N__15732\
        );

    \I__2971\ : LocalMux
    port map (
            O => \N__15732\,
            I => \ppm_encoder_1.elevatorZ0Z_13\
        );

    \I__2970\ : InMux
    port map (
            O => \N__15729\,
            I => \N__15726\
        );

    \I__2969\ : LocalMux
    port map (
            O => \N__15726\,
            I => \N__15723\
        );

    \I__2968\ : Odrv12
    port map (
            O => \N__15723\,
            I => \ppm_encoder_1.un2_throttle_iv_0_1_11\
        );

    \I__2967\ : InMux
    port map (
            O => \N__15720\,
            I => \N__15717\
        );

    \I__2966\ : LocalMux
    port map (
            O => \N__15717\,
            I => \N__15713\
        );

    \I__2965\ : InMux
    port map (
            O => \N__15716\,
            I => \N__15710\
        );

    \I__2964\ : Span4Mux_h
    port map (
            O => \N__15713\,
            I => \N__15707\
        );

    \I__2963\ : LocalMux
    port map (
            O => \N__15710\,
            I => \N__15704\
        );

    \I__2962\ : Span4Mux_v
    port map (
            O => \N__15707\,
            I => \N__15701\
        );

    \I__2961\ : Span4Mux_h
    port map (
            O => \N__15704\,
            I => \N__15698\
        );

    \I__2960\ : Odrv4
    port map (
            O => \N__15701\,
            I => scaler_3_data_11
        );

    \I__2959\ : Odrv4
    port map (
            O => \N__15698\,
            I => scaler_3_data_11
        );

    \I__2958\ : CascadeMux
    port map (
            O => \N__15693\,
            I => \N__15690\
        );

    \I__2957\ : InMux
    port map (
            O => \N__15690\,
            I => \N__15687\
        );

    \I__2956\ : LocalMux
    port map (
            O => \N__15687\,
            I => \N__15684\
        );

    \I__2955\ : Span4Mux_s3_v
    port map (
            O => \N__15684\,
            I => \N__15681\
        );

    \I__2954\ : Odrv4
    port map (
            O => \N__15681\,
            I => \ppm_encoder_1.un1_elevator_cry_10_THRU_CO\
        );

    \I__2953\ : CascadeMux
    port map (
            O => \N__15678\,
            I => \ppm_encoder_1.N_114_cascade_\
        );

    \I__2952\ : InMux
    port map (
            O => \N__15675\,
            I => \N__15670\
        );

    \I__2951\ : InMux
    port map (
            O => \N__15674\,
            I => \N__15667\
        );

    \I__2950\ : InMux
    port map (
            O => \N__15673\,
            I => \N__15664\
        );

    \I__2949\ : LocalMux
    port map (
            O => \N__15670\,
            I => \N__15661\
        );

    \I__2948\ : LocalMux
    port map (
            O => \N__15667\,
            I => \N__15658\
        );

    \I__2947\ : LocalMux
    port map (
            O => \N__15664\,
            I => \ppm_encoder_1.elevatorZ0Z_10\
        );

    \I__2946\ : Odrv4
    port map (
            O => \N__15661\,
            I => \ppm_encoder_1.elevatorZ0Z_10\
        );

    \I__2945\ : Odrv4
    port map (
            O => \N__15658\,
            I => \ppm_encoder_1.elevatorZ0Z_10\
        );

    \I__2944\ : CascadeMux
    port map (
            O => \N__15651\,
            I => \N__15646\
        );

    \I__2943\ : CascadeMux
    port map (
            O => \N__15650\,
            I => \N__15643\
        );

    \I__2942\ : InMux
    port map (
            O => \N__15649\,
            I => \N__15640\
        );

    \I__2941\ : InMux
    port map (
            O => \N__15646\,
            I => \N__15637\
        );

    \I__2940\ : InMux
    port map (
            O => \N__15643\,
            I => \N__15634\
        );

    \I__2939\ : LocalMux
    port map (
            O => \N__15640\,
            I => \N__15629\
        );

    \I__2938\ : LocalMux
    port map (
            O => \N__15637\,
            I => \N__15629\
        );

    \I__2937\ : LocalMux
    port map (
            O => \N__15634\,
            I => \N__15626\
        );

    \I__2936\ : Odrv4
    port map (
            O => \N__15629\,
            I => \ppm_encoder_1.aileronZ0Z_10\
        );

    \I__2935\ : Odrv4
    port map (
            O => \N__15626\,
            I => \ppm_encoder_1.aileronZ0Z_10\
        );

    \I__2934\ : CascadeMux
    port map (
            O => \N__15621\,
            I => \ppm_encoder_1.N_348_cascade_\
        );

    \I__2933\ : InMux
    port map (
            O => \N__15618\,
            I => \N__15615\
        );

    \I__2932\ : LocalMux
    port map (
            O => \N__15615\,
            I => \N__15612\
        );

    \I__2931\ : Odrv4
    port map (
            O => \N__15612\,
            I => \ppm_encoder_1.un1_init_pulses_10_14\
        );

    \I__2930\ : CascadeMux
    port map (
            O => \N__15609\,
            I => \ppm_encoder_1.init_pulses_18_i_0_14_cascade_\
        );

    \I__2929\ : InMux
    port map (
            O => \N__15606\,
            I => \N__15603\
        );

    \I__2928\ : LocalMux
    port map (
            O => \N__15603\,
            I => \ppm_encoder_1.init_pulses_18_i_a2_0_14\
        );

    \I__2927\ : InMux
    port map (
            O => \N__15600\,
            I => \N__15597\
        );

    \I__2926\ : LocalMux
    port map (
            O => \N__15597\,
            I => \N__15594\
        );

    \I__2925\ : Odrv4
    port map (
            O => \N__15594\,
            I => \ppm_encoder_1.un1_init_pulses_10_16\
        );

    \I__2924\ : CascadeMux
    port map (
            O => \N__15591\,
            I => \ppm_encoder_1.N_241_cascade_\
        );

    \I__2923\ : CascadeMux
    port map (
            O => \N__15588\,
            I => \ppm_encoder_1.un1_init_pulses_0_axb_14_cascade_\
        );

    \I__2922\ : CascadeMux
    port map (
            O => \N__15585\,
            I => \N__15582\
        );

    \I__2921\ : InMux
    port map (
            O => \N__15582\,
            I => \N__15579\
        );

    \I__2920\ : LocalMux
    port map (
            O => \N__15579\,
            I => \ppm_encoder_1.init_pulses_RNINK8A6Z0Z_14\
        );

    \I__2919\ : CascadeMux
    port map (
            O => \N__15576\,
            I => \N__15573\
        );

    \I__2918\ : InMux
    port map (
            O => \N__15573\,
            I => \N__15570\
        );

    \I__2917\ : LocalMux
    port map (
            O => \N__15570\,
            I => \N__15567\
        );

    \I__2916\ : Odrv4
    port map (
            O => \N__15567\,
            I => \ppm_encoder_1.init_pulses_RNIJJM71Z0Z_15\
        );

    \I__2915\ : InMux
    port map (
            O => \N__15564\,
            I => \N__15561\
        );

    \I__2914\ : LocalMux
    port map (
            O => \N__15561\,
            I => \N__15558\
        );

    \I__2913\ : Span4Mux_v
    port map (
            O => \N__15558\,
            I => \N__15555\
        );

    \I__2912\ : Odrv4
    port map (
            O => \N__15555\,
            I => \ppm_encoder_1.N_403\
        );

    \I__2911\ : CascadeMux
    port map (
            O => \N__15552\,
            I => \N__15549\
        );

    \I__2910\ : InMux
    port map (
            O => \N__15549\,
            I => \N__15546\
        );

    \I__2909\ : LocalMux
    port map (
            O => \N__15546\,
            I => \N__15543\
        );

    \I__2908\ : Span4Mux_h
    port map (
            O => \N__15543\,
            I => \N__15540\
        );

    \I__2907\ : Odrv4
    port map (
            O => \N__15540\,
            I => \ppm_encoder_1.throttleZ0Z_14\
        );

    \I__2906\ : InMux
    port map (
            O => \N__15537\,
            I => \N__15534\
        );

    \I__2905\ : LocalMux
    port map (
            O => \N__15534\,
            I => \N__15531\
        );

    \I__2904\ : Odrv12
    port map (
            O => \N__15531\,
            I => \ppm_encoder_1.init_pulses_RNIJ2JB5Z0Z_10\
        );

    \I__2903\ : InMux
    port map (
            O => \N__15528\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_9\
        );

    \I__2902\ : InMux
    port map (
            O => \N__15525\,
            I => \N__15522\
        );

    \I__2901\ : LocalMux
    port map (
            O => \N__15522\,
            I => \N__15519\
        );

    \I__2900\ : Odrv12
    port map (
            O => \N__15519\,
            I => \ppm_encoder_1.init_pulses_RNIV8JB5Z0Z_11\
        );

    \I__2899\ : InMux
    port map (
            O => \N__15516\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_10\
        );

    \I__2898\ : InMux
    port map (
            O => \N__15513\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_11\
        );

    \I__2897\ : InMux
    port map (
            O => \N__15510\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_12\
        );

    \I__2896\ : InMux
    port map (
            O => \N__15507\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_13\
        );

    \I__2895\ : InMux
    port map (
            O => \N__15504\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_14\
        );

    \I__2894\ : InMux
    port map (
            O => \N__15501\,
            I => \bfn_7_25_0_\
        );

    \I__2893\ : InMux
    port map (
            O => \N__15498\,
            I => \N__15495\
        );

    \I__2892\ : LocalMux
    port map (
            O => \N__15495\,
            I => \N__15492\
        );

    \I__2891\ : Odrv12
    port map (
            O => \N__15492\,
            I => \ppm_encoder_1.un1_init_pulses_0_axb_17\
        );

    \I__2890\ : InMux
    port map (
            O => \N__15489\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_16\
        );

    \I__2889\ : InMux
    port map (
            O => \N__15486\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_17\
        );

    \I__2888\ : InMux
    port map (
            O => \N__15483\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_1\
        );

    \I__2887\ : InMux
    port map (
            O => \N__15480\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_2\
        );

    \I__2886\ : InMux
    port map (
            O => \N__15477\,
            I => \N__15474\
        );

    \I__2885\ : LocalMux
    port map (
            O => \N__15474\,
            I => \ppm_encoder_1.init_pulses_RNI398E4Z0Z_4\
        );

    \I__2884\ : InMux
    port map (
            O => \N__15471\,
            I => \N__15468\
        );

    \I__2883\ : LocalMux
    port map (
            O => \N__15468\,
            I => \ppm_encoder_1.un1_init_pulses_10_4\
        );

    \I__2882\ : InMux
    port map (
            O => \N__15465\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_3\
        );

    \I__2881\ : InMux
    port map (
            O => \N__15462\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_4\
        );

    \I__2880\ : InMux
    port map (
            O => \N__15459\,
            I => \N__15456\
        );

    \I__2879\ : LocalMux
    port map (
            O => \N__15456\,
            I => \N__15453\
        );

    \I__2878\ : Odrv4
    port map (
            O => \N__15453\,
            I => \ppm_encoder_1.init_pulses_RNI6UPC6Z0Z_6\
        );

    \I__2877\ : InMux
    port map (
            O => \N__15450\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_5\
        );

    \I__2876\ : InMux
    port map (
            O => \N__15447\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_6\
        );

    \I__2875\ : InMux
    port map (
            O => \N__15444\,
            I => \bfn_7_24_0_\
        );

    \I__2874\ : InMux
    port map (
            O => \N__15441\,
            I => \N__15438\
        );

    \I__2873\ : LocalMux
    port map (
            O => \N__15438\,
            I => \N__15435\
        );

    \I__2872\ : Odrv4
    port map (
            O => \N__15435\,
            I => \ppm_encoder_1.init_pulses_RNI31EQ5Z0Z_9\
        );

    \I__2871\ : InMux
    port map (
            O => \N__15432\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_8\
        );

    \I__2870\ : CascadeMux
    port map (
            O => \N__15429\,
            I => \ppm_encoder_1.un1_init_pulses_11_0_cascade_\
        );

    \I__2869\ : InMux
    port map (
            O => \N__15426\,
            I => \N__15423\
        );

    \I__2868\ : LocalMux
    port map (
            O => \N__15423\,
            I => \ppm_encoder_1.un2_throttle_iv_i_i_1_4\
        );

    \I__2867\ : CascadeMux
    port map (
            O => \N__15420\,
            I => \ppm_encoder_1.un1_init_pulses_0_axb_4_cascade_\
        );

    \I__2866\ : InMux
    port map (
            O => \N__15417\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_0\
        );

    \I__2865\ : InMux
    port map (
            O => \N__15414\,
            I => \N__15411\
        );

    \I__2864\ : LocalMux
    port map (
            O => \N__15411\,
            I => \N__15407\
        );

    \I__2863\ : IoInMux
    port map (
            O => \N__15410\,
            I => \N__15404\
        );

    \I__2862\ : Span4Mux_h
    port map (
            O => \N__15407\,
            I => \N__15401\
        );

    \I__2861\ : LocalMux
    port map (
            O => \N__15404\,
            I => \N__15398\
        );

    \I__2860\ : Span4Mux_v
    port map (
            O => \N__15401\,
            I => \N__15395\
        );

    \I__2859\ : IoSpan4Mux
    port map (
            O => \N__15398\,
            I => \N__15392\
        );

    \I__2858\ : Odrv4
    port map (
            O => \N__15395\,
            I => uart_input_c
        );

    \I__2857\ : Odrv4
    port map (
            O => \N__15392\,
            I => uart_input_c
        );

    \I__2856\ : InMux
    port map (
            O => \N__15387\,
            I => \N__15384\
        );

    \I__2855\ : LocalMux
    port map (
            O => \N__15384\,
            I => \N__15381\
        );

    \I__2854\ : Span4Mux_v
    port map (
            O => \N__15381\,
            I => \N__15378\
        );

    \I__2853\ : Odrv4
    port map (
            O => \N__15378\,
            I => \uart_sync.aux_0__0_Z0Z_0\
        );

    \I__2852\ : InMux
    port map (
            O => \N__15375\,
            I => \N__15372\
        );

    \I__2851\ : LocalMux
    port map (
            O => \N__15372\,
            I => \N__15368\
        );

    \I__2850\ : InMux
    port map (
            O => \N__15371\,
            I => \N__15364\
        );

    \I__2849\ : Span4Mux_h
    port map (
            O => \N__15368\,
            I => \N__15361\
        );

    \I__2848\ : InMux
    port map (
            O => \N__15367\,
            I => \N__15358\
        );

    \I__2847\ : LocalMux
    port map (
            O => \N__15364\,
            I => \ppm_encoder_1.throttleZ0Z_6\
        );

    \I__2846\ : Odrv4
    port map (
            O => \N__15361\,
            I => \ppm_encoder_1.throttleZ0Z_6\
        );

    \I__2845\ : LocalMux
    port map (
            O => \N__15358\,
            I => \ppm_encoder_1.throttleZ0Z_6\
        );

    \I__2844\ : CascadeMux
    port map (
            O => \N__15351\,
            I => \N__15348\
        );

    \I__2843\ : InMux
    port map (
            O => \N__15348\,
            I => \N__15345\
        );

    \I__2842\ : LocalMux
    port map (
            O => \N__15345\,
            I => \N__15342\
        );

    \I__2841\ : Span4Mux_h
    port map (
            O => \N__15342\,
            I => \N__15339\
        );

    \I__2840\ : Odrv4
    port map (
            O => \N__15339\,
            I => \ppm_encoder_1.pulses2count_9_0_o2_0_6\
        );

    \I__2839\ : CascadeMux
    port map (
            O => \N__15336\,
            I => \ppm_encoder_1.un1_init_pulses_0_axb_11_cascade_\
        );

    \I__2838\ : InMux
    port map (
            O => \N__15333\,
            I => \N__15330\
        );

    \I__2837\ : LocalMux
    port map (
            O => \N__15330\,
            I => \ppm_encoder_1.un2_throttle_iv_0_2_11\
        );

    \I__2836\ : CascadeMux
    port map (
            O => \N__15327\,
            I => \ppm_encoder_1.un2_throttle_iv_i_i_1_1_4_cascade_\
        );

    \I__2835\ : InMux
    port map (
            O => \N__15324\,
            I => \N__15321\
        );

    \I__2834\ : LocalMux
    port map (
            O => \N__15321\,
            I => \N__15318\
        );

    \I__2833\ : Odrv4
    port map (
            O => \N__15318\,
            I => \ppm_encoder_1.N_462\
        );

    \I__2832\ : InMux
    port map (
            O => \N__15315\,
            I => \N__15312\
        );

    \I__2831\ : LocalMux
    port map (
            O => \N__15312\,
            I => \N__15307\
        );

    \I__2830\ : InMux
    port map (
            O => \N__15311\,
            I => \N__15302\
        );

    \I__2829\ : InMux
    port map (
            O => \N__15310\,
            I => \N__15302\
        );

    \I__2828\ : Odrv4
    port map (
            O => \N__15307\,
            I => \ppm_encoder_1.aileronZ0Z_9\
        );

    \I__2827\ : LocalMux
    port map (
            O => \N__15302\,
            I => \ppm_encoder_1.aileronZ0Z_9\
        );

    \I__2826\ : InMux
    port map (
            O => \N__15297\,
            I => \N__15294\
        );

    \I__2825\ : LocalMux
    port map (
            O => \N__15294\,
            I => \N__15291\
        );

    \I__2824\ : Odrv4
    port map (
            O => \N__15291\,
            I => \ppm_encoder_1.un1_rudder_cry_8_THRU_CO\
        );

    \I__2823\ : InMux
    port map (
            O => \N__15288\,
            I => \N__15285\
        );

    \I__2822\ : LocalMux
    port map (
            O => \N__15285\,
            I => \N__15281\
        );

    \I__2821\ : InMux
    port map (
            O => \N__15284\,
            I => \N__15278\
        );

    \I__2820\ : Span4Mux_v
    port map (
            O => \N__15281\,
            I => \N__15275\
        );

    \I__2819\ : LocalMux
    port map (
            O => \N__15278\,
            I => \N__15272\
        );

    \I__2818\ : Odrv4
    port map (
            O => \N__15275\,
            I => scaler_4_data_9
        );

    \I__2817\ : Odrv4
    port map (
            O => \N__15272\,
            I => scaler_4_data_9
        );

    \I__2816\ : InMux
    port map (
            O => \N__15267\,
            I => \N__15263\
        );

    \I__2815\ : InMux
    port map (
            O => \N__15266\,
            I => \N__15260\
        );

    \I__2814\ : LocalMux
    port map (
            O => \N__15263\,
            I => \N__15257\
        );

    \I__2813\ : LocalMux
    port map (
            O => \N__15260\,
            I => \N__15254\
        );

    \I__2812\ : Span4Mux_v
    port map (
            O => \N__15257\,
            I => \N__15251\
        );

    \I__2811\ : Span4Mux_h
    port map (
            O => \N__15254\,
            I => \N__15248\
        );

    \I__2810\ : Odrv4
    port map (
            O => \N__15251\,
            I => scaler_3_data_10
        );

    \I__2809\ : Odrv4
    port map (
            O => \N__15248\,
            I => scaler_3_data_10
        );

    \I__2808\ : InMux
    port map (
            O => \N__15243\,
            I => \N__15240\
        );

    \I__2807\ : LocalMux
    port map (
            O => \N__15240\,
            I => \ppm_encoder_1.un1_elevator_cry_9_THRU_CO\
        );

    \I__2806\ : InMux
    port map (
            O => \N__15237\,
            I => \N__15234\
        );

    \I__2805\ : LocalMux
    port map (
            O => \N__15234\,
            I => \N__15231\
        );

    \I__2804\ : Span4Mux_v
    port map (
            O => \N__15231\,
            I => \N__15226\
        );

    \I__2803\ : InMux
    port map (
            O => \N__15230\,
            I => \N__15223\
        );

    \I__2802\ : InMux
    port map (
            O => \N__15229\,
            I => \N__15219\
        );

    \I__2801\ : Span4Mux_v
    port map (
            O => \N__15226\,
            I => \N__15214\
        );

    \I__2800\ : LocalMux
    port map (
            O => \N__15223\,
            I => \N__15214\
        );

    \I__2799\ : CascadeMux
    port map (
            O => \N__15222\,
            I => \N__15211\
        );

    \I__2798\ : LocalMux
    port map (
            O => \N__15219\,
            I => \N__15208\
        );

    \I__2797\ : Span4Mux_h
    port map (
            O => \N__15214\,
            I => \N__15205\
        );

    \I__2796\ : InMux
    port map (
            O => \N__15211\,
            I => \N__15202\
        );

    \I__2795\ : Odrv4
    port map (
            O => \N__15208\,
            I => \frame_decoder_OFF2data_0\
        );

    \I__2794\ : Odrv4
    port map (
            O => \N__15205\,
            I => \frame_decoder_OFF2data_0\
        );

    \I__2793\ : LocalMux
    port map (
            O => \N__15202\,
            I => \frame_decoder_OFF2data_0\
        );

    \I__2792\ : InMux
    port map (
            O => \N__15195\,
            I => \N__15191\
        );

    \I__2791\ : InMux
    port map (
            O => \N__15194\,
            I => \N__15188\
        );

    \I__2790\ : LocalMux
    port map (
            O => \N__15191\,
            I => \N__15185\
        );

    \I__2789\ : LocalMux
    port map (
            O => \N__15188\,
            I => \N__15181\
        );

    \I__2788\ : Span4Mux_v
    port map (
            O => \N__15185\,
            I => \N__15178\
        );

    \I__2787\ : InMux
    port map (
            O => \N__15184\,
            I => \N__15175\
        );

    \I__2786\ : Span4Mux_h
    port map (
            O => \N__15181\,
            I => \N__15171\
        );

    \I__2785\ : Span4Mux_h
    port map (
            O => \N__15178\,
            I => \N__15168\
        );

    \I__2784\ : LocalMux
    port map (
            O => \N__15175\,
            I => \N__15165\
        );

    \I__2783\ : InMux
    port map (
            O => \N__15174\,
            I => \N__15162\
        );

    \I__2782\ : Odrv4
    port map (
            O => \N__15171\,
            I => \frame_decoder_CH2data_0\
        );

    \I__2781\ : Odrv4
    port map (
            O => \N__15168\,
            I => \frame_decoder_CH2data_0\
        );

    \I__2780\ : Odrv12
    port map (
            O => \N__15165\,
            I => \frame_decoder_CH2data_0\
        );

    \I__2779\ : LocalMux
    port map (
            O => \N__15162\,
            I => \frame_decoder_CH2data_0\
        );

    \I__2778\ : InMux
    port map (
            O => \N__15153\,
            I => \N__15149\
        );

    \I__2777\ : CascadeMux
    port map (
            O => \N__15152\,
            I => \N__15146\
        );

    \I__2776\ : LocalMux
    port map (
            O => \N__15149\,
            I => \N__15143\
        );

    \I__2775\ : InMux
    port map (
            O => \N__15146\,
            I => \N__15140\
        );

    \I__2774\ : Odrv12
    port map (
            O => \N__15143\,
            I => scaler_2_data_4
        );

    \I__2773\ : LocalMux
    port map (
            O => \N__15140\,
            I => scaler_2_data_4
        );

    \I__2772\ : InMux
    port map (
            O => \N__15135\,
            I => \N__15131\
        );

    \I__2771\ : InMux
    port map (
            O => \N__15134\,
            I => \N__15128\
        );

    \I__2770\ : LocalMux
    port map (
            O => \N__15131\,
            I => \N__15123\
        );

    \I__2769\ : LocalMux
    port map (
            O => \N__15128\,
            I => \N__15123\
        );

    \I__2768\ : Span4Mux_h
    port map (
            O => \N__15123\,
            I => \N__15120\
        );

    \I__2767\ : Odrv4
    port map (
            O => \N__15120\,
            I => scaler_4_data_12
        );

    \I__2766\ : InMux
    port map (
            O => \N__15117\,
            I => \N__15114\
        );

    \I__2765\ : LocalMux
    port map (
            O => \N__15114\,
            I => \N__15111\
        );

    \I__2764\ : Odrv4
    port map (
            O => \N__15111\,
            I => \ppm_encoder_1.un1_rudder_cry_11_THRU_CO\
        );

    \I__2763\ : InMux
    port map (
            O => \N__15108\,
            I => \N__15102\
        );

    \I__2762\ : InMux
    port map (
            O => \N__15107\,
            I => \N__15099\
        );

    \I__2761\ : InMux
    port map (
            O => \N__15106\,
            I => \N__15096\
        );

    \I__2760\ : InMux
    port map (
            O => \N__15105\,
            I => \N__15090\
        );

    \I__2759\ : LocalMux
    port map (
            O => \N__15102\,
            I => \N__15083\
        );

    \I__2758\ : LocalMux
    port map (
            O => \N__15099\,
            I => \N__15083\
        );

    \I__2757\ : LocalMux
    port map (
            O => \N__15096\,
            I => \N__15083\
        );

    \I__2756\ : InMux
    port map (
            O => \N__15095\,
            I => \N__15080\
        );

    \I__2755\ : InMux
    port map (
            O => \N__15094\,
            I => \N__15077\
        );

    \I__2754\ : InMux
    port map (
            O => \N__15093\,
            I => \N__15074\
        );

    \I__2753\ : LocalMux
    port map (
            O => \N__15090\,
            I => \N__15070\
        );

    \I__2752\ : Span4Mux_v
    port map (
            O => \N__15083\,
            I => \N__15061\
        );

    \I__2751\ : LocalMux
    port map (
            O => \N__15080\,
            I => \N__15061\
        );

    \I__2750\ : LocalMux
    port map (
            O => \N__15077\,
            I => \N__15061\
        );

    \I__2749\ : LocalMux
    port map (
            O => \N__15074\,
            I => \N__15061\
        );

    \I__2748\ : InMux
    port map (
            O => \N__15073\,
            I => \N__15058\
        );

    \I__2747\ : Span4Mux_v
    port map (
            O => \N__15070\,
            I => \N__15053\
        );

    \I__2746\ : Span4Mux_v
    port map (
            O => \N__15061\,
            I => \N__15048\
        );

    \I__2745\ : LocalMux
    port map (
            O => \N__15058\,
            I => \N__15048\
        );

    \I__2744\ : InMux
    port map (
            O => \N__15057\,
            I => \N__15045\
        );

    \I__2743\ : InMux
    port map (
            O => \N__15056\,
            I => \N__15042\
        );

    \I__2742\ : Odrv4
    port map (
            O => \N__15053\,
            I => uart_data_4
        );

    \I__2741\ : Odrv4
    port map (
            O => \N__15048\,
            I => uart_data_4
        );

    \I__2740\ : LocalMux
    port map (
            O => \N__15045\,
            I => uart_data_4
        );

    \I__2739\ : LocalMux
    port map (
            O => \N__15042\,
            I => uart_data_4
        );

    \I__2738\ : InMux
    port map (
            O => \N__15033\,
            I => \N__15030\
        );

    \I__2737\ : LocalMux
    port map (
            O => \N__15030\,
            I => \N__15027\
        );

    \I__2736\ : Odrv4
    port map (
            O => \N__15027\,
            I => \frame_decoder_CH1data_4\
        );

    \I__2735\ : CEMux
    port map (
            O => \N__15024\,
            I => \N__15021\
        );

    \I__2734\ : LocalMux
    port map (
            O => \N__15021\,
            I => \N__15018\
        );

    \I__2733\ : Span4Mux_v
    port map (
            O => \N__15018\,
            I => \N__15014\
        );

    \I__2732\ : CEMux
    port map (
            O => \N__15017\,
            I => \N__15011\
        );

    \I__2731\ : Span4Mux_h
    port map (
            O => \N__15014\,
            I => \N__15008\
        );

    \I__2730\ : LocalMux
    port map (
            O => \N__15011\,
            I => \N__15005\
        );

    \I__2729\ : Odrv4
    port map (
            O => \N__15008\,
            I => \uart_frame_decoder.source_CH1data_1_sqmuxa_0\
        );

    \I__2728\ : Odrv12
    port map (
            O => \N__15005\,
            I => \uart_frame_decoder.source_CH1data_1_sqmuxa_0\
        );

    \I__2727\ : InMux
    port map (
            O => \N__15000\,
            I => \N__14997\
        );

    \I__2726\ : LocalMux
    port map (
            O => \N__14997\,
            I => \ppm_encoder_1.un1_throttle_cry_11_THRU_CO\
        );

    \I__2725\ : InMux
    port map (
            O => \N__14994\,
            I => \N__14991\
        );

    \I__2724\ : LocalMux
    port map (
            O => \N__14991\,
            I => \N__14987\
        );

    \I__2723\ : InMux
    port map (
            O => \N__14990\,
            I => \N__14984\
        );

    \I__2722\ : Odrv12
    port map (
            O => \N__14987\,
            I => scaler_1_data_12
        );

    \I__2721\ : LocalMux
    port map (
            O => \N__14984\,
            I => scaler_1_data_12
        );

    \I__2720\ : InMux
    port map (
            O => \N__14979\,
            I => \N__14976\
        );

    \I__2719\ : LocalMux
    port map (
            O => \N__14976\,
            I => \N__14973\
        );

    \I__2718\ : Span4Mux_v
    port map (
            O => \N__14973\,
            I => \N__14969\
        );

    \I__2717\ : InMux
    port map (
            O => \N__14972\,
            I => \N__14966\
        );

    \I__2716\ : Odrv4
    port map (
            O => \N__14969\,
            I => scaler_1_data_13
        );

    \I__2715\ : LocalMux
    port map (
            O => \N__14966\,
            I => scaler_1_data_13
        );

    \I__2714\ : InMux
    port map (
            O => \N__14961\,
            I => \N__14958\
        );

    \I__2713\ : LocalMux
    port map (
            O => \N__14958\,
            I => \ppm_encoder_1.un1_throttle_cry_12_THRU_CO\
        );

    \I__2712\ : IoInMux
    port map (
            O => \N__14955\,
            I => \N__14952\
        );

    \I__2711\ : LocalMux
    port map (
            O => \N__14952\,
            I => \N__14949\
        );

    \I__2710\ : Span12Mux_s8_v
    port map (
            O => \N__14949\,
            I => \N__14943\
        );

    \I__2709\ : InMux
    port map (
            O => \N__14948\,
            I => \N__14940\
        );

    \I__2708\ : InMux
    port map (
            O => \N__14947\,
            I => \N__14934\
        );

    \I__2707\ : InMux
    port map (
            O => \N__14946\,
            I => \N__14934\
        );

    \I__2706\ : Span12Mux_h
    port map (
            O => \N__14943\,
            I => \N__14929\
        );

    \I__2705\ : LocalMux
    port map (
            O => \N__14940\,
            I => \N__14926\
        );

    \I__2704\ : InMux
    port map (
            O => \N__14939\,
            I => \N__14923\
        );

    \I__2703\ : LocalMux
    port map (
            O => \N__14934\,
            I => \N__14920\
        );

    \I__2702\ : InMux
    port map (
            O => \N__14933\,
            I => \N__14917\
        );

    \I__2701\ : CascadeMux
    port map (
            O => \N__14932\,
            I => \N__14913\
        );

    \I__2700\ : Span12Mux_v
    port map (
            O => \N__14929\,
            I => \N__14906\
        );

    \I__2699\ : Sp12to4
    port map (
            O => \N__14926\,
            I => \N__14906\
        );

    \I__2698\ : LocalMux
    port map (
            O => \N__14923\,
            I => \N__14906\
        );

    \I__2697\ : Span4Mux_h
    port map (
            O => \N__14920\,
            I => \N__14901\
        );

    \I__2696\ : LocalMux
    port map (
            O => \N__14917\,
            I => \N__14901\
        );

    \I__2695\ : InMux
    port map (
            O => \N__14916\,
            I => \N__14896\
        );

    \I__2694\ : InMux
    port map (
            O => \N__14913\,
            I => \N__14896\
        );

    \I__2693\ : Span12Mux_s9_v
    port map (
            O => \N__14906\,
            I => \N__14893\
        );

    \I__2692\ : Odrv4
    port map (
            O => \N__14901\,
            I => frame_decoder_dv_c
        );

    \I__2691\ : LocalMux
    port map (
            O => \N__14896\,
            I => frame_decoder_dv_c
        );

    \I__2690\ : Odrv12
    port map (
            O => \N__14893\,
            I => frame_decoder_dv_c
        );

    \I__2689\ : IoInMux
    port map (
            O => \N__14886\,
            I => \N__14883\
        );

    \I__2688\ : LocalMux
    port map (
            O => \N__14883\,
            I => frame_decoder_dv_c_0
        );

    \I__2687\ : InMux
    port map (
            O => \N__14880\,
            I => \N__14877\
        );

    \I__2686\ : LocalMux
    port map (
            O => \N__14877\,
            I => \ppm_encoder_1.N_415\
        );

    \I__2685\ : CascadeMux
    port map (
            O => \N__14874\,
            I => \ppm_encoder_1.N_414_cascade_\
        );

    \I__2684\ : CascadeMux
    port map (
            O => \N__14871\,
            I => \ppm_encoder_1.un2_throttle_iv_0_1_10_cascade_\
        );

    \I__2683\ : CascadeMux
    port map (
            O => \N__14868\,
            I => \ppm_encoder_1.un1_init_pulses_0_axb_10_cascade_\
        );

    \I__2682\ : CascadeMux
    port map (
            O => \N__14865\,
            I => \N__14861\
        );

    \I__2681\ : CascadeMux
    port map (
            O => \N__14864\,
            I => \N__14858\
        );

    \I__2680\ : InMux
    port map (
            O => \N__14861\,
            I => \N__14855\
        );

    \I__2679\ : InMux
    port map (
            O => \N__14858\,
            I => \N__14851\
        );

    \I__2678\ : LocalMux
    port map (
            O => \N__14855\,
            I => \N__14848\
        );

    \I__2677\ : InMux
    port map (
            O => \N__14854\,
            I => \N__14845\
        );

    \I__2676\ : LocalMux
    port map (
            O => \N__14851\,
            I => \ppm_encoder_1.elevatorZ0Z_9\
        );

    \I__2675\ : Odrv12
    port map (
            O => \N__14848\,
            I => \ppm_encoder_1.elevatorZ0Z_9\
        );

    \I__2674\ : LocalMux
    port map (
            O => \N__14845\,
            I => \ppm_encoder_1.elevatorZ0Z_9\
        );

    \I__2673\ : InMux
    port map (
            O => \N__14838\,
            I => \N__14835\
        );

    \I__2672\ : LocalMux
    port map (
            O => \N__14835\,
            I => \ppm_encoder_1.N_412\
        );

    \I__2671\ : CascadeMux
    port map (
            O => \N__14832\,
            I => \ppm_encoder_1.N_411_cascade_\
        );

    \I__2670\ : CascadeMux
    port map (
            O => \N__14829\,
            I => \ppm_encoder_1.un2_throttle_iv_0_1_9_cascade_\
        );

    \I__2669\ : InMux
    port map (
            O => \N__14826\,
            I => \N__14823\
        );

    \I__2668\ : LocalMux
    port map (
            O => \N__14823\,
            I => \ppm_encoder_1.un1_init_pulses_0_axb_9\
        );

    \I__2667\ : InMux
    port map (
            O => \N__14820\,
            I => \N__14817\
        );

    \I__2666\ : LocalMux
    port map (
            O => \N__14817\,
            I => \ppm_encoder_1.un1_aileron_cry_8_THRU_CO\
        );

    \I__2665\ : InMux
    port map (
            O => \N__14814\,
            I => \N__14811\
        );

    \I__2664\ : LocalMux
    port map (
            O => \N__14811\,
            I => \N__14807\
        );

    \I__2663\ : InMux
    port map (
            O => \N__14810\,
            I => \N__14804\
        );

    \I__2662\ : Span4Mux_v
    port map (
            O => \N__14807\,
            I => \N__14801\
        );

    \I__2661\ : LocalMux
    port map (
            O => \N__14804\,
            I => \N__14798\
        );

    \I__2660\ : Odrv4
    port map (
            O => \N__14801\,
            I => scaler_2_data_9
        );

    \I__2659\ : Odrv4
    port map (
            O => \N__14798\,
            I => scaler_2_data_9
        );

    \I__2658\ : InMux
    port map (
            O => \N__14793\,
            I => \N__14789\
        );

    \I__2657\ : InMux
    port map (
            O => \N__14792\,
            I => \N__14786\
        );

    \I__2656\ : LocalMux
    port map (
            O => \N__14789\,
            I => \ppm_encoder_1.elevatorZ0Z_4\
        );

    \I__2655\ : LocalMux
    port map (
            O => \N__14786\,
            I => \ppm_encoder_1.elevatorZ0Z_4\
        );

    \I__2654\ : InMux
    port map (
            O => \N__14781\,
            I => \N__14777\
        );

    \I__2653\ : InMux
    port map (
            O => \N__14780\,
            I => \N__14774\
        );

    \I__2652\ : LocalMux
    port map (
            O => \N__14777\,
            I => \ppm_encoder_1.aileronZ0Z_4\
        );

    \I__2651\ : LocalMux
    port map (
            O => \N__14774\,
            I => \ppm_encoder_1.aileronZ0Z_4\
        );

    \I__2650\ : InMux
    port map (
            O => \N__14769\,
            I => \N__14766\
        );

    \I__2649\ : LocalMux
    port map (
            O => \N__14766\,
            I => \N__14762\
        );

    \I__2648\ : InMux
    port map (
            O => \N__14765\,
            I => \N__14759\
        );

    \I__2647\ : Span4Mux_h
    port map (
            O => \N__14762\,
            I => \N__14754\
        );

    \I__2646\ : LocalMux
    port map (
            O => \N__14759\,
            I => \N__14754\
        );

    \I__2645\ : Span4Mux_v
    port map (
            O => \N__14754\,
            I => \N__14751\
        );

    \I__2644\ : Odrv4
    port map (
            O => \N__14751\,
            I => scaler_2_data_6
        );

    \I__2643\ : InMux
    port map (
            O => \N__14748\,
            I => \N__14742\
        );

    \I__2642\ : InMux
    port map (
            O => \N__14747\,
            I => \N__14742\
        );

    \I__2641\ : LocalMux
    port map (
            O => \N__14742\,
            I => \ppm_encoder_1.aileronZ0Z_6\
        );

    \I__2640\ : CascadeMux
    port map (
            O => \N__14739\,
            I => \N__14736\
        );

    \I__2639\ : InMux
    port map (
            O => \N__14736\,
            I => \N__14732\
        );

    \I__2638\ : InMux
    port map (
            O => \N__14735\,
            I => \N__14729\
        );

    \I__2637\ : LocalMux
    port map (
            O => \N__14732\,
            I => \N__14726\
        );

    \I__2636\ : LocalMux
    port map (
            O => \N__14729\,
            I => \ppm_encoder_1.elevatorZ0Z_6\
        );

    \I__2635\ : Odrv4
    port map (
            O => \N__14726\,
            I => \ppm_encoder_1.elevatorZ0Z_6\
        );

    \I__2634\ : CascadeMux
    port map (
            O => \N__14721\,
            I => \ppm_encoder_1.pulses2count_9_0_o2_0_6_cascade_\
        );

    \I__2633\ : InMux
    port map (
            O => \N__14718\,
            I => \N__14715\
        );

    \I__2632\ : LocalMux
    port map (
            O => \N__14715\,
            I => \ppm_encoder_1.un2_throttle_iv_0_rn_0_6\
        );

    \I__2631\ : CascadeMux
    port map (
            O => \N__14712\,
            I => \ppm_encoder_1.un2_throttle_0_6_cascade_\
        );

    \I__2630\ : CascadeMux
    port map (
            O => \N__14709\,
            I => \ppm_encoder_1.un1_init_pulses_0_axb_6_cascade_\
        );

    \I__2629\ : InMux
    port map (
            O => \N__14706\,
            I => \N__14703\
        );

    \I__2628\ : LocalMux
    port map (
            O => \N__14703\,
            I => \ppm_encoder_1.un2_throttle_iv_0_sn_6\
        );

    \I__2627\ : InMux
    port map (
            O => \N__14700\,
            I => \reset_module_System.count_1_cry_20\
        );

    \I__2626\ : InMux
    port map (
            O => \N__14697\,
            I => \N__14691\
        );

    \I__2625\ : InMux
    port map (
            O => \N__14696\,
            I => \N__14691\
        );

    \I__2624\ : LocalMux
    port map (
            O => \N__14691\,
            I => \reset_module_System.countZ0Z_19\
        );

    \I__2623\ : InMux
    port map (
            O => \N__14688\,
            I => \N__14684\
        );

    \I__2622\ : InMux
    port map (
            O => \N__14687\,
            I => \N__14681\
        );

    \I__2621\ : LocalMux
    port map (
            O => \N__14684\,
            I => \reset_module_System.countZ0Z_15\
        );

    \I__2620\ : LocalMux
    port map (
            O => \N__14681\,
            I => \reset_module_System.countZ0Z_15\
        );

    \I__2619\ : CascadeMux
    port map (
            O => \N__14676\,
            I => \N__14672\
        );

    \I__2618\ : InMux
    port map (
            O => \N__14675\,
            I => \N__14667\
        );

    \I__2617\ : InMux
    port map (
            O => \N__14672\,
            I => \N__14667\
        );

    \I__2616\ : LocalMux
    port map (
            O => \N__14667\,
            I => \reset_module_System.countZ0Z_21\
        );

    \I__2615\ : InMux
    port map (
            O => \N__14664\,
            I => \N__14660\
        );

    \I__2614\ : InMux
    port map (
            O => \N__14663\,
            I => \N__14657\
        );

    \I__2613\ : LocalMux
    port map (
            O => \N__14660\,
            I => \reset_module_System.countZ0Z_13\
        );

    \I__2612\ : LocalMux
    port map (
            O => \N__14657\,
            I => \reset_module_System.countZ0Z_13\
        );

    \I__2611\ : CascadeMux
    port map (
            O => \N__14652\,
            I => \N__14649\
        );

    \I__2610\ : InMux
    port map (
            O => \N__14649\,
            I => \N__14641\
        );

    \I__2609\ : InMux
    port map (
            O => \N__14648\,
            I => \N__14641\
        );

    \I__2608\ : InMux
    port map (
            O => \N__14647\,
            I => \N__14636\
        );

    \I__2607\ : InMux
    port map (
            O => \N__14646\,
            I => \N__14636\
        );

    \I__2606\ : LocalMux
    port map (
            O => \N__14641\,
            I => \N__14631\
        );

    \I__2605\ : LocalMux
    port map (
            O => \N__14636\,
            I => \N__14631\
        );

    \I__2604\ : Odrv4
    port map (
            O => \N__14631\,
            I => \reset_module_System.reset6_15\
        );

    \I__2603\ : InMux
    port map (
            O => \N__14628\,
            I => \N__14625\
        );

    \I__2602\ : LocalMux
    port map (
            O => \N__14625\,
            I => \N__14621\
        );

    \I__2601\ : CascadeMux
    port map (
            O => \N__14624\,
            I => \N__14618\
        );

    \I__2600\ : Span4Mux_v
    port map (
            O => \N__14621\,
            I => \N__14615\
        );

    \I__2599\ : InMux
    port map (
            O => \N__14618\,
            I => \N__14612\
        );

    \I__2598\ : Odrv4
    port map (
            O => \N__14615\,
            I => scaler_3_data_4
        );

    \I__2597\ : LocalMux
    port map (
            O => \N__14612\,
            I => scaler_3_data_4
        );

    \I__2596\ : InMux
    port map (
            O => \N__14607\,
            I => \N__14603\
        );

    \I__2595\ : CascadeMux
    port map (
            O => \N__14606\,
            I => \N__14599\
        );

    \I__2594\ : LocalMux
    port map (
            O => \N__14603\,
            I => \N__14595\
        );

    \I__2593\ : InMux
    port map (
            O => \N__14602\,
            I => \N__14592\
        );

    \I__2592\ : InMux
    port map (
            O => \N__14599\,
            I => \N__14587\
        );

    \I__2591\ : InMux
    port map (
            O => \N__14598\,
            I => \N__14587\
        );

    \I__2590\ : Odrv4
    port map (
            O => \N__14595\,
            I => \scaler_2.un2_source_data_0\
        );

    \I__2589\ : LocalMux
    port map (
            O => \N__14592\,
            I => \scaler_2.un2_source_data_0\
        );

    \I__2588\ : LocalMux
    port map (
            O => \N__14587\,
            I => \scaler_2.un2_source_data_0\
        );

    \I__2587\ : CascadeMux
    port map (
            O => \N__14580\,
            I => \N__14577\
        );

    \I__2586\ : InMux
    port map (
            O => \N__14577\,
            I => \N__14574\
        );

    \I__2585\ : LocalMux
    port map (
            O => \N__14574\,
            I => \N__14571\
        );

    \I__2584\ : Odrv4
    port map (
            O => \N__14571\,
            I => \scaler_2.un2_source_data_0_cry_1_c_RNO_0\
        );

    \I__2583\ : InMux
    port map (
            O => \N__14568\,
            I => \reset_module_System.count_1_cry_12\
        );

    \I__2582\ : InMux
    port map (
            O => \N__14565\,
            I => \N__14561\
        );

    \I__2581\ : InMux
    port map (
            O => \N__14564\,
            I => \N__14558\
        );

    \I__2580\ : LocalMux
    port map (
            O => \N__14561\,
            I => \reset_module_System.countZ0Z_14\
        );

    \I__2579\ : LocalMux
    port map (
            O => \N__14558\,
            I => \reset_module_System.countZ0Z_14\
        );

    \I__2578\ : InMux
    port map (
            O => \N__14553\,
            I => \reset_module_System.count_1_cry_13\
        );

    \I__2577\ : InMux
    port map (
            O => \N__14550\,
            I => \reset_module_System.count_1_cry_14\
        );

    \I__2576\ : InMux
    port map (
            O => \N__14547\,
            I => \N__14543\
        );

    \I__2575\ : InMux
    port map (
            O => \N__14546\,
            I => \N__14540\
        );

    \I__2574\ : LocalMux
    port map (
            O => \N__14543\,
            I => \reset_module_System.countZ0Z_16\
        );

    \I__2573\ : LocalMux
    port map (
            O => \N__14540\,
            I => \reset_module_System.countZ0Z_16\
        );

    \I__2572\ : InMux
    port map (
            O => \N__14535\,
            I => \reset_module_System.count_1_cry_15\
        );

    \I__2571\ : CascadeMux
    port map (
            O => \N__14532\,
            I => \N__14528\
        );

    \I__2570\ : InMux
    port map (
            O => \N__14531\,
            I => \N__14525\
        );

    \I__2569\ : InMux
    port map (
            O => \N__14528\,
            I => \N__14522\
        );

    \I__2568\ : LocalMux
    port map (
            O => \N__14525\,
            I => \reset_module_System.countZ0Z_17\
        );

    \I__2567\ : LocalMux
    port map (
            O => \N__14522\,
            I => \reset_module_System.countZ0Z_17\
        );

    \I__2566\ : InMux
    port map (
            O => \N__14517\,
            I => \bfn_5_19_0_\
        );

    \I__2565\ : CascadeMux
    port map (
            O => \N__14514\,
            I => \N__14511\
        );

    \I__2564\ : InMux
    port map (
            O => \N__14511\,
            I => \N__14507\
        );

    \I__2563\ : InMux
    port map (
            O => \N__14510\,
            I => \N__14504\
        );

    \I__2562\ : LocalMux
    port map (
            O => \N__14507\,
            I => \N__14501\
        );

    \I__2561\ : LocalMux
    port map (
            O => \N__14504\,
            I => \reset_module_System.countZ0Z_18\
        );

    \I__2560\ : Odrv4
    port map (
            O => \N__14501\,
            I => \reset_module_System.countZ0Z_18\
        );

    \I__2559\ : InMux
    port map (
            O => \N__14496\,
            I => \reset_module_System.count_1_cry_17\
        );

    \I__2558\ : InMux
    port map (
            O => \N__14493\,
            I => \reset_module_System.count_1_cry_18\
        );

    \I__2557\ : CascadeMux
    port map (
            O => \N__14490\,
            I => \N__14487\
        );

    \I__2556\ : InMux
    port map (
            O => \N__14487\,
            I => \N__14483\
        );

    \I__2555\ : InMux
    port map (
            O => \N__14486\,
            I => \N__14480\
        );

    \I__2554\ : LocalMux
    port map (
            O => \N__14483\,
            I => \N__14477\
        );

    \I__2553\ : LocalMux
    port map (
            O => \N__14480\,
            I => \reset_module_System.countZ0Z_20\
        );

    \I__2552\ : Odrv4
    port map (
            O => \N__14477\,
            I => \reset_module_System.countZ0Z_20\
        );

    \I__2551\ : InMux
    port map (
            O => \N__14472\,
            I => \reset_module_System.count_1_cry_19\
        );

    \I__2550\ : InMux
    port map (
            O => \N__14469\,
            I => \N__14465\
        );

    \I__2549\ : InMux
    port map (
            O => \N__14468\,
            I => \N__14462\
        );

    \I__2548\ : LocalMux
    port map (
            O => \N__14465\,
            I => \reset_module_System.countZ0Z_4\
        );

    \I__2547\ : LocalMux
    port map (
            O => \N__14462\,
            I => \reset_module_System.countZ0Z_4\
        );

    \I__2546\ : InMux
    port map (
            O => \N__14457\,
            I => \reset_module_System.count_1_cry_3\
        );

    \I__2545\ : InMux
    port map (
            O => \N__14454\,
            I => \N__14450\
        );

    \I__2544\ : InMux
    port map (
            O => \N__14453\,
            I => \N__14447\
        );

    \I__2543\ : LocalMux
    port map (
            O => \N__14450\,
            I => \reset_module_System.countZ0Z_5\
        );

    \I__2542\ : LocalMux
    port map (
            O => \N__14447\,
            I => \reset_module_System.countZ0Z_5\
        );

    \I__2541\ : InMux
    port map (
            O => \N__14442\,
            I => \reset_module_System.count_1_cry_4\
        );

    \I__2540\ : InMux
    port map (
            O => \N__14439\,
            I => \N__14435\
        );

    \I__2539\ : InMux
    port map (
            O => \N__14438\,
            I => \N__14432\
        );

    \I__2538\ : LocalMux
    port map (
            O => \N__14435\,
            I => \reset_module_System.countZ0Z_6\
        );

    \I__2537\ : LocalMux
    port map (
            O => \N__14432\,
            I => \reset_module_System.countZ0Z_6\
        );

    \I__2536\ : InMux
    port map (
            O => \N__14427\,
            I => \reset_module_System.count_1_cry_5\
        );

    \I__2535\ : InMux
    port map (
            O => \N__14424\,
            I => \N__14420\
        );

    \I__2534\ : InMux
    port map (
            O => \N__14423\,
            I => \N__14417\
        );

    \I__2533\ : LocalMux
    port map (
            O => \N__14420\,
            I => \reset_module_System.countZ0Z_7\
        );

    \I__2532\ : LocalMux
    port map (
            O => \N__14417\,
            I => \reset_module_System.countZ0Z_7\
        );

    \I__2531\ : InMux
    port map (
            O => \N__14412\,
            I => \reset_module_System.count_1_cry_6\
        );

    \I__2530\ : InMux
    port map (
            O => \N__14409\,
            I => \N__14405\
        );

    \I__2529\ : InMux
    port map (
            O => \N__14408\,
            I => \N__14402\
        );

    \I__2528\ : LocalMux
    port map (
            O => \N__14405\,
            I => \reset_module_System.countZ0Z_8\
        );

    \I__2527\ : LocalMux
    port map (
            O => \N__14402\,
            I => \reset_module_System.countZ0Z_8\
        );

    \I__2526\ : InMux
    port map (
            O => \N__14397\,
            I => \reset_module_System.count_1_cry_7\
        );

    \I__2525\ : CascadeMux
    port map (
            O => \N__14394\,
            I => \N__14390\
        );

    \I__2524\ : InMux
    port map (
            O => \N__14393\,
            I => \N__14387\
        );

    \I__2523\ : InMux
    port map (
            O => \N__14390\,
            I => \N__14384\
        );

    \I__2522\ : LocalMux
    port map (
            O => \N__14387\,
            I => \reset_module_System.countZ0Z_9\
        );

    \I__2521\ : LocalMux
    port map (
            O => \N__14384\,
            I => \reset_module_System.countZ0Z_9\
        );

    \I__2520\ : InMux
    port map (
            O => \N__14379\,
            I => \bfn_5_18_0_\
        );

    \I__2519\ : InMux
    port map (
            O => \N__14376\,
            I => \N__14372\
        );

    \I__2518\ : InMux
    port map (
            O => \N__14375\,
            I => \N__14369\
        );

    \I__2517\ : LocalMux
    port map (
            O => \N__14372\,
            I => \reset_module_System.countZ0Z_10\
        );

    \I__2516\ : LocalMux
    port map (
            O => \N__14369\,
            I => \reset_module_System.countZ0Z_10\
        );

    \I__2515\ : InMux
    port map (
            O => \N__14364\,
            I => \reset_module_System.count_1_cry_9\
        );

    \I__2514\ : InMux
    port map (
            O => \N__14361\,
            I => \N__14357\
        );

    \I__2513\ : InMux
    port map (
            O => \N__14360\,
            I => \N__14354\
        );

    \I__2512\ : LocalMux
    port map (
            O => \N__14357\,
            I => \reset_module_System.countZ0Z_11\
        );

    \I__2511\ : LocalMux
    port map (
            O => \N__14354\,
            I => \reset_module_System.countZ0Z_11\
        );

    \I__2510\ : InMux
    port map (
            O => \N__14349\,
            I => \reset_module_System.count_1_cry_10\
        );

    \I__2509\ : InMux
    port map (
            O => \N__14346\,
            I => \N__14342\
        );

    \I__2508\ : InMux
    port map (
            O => \N__14345\,
            I => \N__14339\
        );

    \I__2507\ : LocalMux
    port map (
            O => \N__14342\,
            I => \reset_module_System.countZ0Z_12\
        );

    \I__2506\ : LocalMux
    port map (
            O => \N__14339\,
            I => \reset_module_System.countZ0Z_12\
        );

    \I__2505\ : InMux
    port map (
            O => \N__14334\,
            I => \reset_module_System.count_1_cry_11\
        );

    \I__2504\ : InMux
    port map (
            O => \N__14331\,
            I => \uart.un4_timer_Count_1_cry_3\
        );

    \I__2503\ : CascadeMux
    port map (
            O => \N__14328\,
            I => \N__14321\
        );

    \I__2502\ : InMux
    port map (
            O => \N__14327\,
            I => \N__14318\
        );

    \I__2501\ : InMux
    port map (
            O => \N__14326\,
            I => \N__14311\
        );

    \I__2500\ : InMux
    port map (
            O => \N__14325\,
            I => \N__14311\
        );

    \I__2499\ : InMux
    port map (
            O => \N__14324\,
            I => \N__14311\
        );

    \I__2498\ : InMux
    port map (
            O => \N__14321\,
            I => \N__14308\
        );

    \I__2497\ : LocalMux
    port map (
            O => \N__14318\,
            I => \uart.timer_CountZ0Z_5\
        );

    \I__2496\ : LocalMux
    port map (
            O => \N__14311\,
            I => \uart.timer_CountZ0Z_5\
        );

    \I__2495\ : LocalMux
    port map (
            O => \N__14308\,
            I => \uart.timer_CountZ0Z_5\
        );

    \I__2494\ : InMux
    port map (
            O => \N__14301\,
            I => \uart.un4_timer_Count_1_cry_4\
        );

    \I__2493\ : InMux
    port map (
            O => \N__14298\,
            I => \N__14292\
        );

    \I__2492\ : InMux
    port map (
            O => \N__14297\,
            I => \N__14292\
        );

    \I__2491\ : LocalMux
    port map (
            O => \N__14292\,
            I => \N__14286\
        );

    \I__2490\ : CascadeMux
    port map (
            O => \N__14291\,
            I => \N__14283\
        );

    \I__2489\ : CascadeMux
    port map (
            O => \N__14290\,
            I => \N__14280\
        );

    \I__2488\ : InMux
    port map (
            O => \N__14289\,
            I => \N__14276\
        );

    \I__2487\ : Span4Mux_v
    port map (
            O => \N__14286\,
            I => \N__14273\
        );

    \I__2486\ : InMux
    port map (
            O => \N__14283\,
            I => \N__14268\
        );

    \I__2485\ : InMux
    port map (
            O => \N__14280\,
            I => \N__14268\
        );

    \I__2484\ : InMux
    port map (
            O => \N__14279\,
            I => \N__14265\
        );

    \I__2483\ : LocalMux
    port map (
            O => \N__14276\,
            I => \uart.timer_CountZ0Z_6\
        );

    \I__2482\ : Odrv4
    port map (
            O => \N__14273\,
            I => \uart.timer_CountZ0Z_6\
        );

    \I__2481\ : LocalMux
    port map (
            O => \N__14268\,
            I => \uart.timer_CountZ0Z_6\
        );

    \I__2480\ : LocalMux
    port map (
            O => \N__14265\,
            I => \uart.timer_CountZ0Z_6\
        );

    \I__2479\ : InMux
    port map (
            O => \N__14256\,
            I => \uart.un4_timer_Count_1_cry_5\
        );

    \I__2478\ : InMux
    port map (
            O => \N__14253\,
            I => \uart.un4_timer_Count_1_cry_6\
        );

    \I__2477\ : InMux
    port map (
            O => \N__14250\,
            I => \N__14244\
        );

    \I__2476\ : InMux
    port map (
            O => \N__14249\,
            I => \N__14241\
        );

    \I__2475\ : InMux
    port map (
            O => \N__14248\,
            I => \N__14237\
        );

    \I__2474\ : InMux
    port map (
            O => \N__14247\,
            I => \N__14234\
        );

    \I__2473\ : LocalMux
    port map (
            O => \N__14244\,
            I => \N__14228\
        );

    \I__2472\ : LocalMux
    port map (
            O => \N__14241\,
            I => \N__14228\
        );

    \I__2471\ : InMux
    port map (
            O => \N__14240\,
            I => \N__14224\
        );

    \I__2470\ : LocalMux
    port map (
            O => \N__14237\,
            I => \N__14219\
        );

    \I__2469\ : LocalMux
    port map (
            O => \N__14234\,
            I => \N__14219\
        );

    \I__2468\ : InMux
    port map (
            O => \N__14233\,
            I => \N__14214\
        );

    \I__2467\ : Span4Mux_v
    port map (
            O => \N__14228\,
            I => \N__14211\
        );

    \I__2466\ : InMux
    port map (
            O => \N__14227\,
            I => \N__14208\
        );

    \I__2465\ : LocalMux
    port map (
            O => \N__14224\,
            I => \N__14205\
        );

    \I__2464\ : Span4Mux_h
    port map (
            O => \N__14219\,
            I => \N__14202\
        );

    \I__2463\ : InMux
    port map (
            O => \N__14218\,
            I => \N__14197\
        );

    \I__2462\ : InMux
    port map (
            O => \N__14217\,
            I => \N__14197\
        );

    \I__2461\ : LocalMux
    port map (
            O => \N__14214\,
            I => \uart.timer_CountZ0Z_7\
        );

    \I__2460\ : Odrv4
    port map (
            O => \N__14211\,
            I => \uart.timer_CountZ0Z_7\
        );

    \I__2459\ : LocalMux
    port map (
            O => \N__14208\,
            I => \uart.timer_CountZ0Z_7\
        );

    \I__2458\ : Odrv4
    port map (
            O => \N__14205\,
            I => \uart.timer_CountZ0Z_7\
        );

    \I__2457\ : Odrv4
    port map (
            O => \N__14202\,
            I => \uart.timer_CountZ0Z_7\
        );

    \I__2456\ : LocalMux
    port map (
            O => \N__14197\,
            I => \uart.timer_CountZ0Z_7\
        );

    \I__2455\ : SRMux
    port map (
            O => \N__14184\,
            I => \N__14180\
        );

    \I__2454\ : SRMux
    port map (
            O => \N__14183\,
            I => \N__14177\
        );

    \I__2453\ : LocalMux
    port map (
            O => \N__14180\,
            I => \N__14173\
        );

    \I__2452\ : LocalMux
    port map (
            O => \N__14177\,
            I => \N__14170\
        );

    \I__2451\ : SRMux
    port map (
            O => \N__14176\,
            I => \N__14167\
        );

    \I__2450\ : Span4Mux_v
    port map (
            O => \N__14173\,
            I => \N__14164\
        );

    \I__2449\ : Span4Mux_v
    port map (
            O => \N__14170\,
            I => \N__14159\
        );

    \I__2448\ : LocalMux
    port map (
            O => \N__14167\,
            I => \N__14159\
        );

    \I__2447\ : Span4Mux_h
    port map (
            O => \N__14164\,
            I => \N__14156\
        );

    \I__2446\ : Span4Mux_h
    port map (
            O => \N__14159\,
            I => \N__14153\
        );

    \I__2445\ : Odrv4
    port map (
            O => \N__14156\,
            I => \uart.timer_Count_1_sqmuxa_i\
        );

    \I__2444\ : Odrv4
    port map (
            O => \N__14153\,
            I => \uart.timer_Count_1_sqmuxa_i\
        );

    \I__2443\ : CascadeMux
    port map (
            O => \N__14148\,
            I => \N__14145\
        );

    \I__2442\ : InMux
    port map (
            O => \N__14145\,
            I => \N__14139\
        );

    \I__2441\ : InMux
    port map (
            O => \N__14144\,
            I => \N__14136\
        );

    \I__2440\ : InMux
    port map (
            O => \N__14143\,
            I => \N__14133\
        );

    \I__2439\ : InMux
    port map (
            O => \N__14142\,
            I => \N__14130\
        );

    \I__2438\ : LocalMux
    port map (
            O => \N__14139\,
            I => \N__14125\
        );

    \I__2437\ : LocalMux
    port map (
            O => \N__14136\,
            I => \N__14125\
        );

    \I__2436\ : LocalMux
    port map (
            O => \N__14133\,
            I => \uart.timer_CountZ0Z_0\
        );

    \I__2435\ : LocalMux
    port map (
            O => \N__14130\,
            I => \uart.timer_CountZ0Z_0\
        );

    \I__2434\ : Odrv4
    port map (
            O => \N__14125\,
            I => \uart.timer_CountZ0Z_0\
        );

    \I__2433\ : InMux
    port map (
            O => \N__14118\,
            I => \N__14111\
        );

    \I__2432\ : InMux
    port map (
            O => \N__14117\,
            I => \N__14108\
        );

    \I__2431\ : InMux
    port map (
            O => \N__14116\,
            I => \N__14103\
        );

    \I__2430\ : InMux
    port map (
            O => \N__14115\,
            I => \N__14103\
        );

    \I__2429\ : InMux
    port map (
            O => \N__14114\,
            I => \N__14100\
        );

    \I__2428\ : LocalMux
    port map (
            O => \N__14111\,
            I => \uart.timer_CountZ0Z_4\
        );

    \I__2427\ : LocalMux
    port map (
            O => \N__14108\,
            I => \uart.timer_CountZ0Z_4\
        );

    \I__2426\ : LocalMux
    port map (
            O => \N__14103\,
            I => \uart.timer_CountZ0Z_4\
        );

    \I__2425\ : LocalMux
    port map (
            O => \N__14100\,
            I => \uart.timer_CountZ0Z_4\
        );

    \I__2424\ : InMux
    port map (
            O => \N__14091\,
            I => \N__14088\
        );

    \I__2423\ : LocalMux
    port map (
            O => \N__14088\,
            I => \uart.un1_state_2_0_a3_0\
        );

    \I__2422\ : InMux
    port map (
            O => \N__14085\,
            I => \N__14082\
        );

    \I__2421\ : LocalMux
    port map (
            O => \N__14082\,
            I => \N__14076\
        );

    \I__2420\ : InMux
    port map (
            O => \N__14081\,
            I => \N__14073\
        );

    \I__2419\ : InMux
    port map (
            O => \N__14080\,
            I => \N__14070\
        );

    \I__2418\ : InMux
    port map (
            O => \N__14079\,
            I => \N__14067\
        );

    \I__2417\ : Odrv4
    port map (
            O => \N__14076\,
            I => \reset_module_System.countZ0Z_0\
        );

    \I__2416\ : LocalMux
    port map (
            O => \N__14073\,
            I => \reset_module_System.countZ0Z_0\
        );

    \I__2415\ : LocalMux
    port map (
            O => \N__14070\,
            I => \reset_module_System.countZ0Z_0\
        );

    \I__2414\ : LocalMux
    port map (
            O => \N__14067\,
            I => \reset_module_System.countZ0Z_0\
        );

    \I__2413\ : InMux
    port map (
            O => \N__14058\,
            I => \N__14053\
        );

    \I__2412\ : CascadeMux
    port map (
            O => \N__14057\,
            I => \N__14050\
        );

    \I__2411\ : InMux
    port map (
            O => \N__14056\,
            I => \N__14047\
        );

    \I__2410\ : LocalMux
    port map (
            O => \N__14053\,
            I => \N__14044\
        );

    \I__2409\ : InMux
    port map (
            O => \N__14050\,
            I => \N__14041\
        );

    \I__2408\ : LocalMux
    port map (
            O => \N__14047\,
            I => \reset_module_System.countZ0Z_1\
        );

    \I__2407\ : Odrv12
    port map (
            O => \N__14044\,
            I => \reset_module_System.countZ0Z_1\
        );

    \I__2406\ : LocalMux
    port map (
            O => \N__14041\,
            I => \reset_module_System.countZ0Z_1\
        );

    \I__2405\ : InMux
    port map (
            O => \N__14034\,
            I => \N__14030\
        );

    \I__2404\ : InMux
    port map (
            O => \N__14033\,
            I => \N__14027\
        );

    \I__2403\ : LocalMux
    port map (
            O => \N__14030\,
            I => \reset_module_System.countZ0Z_2\
        );

    \I__2402\ : LocalMux
    port map (
            O => \N__14027\,
            I => \reset_module_System.countZ0Z_2\
        );

    \I__2401\ : InMux
    port map (
            O => \N__14022\,
            I => \N__14019\
        );

    \I__2400\ : LocalMux
    port map (
            O => \N__14019\,
            I => \reset_module_System.count_1_2\
        );

    \I__2399\ : InMux
    port map (
            O => \N__14016\,
            I => \reset_module_System.count_1_cry_1\
        );

    \I__2398\ : InMux
    port map (
            O => \N__14013\,
            I => \N__14009\
        );

    \I__2397\ : InMux
    port map (
            O => \N__14012\,
            I => \N__14006\
        );

    \I__2396\ : LocalMux
    port map (
            O => \N__14009\,
            I => \reset_module_System.countZ0Z_3\
        );

    \I__2395\ : LocalMux
    port map (
            O => \N__14006\,
            I => \reset_module_System.countZ0Z_3\
        );

    \I__2394\ : InMux
    port map (
            O => \N__14001\,
            I => \reset_module_System.count_1_cry_2\
        );

    \I__2393\ : InMux
    port map (
            O => \N__13998\,
            I => \ppm_encoder_1.un1_throttle_cry_10\
        );

    \I__2392\ : InMux
    port map (
            O => \N__13995\,
            I => \ppm_encoder_1.un1_throttle_cry_11\
        );

    \I__2391\ : InMux
    port map (
            O => \N__13992\,
            I => \ppm_encoder_1.un1_throttle_cry_12\
        );

    \I__2390\ : InMux
    port map (
            O => \N__13989\,
            I => \N__13986\
        );

    \I__2389\ : LocalMux
    port map (
            O => \N__13986\,
            I => scaler_1_data_14
        );

    \I__2388\ : InMux
    port map (
            O => \N__13983\,
            I => \bfn_4_30_0_\
        );

    \I__2387\ : InMux
    port map (
            O => \N__13980\,
            I => \N__13977\
        );

    \I__2386\ : LocalMux
    port map (
            O => \N__13977\,
            I => \uart_sync.aux_1__0_Z0Z_0\
        );

    \I__2385\ : InMux
    port map (
            O => \N__13974\,
            I => \N__13969\
        );

    \I__2384\ : InMux
    port map (
            O => \N__13973\,
            I => \N__13966\
        );

    \I__2383\ : InMux
    port map (
            O => \N__13972\,
            I => \N__13963\
        );

    \I__2382\ : LocalMux
    port map (
            O => \N__13969\,
            I => \N__13960\
        );

    \I__2381\ : LocalMux
    port map (
            O => \N__13966\,
            I => \N__13957\
        );

    \I__2380\ : LocalMux
    port map (
            O => \N__13963\,
            I => \uart.timer_CountZ0Z_1\
        );

    \I__2379\ : Odrv4
    port map (
            O => \N__13960\,
            I => \uart.timer_CountZ0Z_1\
        );

    \I__2378\ : Odrv4
    port map (
            O => \N__13957\,
            I => \uart.timer_CountZ0Z_1\
        );

    \I__2377\ : InMux
    port map (
            O => \N__13950\,
            I => \N__13944\
        );

    \I__2376\ : InMux
    port map (
            O => \N__13949\,
            I => \N__13941\
        );

    \I__2375\ : InMux
    port map (
            O => \N__13948\,
            I => \N__13936\
        );

    \I__2374\ : InMux
    port map (
            O => \N__13947\,
            I => \N__13936\
        );

    \I__2373\ : LocalMux
    port map (
            O => \N__13944\,
            I => \uart.timer_CountZ0Z_2\
        );

    \I__2372\ : LocalMux
    port map (
            O => \N__13941\,
            I => \uart.timer_CountZ0Z_2\
        );

    \I__2371\ : LocalMux
    port map (
            O => \N__13936\,
            I => \uart.timer_CountZ0Z_2\
        );

    \I__2370\ : InMux
    port map (
            O => \N__13929\,
            I => \uart.un4_timer_Count_1_cry_1\
        );

    \I__2369\ : CascadeMux
    port map (
            O => \N__13926\,
            I => \N__13921\
        );

    \I__2368\ : InMux
    port map (
            O => \N__13925\,
            I => \N__13917\
        );

    \I__2367\ : InMux
    port map (
            O => \N__13924\,
            I => \N__13914\
        );

    \I__2366\ : InMux
    port map (
            O => \N__13921\,
            I => \N__13909\
        );

    \I__2365\ : InMux
    port map (
            O => \N__13920\,
            I => \N__13909\
        );

    \I__2364\ : LocalMux
    port map (
            O => \N__13917\,
            I => \uart.timer_CountZ0Z_3\
        );

    \I__2363\ : LocalMux
    port map (
            O => \N__13914\,
            I => \uart.timer_CountZ0Z_3\
        );

    \I__2362\ : LocalMux
    port map (
            O => \N__13909\,
            I => \uart.timer_CountZ0Z_3\
        );

    \I__2361\ : InMux
    port map (
            O => \N__13902\,
            I => \uart.un4_timer_Count_1_cry_2\
        );

    \I__2360\ : InMux
    port map (
            O => \N__13899\,
            I => \N__13895\
        );

    \I__2359\ : InMux
    port map (
            O => \N__13898\,
            I => \N__13892\
        );

    \I__2358\ : LocalMux
    port map (
            O => \N__13895\,
            I => \N__13889\
        );

    \I__2357\ : LocalMux
    port map (
            O => \N__13892\,
            I => \N__13886\
        );

    \I__2356\ : Span4Mux_h
    port map (
            O => \N__13889\,
            I => \N__13883\
        );

    \I__2355\ : Span4Mux_h
    port map (
            O => \N__13886\,
            I => \N__13880\
        );

    \I__2354\ : Odrv4
    port map (
            O => \N__13883\,
            I => scaler_3_data_12
        );

    \I__2353\ : Odrv4
    port map (
            O => \N__13880\,
            I => scaler_3_data_12
        );

    \I__2352\ : InMux
    port map (
            O => \N__13875\,
            I => \N__13872\
        );

    \I__2351\ : LocalMux
    port map (
            O => \N__13872\,
            I => \ppm_encoder_1.un1_elevator_cry_11_THRU_CO\
        );

    \I__2350\ : InMux
    port map (
            O => \N__13869\,
            I => \ppm_encoder_1.un1_elevator_cry_11\
        );

    \I__2349\ : InMux
    port map (
            O => \N__13866\,
            I => \ppm_encoder_1.un1_elevator_cry_12\
        );

    \I__2348\ : InMux
    port map (
            O => \N__13863\,
            I => \N__13860\
        );

    \I__2347\ : LocalMux
    port map (
            O => \N__13860\,
            I => \N__13857\
        );

    \I__2346\ : Span4Mux_v
    port map (
            O => \N__13857\,
            I => \N__13854\
        );

    \I__2345\ : Odrv4
    port map (
            O => \N__13854\,
            I => scaler_3_data_14
        );

    \I__2344\ : InMux
    port map (
            O => \N__13851\,
            I => \bfn_4_28_0_\
        );

    \I__2343\ : InMux
    port map (
            O => \N__13848\,
            I => \N__13845\
        );

    \I__2342\ : LocalMux
    port map (
            O => \N__13845\,
            I => \N__13842\
        );

    \I__2341\ : Span4Mux_v
    port map (
            O => \N__13842\,
            I => \N__13838\
        );

    \I__2340\ : InMux
    port map (
            O => \N__13841\,
            I => \N__13835\
        );

    \I__2339\ : Odrv4
    port map (
            O => \N__13838\,
            I => scaler_1_data_6
        );

    \I__2338\ : LocalMux
    port map (
            O => \N__13835\,
            I => scaler_1_data_6
        );

    \I__2337\ : InMux
    port map (
            O => \N__13830\,
            I => \ppm_encoder_1.un1_throttle_cry_6\
        );

    \I__2336\ : InMux
    port map (
            O => \N__13827\,
            I => \ppm_encoder_1.un1_throttle_cry_7\
        );

    \I__2335\ : InMux
    port map (
            O => \N__13824\,
            I => \N__13821\
        );

    \I__2334\ : LocalMux
    port map (
            O => \N__13821\,
            I => \N__13817\
        );

    \I__2333\ : InMux
    port map (
            O => \N__13820\,
            I => \N__13814\
        );

    \I__2332\ : Odrv4
    port map (
            O => \N__13817\,
            I => scaler_1_data_9
        );

    \I__2331\ : LocalMux
    port map (
            O => \N__13814\,
            I => scaler_1_data_9
        );

    \I__2330\ : InMux
    port map (
            O => \N__13809\,
            I => \N__13806\
        );

    \I__2329\ : LocalMux
    port map (
            O => \N__13806\,
            I => \N__13803\
        );

    \I__2328\ : Odrv4
    port map (
            O => \N__13803\,
            I => \ppm_encoder_1.un1_throttle_cry_8_THRU_CO\
        );

    \I__2327\ : InMux
    port map (
            O => \N__13800\,
            I => \ppm_encoder_1.un1_throttle_cry_8\
        );

    \I__2326\ : InMux
    port map (
            O => \N__13797\,
            I => \N__13794\
        );

    \I__2325\ : LocalMux
    port map (
            O => \N__13794\,
            I => \N__13790\
        );

    \I__2324\ : InMux
    port map (
            O => \N__13793\,
            I => \N__13787\
        );

    \I__2323\ : Odrv4
    port map (
            O => \N__13790\,
            I => scaler_1_data_10
        );

    \I__2322\ : LocalMux
    port map (
            O => \N__13787\,
            I => scaler_1_data_10
        );

    \I__2321\ : InMux
    port map (
            O => \N__13782\,
            I => \N__13779\
        );

    \I__2320\ : LocalMux
    port map (
            O => \N__13779\,
            I => \N__13776\
        );

    \I__2319\ : Odrv4
    port map (
            O => \N__13776\,
            I => \ppm_encoder_1.un1_throttle_cry_9_THRU_CO\
        );

    \I__2318\ : InMux
    port map (
            O => \N__13773\,
            I => \ppm_encoder_1.un1_throttle_cry_9\
        );

    \I__2317\ : InMux
    port map (
            O => \N__13770\,
            I => \N__13766\
        );

    \I__2316\ : InMux
    port map (
            O => \N__13769\,
            I => \N__13763\
        );

    \I__2315\ : LocalMux
    port map (
            O => \N__13766\,
            I => \N__13760\
        );

    \I__2314\ : LocalMux
    port map (
            O => \N__13763\,
            I => \N__13757\
        );

    \I__2313\ : Span4Mux_h
    port map (
            O => \N__13760\,
            I => \N__13752\
        );

    \I__2312\ : Span4Mux_h
    port map (
            O => \N__13757\,
            I => \N__13752\
        );

    \I__2311\ : Odrv4
    port map (
            O => \N__13752\,
            I => scaler_3_data_6
        );

    \I__2310\ : InMux
    port map (
            O => \N__13749\,
            I => \N__13745\
        );

    \I__2309\ : InMux
    port map (
            O => \N__13748\,
            I => \N__13742\
        );

    \I__2308\ : LocalMux
    port map (
            O => \N__13745\,
            I => \N__13739\
        );

    \I__2307\ : LocalMux
    port map (
            O => \N__13742\,
            I => \N__13736\
        );

    \I__2306\ : Span4Mux_v
    port map (
            O => \N__13739\,
            I => \N__13731\
        );

    \I__2305\ : Span4Mux_v
    port map (
            O => \N__13736\,
            I => \N__13731\
        );

    \I__2304\ : Odrv4
    port map (
            O => \N__13731\,
            I => scaler_3_data_7
        );

    \I__2303\ : InMux
    port map (
            O => \N__13728\,
            I => \N__13725\
        );

    \I__2302\ : LocalMux
    port map (
            O => \N__13725\,
            I => \N__13722\
        );

    \I__2301\ : Odrv12
    port map (
            O => \N__13722\,
            I => \ppm_encoder_1.un1_elevator_cry_6_THRU_CO\
        );

    \I__2300\ : InMux
    port map (
            O => \N__13719\,
            I => \ppm_encoder_1.un1_elevator_cry_6\
        );

    \I__2299\ : InMux
    port map (
            O => \N__13716\,
            I => \ppm_encoder_1.un1_elevator_cry_7\
        );

    \I__2298\ : InMux
    port map (
            O => \N__13713\,
            I => \N__13710\
        );

    \I__2297\ : LocalMux
    port map (
            O => \N__13710\,
            I => \N__13706\
        );

    \I__2296\ : InMux
    port map (
            O => \N__13709\,
            I => \N__13703\
        );

    \I__2295\ : Span4Mux_v
    port map (
            O => \N__13706\,
            I => \N__13698\
        );

    \I__2294\ : LocalMux
    port map (
            O => \N__13703\,
            I => \N__13698\
        );

    \I__2293\ : Span4Mux_h
    port map (
            O => \N__13698\,
            I => \N__13695\
        );

    \I__2292\ : Odrv4
    port map (
            O => \N__13695\,
            I => scaler_3_data_9
        );

    \I__2291\ : InMux
    port map (
            O => \N__13692\,
            I => \N__13689\
        );

    \I__2290\ : LocalMux
    port map (
            O => \N__13689\,
            I => \ppm_encoder_1.un1_elevator_cry_8_THRU_CO\
        );

    \I__2289\ : InMux
    port map (
            O => \N__13686\,
            I => \ppm_encoder_1.un1_elevator_cry_8\
        );

    \I__2288\ : InMux
    port map (
            O => \N__13683\,
            I => \ppm_encoder_1.un1_elevator_cry_9\
        );

    \I__2287\ : InMux
    port map (
            O => \N__13680\,
            I => \ppm_encoder_1.un1_elevator_cry_10\
        );

    \I__2286\ : InMux
    port map (
            O => \N__13677\,
            I => \ppm_encoder_1.un1_aileron_cry_9\
        );

    \I__2285\ : InMux
    port map (
            O => \N__13674\,
            I => \N__13670\
        );

    \I__2284\ : InMux
    port map (
            O => \N__13673\,
            I => \N__13667\
        );

    \I__2283\ : LocalMux
    port map (
            O => \N__13670\,
            I => \N__13662\
        );

    \I__2282\ : LocalMux
    port map (
            O => \N__13667\,
            I => \N__13662\
        );

    \I__2281\ : Span4Mux_v
    port map (
            O => \N__13662\,
            I => \N__13659\
        );

    \I__2280\ : Odrv4
    port map (
            O => \N__13659\,
            I => scaler_2_data_11
        );

    \I__2279\ : InMux
    port map (
            O => \N__13656\,
            I => \N__13653\
        );

    \I__2278\ : LocalMux
    port map (
            O => \N__13653\,
            I => \ppm_encoder_1.un1_aileron_cry_10_THRU_CO\
        );

    \I__2277\ : InMux
    port map (
            O => \N__13650\,
            I => \ppm_encoder_1.un1_aileron_cry_10\
        );

    \I__2276\ : InMux
    port map (
            O => \N__13647\,
            I => \ppm_encoder_1.un1_aileron_cry_11\
        );

    \I__2275\ : InMux
    port map (
            O => \N__13644\,
            I => \ppm_encoder_1.un1_aileron_cry_12\
        );

    \I__2274\ : InMux
    port map (
            O => \N__13641\,
            I => \N__13638\
        );

    \I__2273\ : LocalMux
    port map (
            O => \N__13638\,
            I => \N__13635\
        );

    \I__2272\ : Span4Mux_v
    port map (
            O => \N__13635\,
            I => \N__13632\
        );

    \I__2271\ : Odrv4
    port map (
            O => \N__13632\,
            I => scaler_2_data_14
        );

    \I__2270\ : InMux
    port map (
            O => \N__13629\,
            I => \bfn_4_25_0_\
        );

    \I__2269\ : InMux
    port map (
            O => \N__13626\,
            I => \N__13623\
        );

    \I__2268\ : LocalMux
    port map (
            O => \N__13623\,
            I => \ppm_encoder_1.un1_rudder_cry_9_THRU_CO\
        );

    \I__2267\ : InMux
    port map (
            O => \N__13620\,
            I => \N__13617\
        );

    \I__2266\ : LocalMux
    port map (
            O => \N__13617\,
            I => \N__13613\
        );

    \I__2265\ : CascadeMux
    port map (
            O => \N__13616\,
            I => \N__13610\
        );

    \I__2264\ : Span4Mux_v
    port map (
            O => \N__13613\,
            I => \N__13607\
        );

    \I__2263\ : InMux
    port map (
            O => \N__13610\,
            I => \N__13604\
        );

    \I__2262\ : Span4Mux_s1_v
    port map (
            O => \N__13607\,
            I => \N__13601\
        );

    \I__2261\ : LocalMux
    port map (
            O => \N__13604\,
            I => \N__13598\
        );

    \I__2260\ : Odrv4
    port map (
            O => \N__13601\,
            I => scaler_4_data_10
        );

    \I__2259\ : Odrv4
    port map (
            O => \N__13598\,
            I => scaler_4_data_10
        );

    \I__2258\ : InMux
    port map (
            O => \N__13593\,
            I => \N__13590\
        );

    \I__2257\ : LocalMux
    port map (
            O => \N__13590\,
            I => \N__13586\
        );

    \I__2256\ : InMux
    port map (
            O => \N__13589\,
            I => \N__13583\
        );

    \I__2255\ : Span4Mux_v
    port map (
            O => \N__13586\,
            I => \N__13580\
        );

    \I__2254\ : LocalMux
    port map (
            O => \N__13583\,
            I => \N__13577\
        );

    \I__2253\ : Odrv4
    port map (
            O => \N__13580\,
            I => scaler_2_data_10
        );

    \I__2252\ : Odrv4
    port map (
            O => \N__13577\,
            I => scaler_2_data_10
        );

    \I__2251\ : InMux
    port map (
            O => \N__13572\,
            I => \N__13569\
        );

    \I__2250\ : LocalMux
    port map (
            O => \N__13569\,
            I => \N__13566\
        );

    \I__2249\ : Odrv4
    port map (
            O => \N__13566\,
            I => \ppm_encoder_1.un1_aileron_cry_9_THRU_CO\
        );

    \I__2248\ : InMux
    port map (
            O => \N__13563\,
            I => \N__13560\
        );

    \I__2247\ : LocalMux
    port map (
            O => \N__13560\,
            I => \N__13556\
        );

    \I__2246\ : InMux
    port map (
            O => \N__13559\,
            I => \N__13553\
        );

    \I__2245\ : Span4Mux_h
    port map (
            O => \N__13556\,
            I => \N__13550\
        );

    \I__2244\ : LocalMux
    port map (
            O => \N__13553\,
            I => \N__13547\
        );

    \I__2243\ : Span4Mux_s2_h
    port map (
            O => \N__13550\,
            I => \N__13542\
        );

    \I__2242\ : Span4Mux_h
    port map (
            O => \N__13547\,
            I => \N__13542\
        );

    \I__2241\ : Odrv4
    port map (
            O => \N__13542\,
            I => scaler_4_data_13
        );

    \I__2240\ : InMux
    port map (
            O => \N__13539\,
            I => \N__13536\
        );

    \I__2239\ : LocalMux
    port map (
            O => \N__13536\,
            I => \ppm_encoder_1.un1_rudder_cry_12_THRU_CO\
        );

    \I__2238\ : InMux
    port map (
            O => \N__13533\,
            I => \N__13530\
        );

    \I__2237\ : LocalMux
    port map (
            O => \N__13530\,
            I => \N__13527\
        );

    \I__2236\ : Span4Mux_h
    port map (
            O => \N__13527\,
            I => \N__13523\
        );

    \I__2235\ : InMux
    port map (
            O => \N__13526\,
            I => \N__13520\
        );

    \I__2234\ : Span4Mux_v
    port map (
            O => \N__13523\,
            I => \N__13517\
        );

    \I__2233\ : LocalMux
    port map (
            O => \N__13520\,
            I => \N__13514\
        );

    \I__2232\ : Odrv4
    port map (
            O => \N__13517\,
            I => scaler_4_data_6
        );

    \I__2231\ : Odrv4
    port map (
            O => \N__13514\,
            I => scaler_4_data_6
        );

    \I__2230\ : InMux
    port map (
            O => \N__13509\,
            I => \N__13506\
        );

    \I__2229\ : LocalMux
    port map (
            O => \N__13506\,
            I => \N__13500\
        );

    \I__2228\ : InMux
    port map (
            O => \N__13505\,
            I => \N__13497\
        );

    \I__2227\ : InMux
    port map (
            O => \N__13504\,
            I => \N__13494\
        );

    \I__2226\ : CascadeMux
    port map (
            O => \N__13503\,
            I => \N__13491\
        );

    \I__2225\ : Span4Mux_v
    port map (
            O => \N__13500\,
            I => \N__13486\
        );

    \I__2224\ : LocalMux
    port map (
            O => \N__13497\,
            I => \N__13486\
        );

    \I__2223\ : LocalMux
    port map (
            O => \N__13494\,
            I => \N__13483\
        );

    \I__2222\ : InMux
    port map (
            O => \N__13491\,
            I => \N__13480\
        );

    \I__2221\ : Odrv4
    port map (
            O => \N__13486\,
            I => \frame_decoder_OFF3data_0\
        );

    \I__2220\ : Odrv4
    port map (
            O => \N__13483\,
            I => \frame_decoder_OFF3data_0\
        );

    \I__2219\ : LocalMux
    port map (
            O => \N__13480\,
            I => \frame_decoder_OFF3data_0\
        );

    \I__2218\ : InMux
    port map (
            O => \N__13473\,
            I => \N__13469\
        );

    \I__2217\ : InMux
    port map (
            O => \N__13472\,
            I => \N__13466\
        );

    \I__2216\ : LocalMux
    port map (
            O => \N__13469\,
            I => \N__13461\
        );

    \I__2215\ : LocalMux
    port map (
            O => \N__13466\,
            I => \N__13461\
        );

    \I__2214\ : Span4Mux_v
    port map (
            O => \N__13461\,
            I => \N__13456\
        );

    \I__2213\ : InMux
    port map (
            O => \N__13460\,
            I => \N__13453\
        );

    \I__2212\ : InMux
    port map (
            O => \N__13459\,
            I => \N__13450\
        );

    \I__2211\ : Odrv4
    port map (
            O => \N__13456\,
            I => \frame_decoder_CH3data_0\
        );

    \I__2210\ : LocalMux
    port map (
            O => \N__13453\,
            I => \frame_decoder_CH3data_0\
        );

    \I__2209\ : LocalMux
    port map (
            O => \N__13450\,
            I => \frame_decoder_CH3data_0\
        );

    \I__2208\ : InMux
    port map (
            O => \N__13443\,
            I => \ppm_encoder_1.un1_aileron_cry_6\
        );

    \I__2207\ : InMux
    port map (
            O => \N__13440\,
            I => \ppm_encoder_1.un1_aileron_cry_7\
        );

    \I__2206\ : InMux
    port map (
            O => \N__13437\,
            I => \ppm_encoder_1.un1_aileron_cry_8\
        );

    \I__2205\ : InMux
    port map (
            O => \N__13434\,
            I => \N__13431\
        );

    \I__2204\ : LocalMux
    port map (
            O => \N__13431\,
            I => \N__13427\
        );

    \I__2203\ : InMux
    port map (
            O => \N__13430\,
            I => \N__13424\
        );

    \I__2202\ : Span4Mux_h
    port map (
            O => \N__13427\,
            I => \N__13421\
        );

    \I__2201\ : LocalMux
    port map (
            O => \N__13424\,
            I => \uart_frame_decoder.state_1Z0Z_6\
        );

    \I__2200\ : Odrv4
    port map (
            O => \N__13421\,
            I => \uart_frame_decoder.state_1Z0Z_6\
        );

    \I__2199\ : InMux
    port map (
            O => \N__13416\,
            I => \N__13413\
        );

    \I__2198\ : LocalMux
    port map (
            O => \N__13413\,
            I => \N__13410\
        );

    \I__2197\ : Span4Mux_h
    port map (
            O => \N__13410\,
            I => \N__13407\
        );

    \I__2196\ : Odrv4
    port map (
            O => \N__13407\,
            I => \uart_frame_decoder.source_offset1data_1_sqmuxa\
        );

    \I__2195\ : CascadeMux
    port map (
            O => \N__13404\,
            I => \uart_frame_decoder.source_offset1data_1_sqmuxa_cascade_\
        );

    \I__2194\ : CEMux
    port map (
            O => \N__13401\,
            I => \N__13398\
        );

    \I__2193\ : LocalMux
    port map (
            O => \N__13398\,
            I => \N__13395\
        );

    \I__2192\ : Span4Mux_h
    port map (
            O => \N__13395\,
            I => \N__13392\
        );

    \I__2191\ : Span4Mux_v
    port map (
            O => \N__13392\,
            I => \N__13389\
        );

    \I__2190\ : Odrv4
    port map (
            O => \N__13389\,
            I => \uart_frame_decoder.source_offset1data_1_sqmuxa_0\
        );

    \I__2189\ : InMux
    port map (
            O => \N__13386\,
            I => \N__13368\
        );

    \I__2188\ : InMux
    port map (
            O => \N__13385\,
            I => \N__13368\
        );

    \I__2187\ : InMux
    port map (
            O => \N__13384\,
            I => \N__13368\
        );

    \I__2186\ : InMux
    port map (
            O => \N__13383\,
            I => \N__13368\
        );

    \I__2185\ : InMux
    port map (
            O => \N__13382\,
            I => \N__13368\
        );

    \I__2184\ : InMux
    port map (
            O => \N__13381\,
            I => \N__13361\
        );

    \I__2183\ : InMux
    port map (
            O => \N__13380\,
            I => \N__13361\
        );

    \I__2182\ : InMux
    port map (
            O => \N__13379\,
            I => \N__13361\
        );

    \I__2181\ : LocalMux
    port map (
            O => \N__13368\,
            I => \N__13355\
        );

    \I__2180\ : LocalMux
    port map (
            O => \N__13361\,
            I => \N__13355\
        );

    \I__2179\ : InMux
    port map (
            O => \N__13360\,
            I => \N__13352\
        );

    \I__2178\ : Odrv4
    port map (
            O => \N__13355\,
            I => \uart.data_rdyc_1\
        );

    \I__2177\ : LocalMux
    port map (
            O => \N__13352\,
            I => \uart.data_rdyc_1\
        );

    \I__2176\ : InMux
    port map (
            O => \N__13347\,
            I => \N__13343\
        );

    \I__2175\ : CascadeMux
    port map (
            O => \N__13346\,
            I => \N__13340\
        );

    \I__2174\ : LocalMux
    port map (
            O => \N__13343\,
            I => \N__13337\
        );

    \I__2173\ : InMux
    port map (
            O => \N__13340\,
            I => \N__13334\
        );

    \I__2172\ : Odrv4
    port map (
            O => \N__13337\,
            I => \uart.data_AuxZ0Z_4\
        );

    \I__2171\ : LocalMux
    port map (
            O => \N__13334\,
            I => \uart.data_AuxZ0Z_4\
        );

    \I__2170\ : SRMux
    port map (
            O => \N__13329\,
            I => \N__13326\
        );

    \I__2169\ : LocalMux
    port map (
            O => \N__13326\,
            I => \N__13322\
        );

    \I__2168\ : SRMux
    port map (
            O => \N__13325\,
            I => \N__13319\
        );

    \I__2167\ : Span4Mux_h
    port map (
            O => \N__13322\,
            I => \N__13316\
        );

    \I__2166\ : LocalMux
    port map (
            O => \N__13319\,
            I => \N__13313\
        );

    \I__2165\ : Odrv4
    port map (
            O => \N__13316\,
            I => \uart.state_RNIQABT2Z0Z_4\
        );

    \I__2164\ : Odrv12
    port map (
            O => \N__13313\,
            I => \uart.state_RNIQABT2Z0Z_4\
        );

    \I__2163\ : InMux
    port map (
            O => \N__13308\,
            I => \N__13305\
        );

    \I__2162\ : LocalMux
    port map (
            O => \N__13305\,
            I => \N__13302\
        );

    \I__2161\ : Span4Mux_h
    port map (
            O => \N__13302\,
            I => \N__13298\
        );

    \I__2160\ : InMux
    port map (
            O => \N__13301\,
            I => \N__13295\
        );

    \I__2159\ : Odrv4
    port map (
            O => \N__13298\,
            I => \uart_frame_decoder.state_1_ns_0_i_o2_0_10\
        );

    \I__2158\ : LocalMux
    port map (
            O => \N__13295\,
            I => \uart_frame_decoder.state_1_ns_0_i_o2_0_10\
        );

    \I__2157\ : CascadeMux
    port map (
            O => \N__13290\,
            I => \N__13286\
        );

    \I__2156\ : InMux
    port map (
            O => \N__13289\,
            I => \N__13283\
        );

    \I__2155\ : InMux
    port map (
            O => \N__13286\,
            I => \N__13280\
        );

    \I__2154\ : LocalMux
    port map (
            O => \N__13283\,
            I => \N__13277\
        );

    \I__2153\ : LocalMux
    port map (
            O => \N__13280\,
            I => \N__13274\
        );

    \I__2152\ : Span4Mux_v
    port map (
            O => \N__13277\,
            I => \N__13271\
        );

    \I__2151\ : Odrv4
    port map (
            O => \N__13274\,
            I => \uart_frame_decoder.source_offset4data_1_sqmuxa\
        );

    \I__2150\ : Odrv4
    port map (
            O => \N__13271\,
            I => \uart_frame_decoder.source_offset4data_1_sqmuxa\
        );

    \I__2149\ : InMux
    port map (
            O => \N__13266\,
            I => \N__13254\
        );

    \I__2148\ : InMux
    port map (
            O => \N__13265\,
            I => \N__13254\
        );

    \I__2147\ : InMux
    port map (
            O => \N__13264\,
            I => \N__13254\
        );

    \I__2146\ : InMux
    port map (
            O => \N__13263\,
            I => \N__13254\
        );

    \I__2145\ : LocalMux
    port map (
            O => \N__13254\,
            I => \N__13250\
        );

    \I__2144\ : InMux
    port map (
            O => \N__13253\,
            I => \N__13247\
        );

    \I__2143\ : Span4Mux_v
    port map (
            O => \N__13250\,
            I => \N__13241\
        );

    \I__2142\ : LocalMux
    port map (
            O => \N__13247\,
            I => \N__13241\
        );

    \I__2141\ : InMux
    port map (
            O => \N__13246\,
            I => \N__13238\
        );

    \I__2140\ : Span4Mux_v
    port map (
            O => \N__13241\,
            I => \N__13231\
        );

    \I__2139\ : LocalMux
    port map (
            O => \N__13238\,
            I => \N__13228\
        );

    \I__2138\ : InMux
    port map (
            O => \N__13237\,
            I => \N__13225\
        );

    \I__2137\ : InMux
    port map (
            O => \N__13236\,
            I => \N__13218\
        );

    \I__2136\ : InMux
    port map (
            O => \N__13235\,
            I => \N__13218\
        );

    \I__2135\ : InMux
    port map (
            O => \N__13234\,
            I => \N__13218\
        );

    \I__2134\ : Odrv4
    port map (
            O => \N__13231\,
            I => \uart_frame_decoder.WDT_RNIJUEI2Z0Z_15\
        );

    \I__2133\ : Odrv4
    port map (
            O => \N__13228\,
            I => \uart_frame_decoder.WDT_RNIJUEI2Z0Z_15\
        );

    \I__2132\ : LocalMux
    port map (
            O => \N__13225\,
            I => \uart_frame_decoder.WDT_RNIJUEI2Z0Z_15\
        );

    \I__2131\ : LocalMux
    port map (
            O => \N__13218\,
            I => \uart_frame_decoder.WDT_RNIJUEI2Z0Z_15\
        );

    \I__2130\ : InMux
    port map (
            O => \N__13209\,
            I => \N__13205\
        );

    \I__2129\ : InMux
    port map (
            O => \N__13208\,
            I => \N__13202\
        );

    \I__2128\ : LocalMux
    port map (
            O => \N__13205\,
            I => \N__13199\
        );

    \I__2127\ : LocalMux
    port map (
            O => \N__13202\,
            I => \N__13196\
        );

    \I__2126\ : Span12Mux_v
    port map (
            O => \N__13199\,
            I => \N__13193\
        );

    \I__2125\ : Span4Mux_h
    port map (
            O => \N__13196\,
            I => \N__13190\
        );

    \I__2124\ : Odrv12
    port map (
            O => \N__13193\,
            I => scaler_4_data_11
        );

    \I__2123\ : Odrv4
    port map (
            O => \N__13190\,
            I => scaler_4_data_11
        );

    \I__2122\ : InMux
    port map (
            O => \N__13185\,
            I => \N__13182\
        );

    \I__2121\ : LocalMux
    port map (
            O => \N__13182\,
            I => \N__13179\
        );

    \I__2120\ : Span4Mux_v
    port map (
            O => \N__13179\,
            I => \N__13176\
        );

    \I__2119\ : Odrv4
    port map (
            O => \N__13176\,
            I => \ppm_encoder_1.un1_rudder_cry_10_THRU_CO\
        );

    \I__2118\ : CascadeMux
    port map (
            O => \N__13173\,
            I => \N__13169\
        );

    \I__2117\ : InMux
    port map (
            O => \N__13172\,
            I => \N__13165\
        );

    \I__2116\ : InMux
    port map (
            O => \N__13169\,
            I => \N__13162\
        );

    \I__2115\ : CascadeMux
    port map (
            O => \N__13168\,
            I => \N__13158\
        );

    \I__2114\ : LocalMux
    port map (
            O => \N__13165\,
            I => \N__13149\
        );

    \I__2113\ : LocalMux
    port map (
            O => \N__13162\,
            I => \N__13149\
        );

    \I__2112\ : InMux
    port map (
            O => \N__13161\,
            I => \N__13140\
        );

    \I__2111\ : InMux
    port map (
            O => \N__13158\,
            I => \N__13140\
        );

    \I__2110\ : InMux
    port map (
            O => \N__13157\,
            I => \N__13140\
        );

    \I__2109\ : InMux
    port map (
            O => \N__13156\,
            I => \N__13140\
        );

    \I__2108\ : InMux
    port map (
            O => \N__13155\,
            I => \N__13137\
        );

    \I__2107\ : InMux
    port map (
            O => \N__13154\,
            I => \N__13134\
        );

    \I__2106\ : Span4Mux_v
    port map (
            O => \N__13149\,
            I => \N__13131\
        );

    \I__2105\ : LocalMux
    port map (
            O => \N__13140\,
            I => \N__13128\
        );

    \I__2104\ : LocalMux
    port map (
            O => \N__13137\,
            I => \uart_frame_decoder.state_1Z0Z_10\
        );

    \I__2103\ : LocalMux
    port map (
            O => \N__13134\,
            I => \uart_frame_decoder.state_1Z0Z_10\
        );

    \I__2102\ : Odrv4
    port map (
            O => \N__13131\,
            I => \uart_frame_decoder.state_1Z0Z_10\
        );

    \I__2101\ : Odrv4
    port map (
            O => \N__13128\,
            I => \uart_frame_decoder.state_1Z0Z_10\
        );

    \I__2100\ : CascadeMux
    port map (
            O => \N__13119\,
            I => \N__13113\
        );

    \I__2099\ : InMux
    port map (
            O => \N__13118\,
            I => \N__13107\
        );

    \I__2098\ : InMux
    port map (
            O => \N__13117\,
            I => \N__13103\
        );

    \I__2097\ : InMux
    port map (
            O => \N__13116\,
            I => \N__13100\
        );

    \I__2096\ : InMux
    port map (
            O => \N__13113\,
            I => \N__13094\
        );

    \I__2095\ : InMux
    port map (
            O => \N__13112\,
            I => \N__13094\
        );

    \I__2094\ : InMux
    port map (
            O => \N__13111\,
            I => \N__13084\
        );

    \I__2093\ : InMux
    port map (
            O => \N__13110\,
            I => \N__13084\
        );

    \I__2092\ : LocalMux
    port map (
            O => \N__13107\,
            I => \N__13081\
        );

    \I__2091\ : InMux
    port map (
            O => \N__13106\,
            I => \N__13078\
        );

    \I__2090\ : LocalMux
    port map (
            O => \N__13103\,
            I => \N__13075\
        );

    \I__2089\ : LocalMux
    port map (
            O => \N__13100\,
            I => \N__13072\
        );

    \I__2088\ : InMux
    port map (
            O => \N__13099\,
            I => \N__13069\
        );

    \I__2087\ : LocalMux
    port map (
            O => \N__13094\,
            I => \N__13066\
        );

    \I__2086\ : InMux
    port map (
            O => \N__13093\,
            I => \N__13063\
        );

    \I__2085\ : InMux
    port map (
            O => \N__13092\,
            I => \N__13054\
        );

    \I__2084\ : InMux
    port map (
            O => \N__13091\,
            I => \N__13054\
        );

    \I__2083\ : InMux
    port map (
            O => \N__13090\,
            I => \N__13054\
        );

    \I__2082\ : InMux
    port map (
            O => \N__13089\,
            I => \N__13051\
        );

    \I__2081\ : LocalMux
    port map (
            O => \N__13084\,
            I => \N__13044\
        );

    \I__2080\ : Span4Mux_s3_h
    port map (
            O => \N__13081\,
            I => \N__13044\
        );

    \I__2079\ : LocalMux
    port map (
            O => \N__13078\,
            I => \N__13044\
        );

    \I__2078\ : Span4Mux_v
    port map (
            O => \N__13075\,
            I => \N__13039\
        );

    \I__2077\ : Span4Mux_v
    port map (
            O => \N__13072\,
            I => \N__13039\
        );

    \I__2076\ : LocalMux
    port map (
            O => \N__13069\,
            I => \N__13032\
        );

    \I__2075\ : Span4Mux_h
    port map (
            O => \N__13066\,
            I => \N__13032\
        );

    \I__2074\ : LocalMux
    port map (
            O => \N__13063\,
            I => \N__13032\
        );

    \I__2073\ : InMux
    port map (
            O => \N__13062\,
            I => \N__13027\
        );

    \I__2072\ : InMux
    port map (
            O => \N__13061\,
            I => \N__13027\
        );

    \I__2071\ : LocalMux
    port map (
            O => \N__13054\,
            I => \N__13020\
        );

    \I__2070\ : LocalMux
    port map (
            O => \N__13051\,
            I => \N__13020\
        );

    \I__2069\ : Span4Mux_v
    port map (
            O => \N__13044\,
            I => \N__13020\
        );

    \I__2068\ : Odrv4
    port map (
            O => \N__13039\,
            I => uart_data_rdy
        );

    \I__2067\ : Odrv4
    port map (
            O => \N__13032\,
            I => uart_data_rdy
        );

    \I__2066\ : LocalMux
    port map (
            O => \N__13027\,
            I => uart_data_rdy
        );

    \I__2065\ : Odrv4
    port map (
            O => \N__13020\,
            I => uart_data_rdy
        );

    \I__2064\ : InMux
    port map (
            O => \N__13011\,
            I => \N__13008\
        );

    \I__2063\ : LocalMux
    port map (
            O => \N__13008\,
            I => \N__13005\
        );

    \I__2062\ : Span4Mux_v
    port map (
            O => \N__13005\,
            I => \N__13001\
        );

    \I__2061\ : InMux
    port map (
            O => \N__13004\,
            I => \N__12998\
        );

    \I__2060\ : Odrv4
    port map (
            O => \N__13001\,
            I => \uart_frame_decoder.count8_THRU_CO\
        );

    \I__2059\ : LocalMux
    port map (
            O => \N__12998\,
            I => \uart_frame_decoder.count8_THRU_CO\
        );

    \I__2058\ : InMux
    port map (
            O => \N__12993\,
            I => \N__12987\
        );

    \I__2057\ : InMux
    port map (
            O => \N__12992\,
            I => \N__12987\
        );

    \I__2056\ : LocalMux
    port map (
            O => \N__12987\,
            I => \N__12982\
        );

    \I__2055\ : CascadeMux
    port map (
            O => \N__12986\,
            I => \N__12978\
        );

    \I__2054\ : InMux
    port map (
            O => \N__12985\,
            I => \N__12970\
        );

    \I__2053\ : Span4Mux_h
    port map (
            O => \N__12982\,
            I => \N__12967\
        );

    \I__2052\ : InMux
    port map (
            O => \N__12981\,
            I => \N__12964\
        );

    \I__2051\ : InMux
    port map (
            O => \N__12978\,
            I => \N__12961\
        );

    \I__2050\ : InMux
    port map (
            O => \N__12977\,
            I => \N__12950\
        );

    \I__2049\ : InMux
    port map (
            O => \N__12976\,
            I => \N__12950\
        );

    \I__2048\ : InMux
    port map (
            O => \N__12975\,
            I => \N__12950\
        );

    \I__2047\ : InMux
    port map (
            O => \N__12974\,
            I => \N__12950\
        );

    \I__2046\ : InMux
    port map (
            O => \N__12973\,
            I => \N__12950\
        );

    \I__2045\ : LocalMux
    port map (
            O => \N__12970\,
            I => \uart.bit_CountZ0Z_2\
        );

    \I__2044\ : Odrv4
    port map (
            O => \N__12967\,
            I => \uart.bit_CountZ0Z_2\
        );

    \I__2043\ : LocalMux
    port map (
            O => \N__12964\,
            I => \uart.bit_CountZ0Z_2\
        );

    \I__2042\ : LocalMux
    port map (
            O => \N__12961\,
            I => \uart.bit_CountZ0Z_2\
        );

    \I__2041\ : LocalMux
    port map (
            O => \N__12950\,
            I => \uart.bit_CountZ0Z_2\
        );

    \I__2040\ : CascadeMux
    port map (
            O => \N__12939\,
            I => \N__12936\
        );

    \I__2039\ : InMux
    port map (
            O => \N__12936\,
            I => \N__12930\
        );

    \I__2038\ : InMux
    port map (
            O => \N__12935\,
            I => \N__12930\
        );

    \I__2037\ : LocalMux
    port map (
            O => \N__12930\,
            I => \N__12926\
        );

    \I__2036\ : InMux
    port map (
            O => \N__12929\,
            I => \N__12915\
        );

    \I__2035\ : Span4Mux_h
    port map (
            O => \N__12926\,
            I => \N__12912\
        );

    \I__2034\ : InMux
    port map (
            O => \N__12925\,
            I => \N__12907\
        );

    \I__2033\ : InMux
    port map (
            O => \N__12924\,
            I => \N__12907\
        );

    \I__2032\ : InMux
    port map (
            O => \N__12923\,
            I => \N__12904\
        );

    \I__2031\ : InMux
    port map (
            O => \N__12922\,
            I => \N__12899\
        );

    \I__2030\ : InMux
    port map (
            O => \N__12921\,
            I => \N__12899\
        );

    \I__2029\ : InMux
    port map (
            O => \N__12920\,
            I => \N__12892\
        );

    \I__2028\ : InMux
    port map (
            O => \N__12919\,
            I => \N__12892\
        );

    \I__2027\ : InMux
    port map (
            O => \N__12918\,
            I => \N__12892\
        );

    \I__2026\ : LocalMux
    port map (
            O => \N__12915\,
            I => \uart.bit_CountZ0Z_1\
        );

    \I__2025\ : Odrv4
    port map (
            O => \N__12912\,
            I => \uart.bit_CountZ0Z_1\
        );

    \I__2024\ : LocalMux
    port map (
            O => \N__12907\,
            I => \uart.bit_CountZ0Z_1\
        );

    \I__2023\ : LocalMux
    port map (
            O => \N__12904\,
            I => \uart.bit_CountZ0Z_1\
        );

    \I__2022\ : LocalMux
    port map (
            O => \N__12899\,
            I => \uart.bit_CountZ0Z_1\
        );

    \I__2021\ : LocalMux
    port map (
            O => \N__12892\,
            I => \uart.bit_CountZ0Z_1\
        );

    \I__2020\ : InMux
    port map (
            O => \N__12879\,
            I => \N__12871\
        );

    \I__2019\ : InMux
    port map (
            O => \N__12878\,
            I => \N__12871\
        );

    \I__2018\ : InMux
    port map (
            O => \N__12877\,
            I => \N__12866\
        );

    \I__2017\ : InMux
    port map (
            O => \N__12876\,
            I => \N__12866\
        );

    \I__2016\ : LocalMux
    port map (
            O => \N__12871\,
            I => \N__12863\
        );

    \I__2015\ : LocalMux
    port map (
            O => \N__12866\,
            I => \N__12850\
        );

    \I__2014\ : Span4Mux_v
    port map (
            O => \N__12863\,
            I => \N__12850\
        );

    \I__2013\ : InMux
    port map (
            O => \N__12862\,
            I => \N__12847\
        );

    \I__2012\ : InMux
    port map (
            O => \N__12861\,
            I => \N__12842\
        );

    \I__2011\ : InMux
    port map (
            O => \N__12860\,
            I => \N__12842\
        );

    \I__2010\ : InMux
    port map (
            O => \N__12859\,
            I => \N__12831\
        );

    \I__2009\ : InMux
    port map (
            O => \N__12858\,
            I => \N__12831\
        );

    \I__2008\ : InMux
    port map (
            O => \N__12857\,
            I => \N__12831\
        );

    \I__2007\ : InMux
    port map (
            O => \N__12856\,
            I => \N__12831\
        );

    \I__2006\ : InMux
    port map (
            O => \N__12855\,
            I => \N__12831\
        );

    \I__2005\ : Odrv4
    port map (
            O => \N__12850\,
            I => \uart.bit_CountZ0Z_0\
        );

    \I__2004\ : LocalMux
    port map (
            O => \N__12847\,
            I => \uart.bit_CountZ0Z_0\
        );

    \I__2003\ : LocalMux
    port map (
            O => \N__12842\,
            I => \uart.bit_CountZ0Z_0\
        );

    \I__2002\ : LocalMux
    port map (
            O => \N__12831\,
            I => \uart.bit_CountZ0Z_0\
        );

    \I__2001\ : InMux
    port map (
            O => \N__12822\,
            I => \N__12819\
        );

    \I__2000\ : LocalMux
    port map (
            O => \N__12819\,
            I => \uart.data_Auxce_0_0_2\
        );

    \I__1999\ : InMux
    port map (
            O => \N__12816\,
            I => \N__12813\
        );

    \I__1998\ : LocalMux
    port map (
            O => \N__12813\,
            I => \N__12810\
        );

    \I__1997\ : Odrv4
    port map (
            O => \N__12810\,
            I => \reset_module_System.reset6_13\
        );

    \I__1996\ : InMux
    port map (
            O => \N__12807\,
            I => \N__12804\
        );

    \I__1995\ : LocalMux
    port map (
            O => \N__12804\,
            I => \reset_module_System.reset6_3\
        );

    \I__1994\ : InMux
    port map (
            O => \N__12801\,
            I => \N__12798\
        );

    \I__1993\ : LocalMux
    port map (
            O => \N__12798\,
            I => \N__12795\
        );

    \I__1992\ : Odrv4
    port map (
            O => \N__12795\,
            I => \reset_module_System.reset6_17\
        );

    \I__1991\ : InMux
    port map (
            O => \N__12792\,
            I => \N__12789\
        );

    \I__1990\ : LocalMux
    port map (
            O => \N__12789\,
            I => \N__12783\
        );

    \I__1989\ : InMux
    port map (
            O => \N__12788\,
            I => \N__12780\
        );

    \I__1988\ : InMux
    port map (
            O => \N__12787\,
            I => \N__12774\
        );

    \I__1987\ : InMux
    port map (
            O => \N__12786\,
            I => \N__12771\
        );

    \I__1986\ : Span4Mux_s1_v
    port map (
            O => \N__12783\,
            I => \N__12766\
        );

    \I__1985\ : LocalMux
    port map (
            O => \N__12780\,
            I => \N__12766\
        );

    \I__1984\ : InMux
    port map (
            O => \N__12779\,
            I => \N__12763\
        );

    \I__1983\ : InMux
    port map (
            O => \N__12778\,
            I => \N__12760\
        );

    \I__1982\ : InMux
    port map (
            O => \N__12777\,
            I => \N__12757\
        );

    \I__1981\ : LocalMux
    port map (
            O => \N__12774\,
            I => \N__12752\
        );

    \I__1980\ : LocalMux
    port map (
            O => \N__12771\,
            I => \N__12752\
        );

    \I__1979\ : Span4Mux_v
    port map (
            O => \N__12766\,
            I => \N__12745\
        );

    \I__1978\ : LocalMux
    port map (
            O => \N__12763\,
            I => \N__12745\
        );

    \I__1977\ : LocalMux
    port map (
            O => \N__12760\,
            I => \N__12745\
        );

    \I__1976\ : LocalMux
    port map (
            O => \N__12757\,
            I => \N__12742\
        );

    \I__1975\ : Span12Mux_s10_v
    port map (
            O => \N__12752\,
            I => \N__12736\
        );

    \I__1974\ : Span4Mux_v
    port map (
            O => \N__12745\,
            I => \N__12731\
        );

    \I__1973\ : Span4Mux_s3_h
    port map (
            O => \N__12742\,
            I => \N__12731\
        );

    \I__1972\ : InMux
    port map (
            O => \N__12741\,
            I => \N__12728\
        );

    \I__1971\ : InMux
    port map (
            O => \N__12740\,
            I => \N__12725\
        );

    \I__1970\ : InMux
    port map (
            O => \N__12739\,
            I => \N__12722\
        );

    \I__1969\ : Odrv12
    port map (
            O => \N__12736\,
            I => uart_data_1
        );

    \I__1968\ : Odrv4
    port map (
            O => \N__12731\,
            I => uart_data_1
        );

    \I__1967\ : LocalMux
    port map (
            O => \N__12728\,
            I => uart_data_1
        );

    \I__1966\ : LocalMux
    port map (
            O => \N__12725\,
            I => uart_data_1
        );

    \I__1965\ : LocalMux
    port map (
            O => \N__12722\,
            I => uart_data_1
        );

    \I__1964\ : CascadeMux
    port map (
            O => \N__12711\,
            I => \uart_frame_decoder.state_1_ns_0_i_a2_1_1Z0Z_2_cascade_\
        );

    \I__1963\ : CascadeMux
    port map (
            O => \N__12708\,
            I => \N__12705\
        );

    \I__1962\ : InMux
    port map (
            O => \N__12705\,
            I => \N__12699\
        );

    \I__1961\ : InMux
    port map (
            O => \N__12704\,
            I => \N__12699\
        );

    \I__1960\ : LocalMux
    port map (
            O => \N__12699\,
            I => \N__12695\
        );

    \I__1959\ : InMux
    port map (
            O => \N__12698\,
            I => \N__12692\
        );

    \I__1958\ : Span4Mux_h
    port map (
            O => \N__12695\,
            I => \N__12689\
        );

    \I__1957\ : LocalMux
    port map (
            O => \N__12692\,
            I => \N__12686\
        );

    \I__1956\ : Odrv4
    port map (
            O => \N__12689\,
            I => \uart_frame_decoder.state_1_ns_0_i_a2_1Z0Z_2\
        );

    \I__1955\ : Odrv4
    port map (
            O => \N__12686\,
            I => \uart_frame_decoder.state_1_ns_0_i_a2_1Z0Z_2\
        );

    \I__1954\ : InMux
    port map (
            O => \N__12681\,
            I => \N__12677\
        );

    \I__1953\ : InMux
    port map (
            O => \N__12680\,
            I => \N__12674\
        );

    \I__1952\ : LocalMux
    port map (
            O => \N__12677\,
            I => \N__12671\
        );

    \I__1951\ : LocalMux
    port map (
            O => \N__12674\,
            I => \uart.stateZ0Z_0\
        );

    \I__1950\ : Odrv4
    port map (
            O => \N__12671\,
            I => \uart.stateZ0Z_0\
        );

    \I__1949\ : CascadeMux
    port map (
            O => \N__12666\,
            I => \N__12663\
        );

    \I__1948\ : InMux
    port map (
            O => \N__12663\,
            I => \N__12660\
        );

    \I__1947\ : LocalMux
    port map (
            O => \N__12660\,
            I => \N__12655\
        );

    \I__1946\ : InMux
    port map (
            O => \N__12659\,
            I => \N__12652\
        );

    \I__1945\ : InMux
    port map (
            O => \N__12658\,
            I => \N__12649\
        );

    \I__1944\ : Sp12to4
    port map (
            O => \N__12655\,
            I => \N__12644\
        );

    \I__1943\ : LocalMux
    port map (
            O => \N__12652\,
            I => \N__12644\
        );

    \I__1942\ : LocalMux
    port map (
            O => \N__12649\,
            I => \uart.stateZ0Z_1\
        );

    \I__1941\ : Odrv12
    port map (
            O => \N__12644\,
            I => \uart.stateZ0Z_1\
        );

    \I__1940\ : CascadeMux
    port map (
            O => \N__12639\,
            I => \N__12634\
        );

    \I__1939\ : CascadeMux
    port map (
            O => \N__12638\,
            I => \N__12623\
        );

    \I__1938\ : CascadeMux
    port map (
            O => \N__12637\,
            I => \N__12620\
        );

    \I__1937\ : InMux
    port map (
            O => \N__12634\,
            I => \N__12603\
        );

    \I__1936\ : InMux
    port map (
            O => \N__12633\,
            I => \N__12603\
        );

    \I__1935\ : InMux
    port map (
            O => \N__12632\,
            I => \N__12603\
        );

    \I__1934\ : InMux
    port map (
            O => \N__12631\,
            I => \N__12603\
        );

    \I__1933\ : InMux
    port map (
            O => \N__12630\,
            I => \N__12603\
        );

    \I__1932\ : InMux
    port map (
            O => \N__12629\,
            I => \N__12603\
        );

    \I__1931\ : InMux
    port map (
            O => \N__12628\,
            I => \N__12603\
        );

    \I__1930\ : InMux
    port map (
            O => \N__12627\,
            I => \N__12603\
        );

    \I__1929\ : InMux
    port map (
            O => \N__12626\,
            I => \N__12600\
        );

    \I__1928\ : InMux
    port map (
            O => \N__12623\,
            I => \N__12596\
        );

    \I__1927\ : InMux
    port map (
            O => \N__12620\,
            I => \N__12592\
        );

    \I__1926\ : LocalMux
    port map (
            O => \N__12603\,
            I => \N__12587\
        );

    \I__1925\ : LocalMux
    port map (
            O => \N__12600\,
            I => \N__12587\
        );

    \I__1924\ : InMux
    port map (
            O => \N__12599\,
            I => \N__12584\
        );

    \I__1923\ : LocalMux
    port map (
            O => \N__12596\,
            I => \N__12581\
        );

    \I__1922\ : InMux
    port map (
            O => \N__12595\,
            I => \N__12578\
        );

    \I__1921\ : LocalMux
    port map (
            O => \N__12592\,
            I => \N__12571\
        );

    \I__1920\ : Sp12to4
    port map (
            O => \N__12587\,
            I => \N__12571\
        );

    \I__1919\ : LocalMux
    port map (
            O => \N__12584\,
            I => \N__12571\
        );

    \I__1918\ : Odrv4
    port map (
            O => \N__12581\,
            I => uart_input_sync
        );

    \I__1917\ : LocalMux
    port map (
            O => \N__12578\,
            I => uart_input_sync
        );

    \I__1916\ : Odrv12
    port map (
            O => \N__12571\,
            I => uart_input_sync
        );

    \I__1915\ : InMux
    port map (
            O => \N__12564\,
            I => \N__12560\
        );

    \I__1914\ : CascadeMux
    port map (
            O => \N__12563\,
            I => \N__12557\
        );

    \I__1913\ : LocalMux
    port map (
            O => \N__12560\,
            I => \N__12554\
        );

    \I__1912\ : InMux
    port map (
            O => \N__12557\,
            I => \N__12551\
        );

    \I__1911\ : Odrv4
    port map (
            O => \N__12554\,
            I => \uart.data_AuxZ0Z_3\
        );

    \I__1910\ : LocalMux
    port map (
            O => \N__12551\,
            I => \uart.data_AuxZ0Z_3\
        );

    \I__1909\ : InMux
    port map (
            O => \N__12546\,
            I => \N__12540\
        );

    \I__1908\ : InMux
    port map (
            O => \N__12545\,
            I => \N__12537\
        );

    \I__1907\ : InMux
    port map (
            O => \N__12544\,
            I => \N__12534\
        );

    \I__1906\ : InMux
    port map (
            O => \N__12543\,
            I => \N__12531\
        );

    \I__1905\ : LocalMux
    port map (
            O => \N__12540\,
            I => \N__12519\
        );

    \I__1904\ : LocalMux
    port map (
            O => \N__12537\,
            I => \N__12519\
        );

    \I__1903\ : LocalMux
    port map (
            O => \N__12534\,
            I => \N__12519\
        );

    \I__1902\ : LocalMux
    port map (
            O => \N__12531\,
            I => \N__12519\
        );

    \I__1901\ : InMux
    port map (
            O => \N__12530\,
            I => \N__12516\
        );

    \I__1900\ : InMux
    port map (
            O => \N__12529\,
            I => \N__12513\
        );

    \I__1899\ : InMux
    port map (
            O => \N__12528\,
            I => \N__12510\
        );

    \I__1898\ : Span4Mux_v
    port map (
            O => \N__12519\,
            I => \N__12500\
        );

    \I__1897\ : LocalMux
    port map (
            O => \N__12516\,
            I => \N__12500\
        );

    \I__1896\ : LocalMux
    port map (
            O => \N__12513\,
            I => \N__12500\
        );

    \I__1895\ : LocalMux
    port map (
            O => \N__12510\,
            I => \N__12500\
        );

    \I__1894\ : InMux
    port map (
            O => \N__12509\,
            I => \N__12497\
        );

    \I__1893\ : Span4Mux_v
    port map (
            O => \N__12500\,
            I => \N__12490\
        );

    \I__1892\ : LocalMux
    port map (
            O => \N__12497\,
            I => \N__12490\
        );

    \I__1891\ : InMux
    port map (
            O => \N__12496\,
            I => \N__12487\
        );

    \I__1890\ : InMux
    port map (
            O => \N__12495\,
            I => \N__12484\
        );

    \I__1889\ : Odrv4
    port map (
            O => \N__12490\,
            I => uart_data_3
        );

    \I__1888\ : LocalMux
    port map (
            O => \N__12487\,
            I => uart_data_3
        );

    \I__1887\ : LocalMux
    port map (
            O => \N__12484\,
            I => uart_data_3
        );

    \I__1886\ : InMux
    port map (
            O => \N__12477\,
            I => \N__12474\
        );

    \I__1885\ : LocalMux
    port map (
            O => \N__12474\,
            I => \N__12471\
        );

    \I__1884\ : Span4Mux_v
    port map (
            O => \N__12471\,
            I => \N__12467\
        );

    \I__1883\ : InMux
    port map (
            O => \N__12470\,
            I => \N__12464\
        );

    \I__1882\ : Odrv4
    port map (
            O => \N__12467\,
            I => \uart.data_AuxZ0Z_6\
        );

    \I__1881\ : LocalMux
    port map (
            O => \N__12464\,
            I => \uart.data_AuxZ0Z_6\
        );

    \I__1880\ : InMux
    port map (
            O => \N__12459\,
            I => \N__12452\
        );

    \I__1879\ : InMux
    port map (
            O => \N__12458\,
            I => \N__12449\
        );

    \I__1878\ : InMux
    port map (
            O => \N__12457\,
            I => \N__12446\
        );

    \I__1877\ : InMux
    port map (
            O => \N__12456\,
            I => \N__12443\
        );

    \I__1876\ : InMux
    port map (
            O => \N__12455\,
            I => \N__12440\
        );

    \I__1875\ : LocalMux
    port map (
            O => \N__12452\,
            I => \N__12435\
        );

    \I__1874\ : LocalMux
    port map (
            O => \N__12449\,
            I => \N__12432\
        );

    \I__1873\ : LocalMux
    port map (
            O => \N__12446\,
            I => \N__12427\
        );

    \I__1872\ : LocalMux
    port map (
            O => \N__12443\,
            I => \N__12427\
        );

    \I__1871\ : LocalMux
    port map (
            O => \N__12440\,
            I => \N__12424\
        );

    \I__1870\ : InMux
    port map (
            O => \N__12439\,
            I => \N__12421\
        );

    \I__1869\ : InMux
    port map (
            O => \N__12438\,
            I => \N__12418\
        );

    \I__1868\ : Span4Mux_v
    port map (
            O => \N__12435\,
            I => \N__12414\
        );

    \I__1867\ : Span4Mux_h
    port map (
            O => \N__12432\,
            I => \N__12411\
        );

    \I__1866\ : Span4Mux_v
    port map (
            O => \N__12427\,
            I => \N__12402\
        );

    \I__1865\ : Span4Mux_h
    port map (
            O => \N__12424\,
            I => \N__12402\
        );

    \I__1864\ : LocalMux
    port map (
            O => \N__12421\,
            I => \N__12402\
        );

    \I__1863\ : LocalMux
    port map (
            O => \N__12418\,
            I => \N__12402\
        );

    \I__1862\ : InMux
    port map (
            O => \N__12417\,
            I => \N__12399\
        );

    \I__1861\ : Span4Mux_v
    port map (
            O => \N__12414\,
            I => \N__12394\
        );

    \I__1860\ : Span4Mux_v
    port map (
            O => \N__12411\,
            I => \N__12391\
        );

    \I__1859\ : Span4Mux_v
    port map (
            O => \N__12402\,
            I => \N__12386\
        );

    \I__1858\ : LocalMux
    port map (
            O => \N__12399\,
            I => \N__12386\
        );

    \I__1857\ : InMux
    port map (
            O => \N__12398\,
            I => \N__12383\
        );

    \I__1856\ : InMux
    port map (
            O => \N__12397\,
            I => \N__12380\
        );

    \I__1855\ : Odrv4
    port map (
            O => \N__12394\,
            I => uart_data_6
        );

    \I__1854\ : Odrv4
    port map (
            O => \N__12391\,
            I => uart_data_6
        );

    \I__1853\ : Odrv4
    port map (
            O => \N__12386\,
            I => uart_data_6
        );

    \I__1852\ : LocalMux
    port map (
            O => \N__12383\,
            I => uart_data_6
        );

    \I__1851\ : LocalMux
    port map (
            O => \N__12380\,
            I => uart_data_6
        );

    \I__1850\ : CascadeMux
    port map (
            O => \N__12369\,
            I => \reset_module_System.reset6_11_cascade_\
        );

    \I__1849\ : InMux
    port map (
            O => \N__12366\,
            I => \N__12361\
        );

    \I__1848\ : InMux
    port map (
            O => \N__12365\,
            I => \N__12356\
        );

    \I__1847\ : InMux
    port map (
            O => \N__12364\,
            I => \N__12356\
        );

    \I__1846\ : LocalMux
    port map (
            O => \N__12361\,
            I => \reset_module_System.reset6_19\
        );

    \I__1845\ : LocalMux
    port map (
            O => \N__12356\,
            I => \reset_module_System.reset6_19\
        );

    \I__1844\ : CascadeMux
    port map (
            O => \N__12351\,
            I => \reset_module_System.reset6_19_cascade_\
        );

    \I__1843\ : InMux
    port map (
            O => \N__12348\,
            I => \N__12345\
        );

    \I__1842\ : LocalMux
    port map (
            O => \N__12345\,
            I => \uart.data_Auxce_0_0_4\
        );

    \I__1841\ : InMux
    port map (
            O => \N__12342\,
            I => \N__12334\
        );

    \I__1840\ : InMux
    port map (
            O => \N__12341\,
            I => \N__12334\
        );

    \I__1839\ : InMux
    port map (
            O => \N__12340\,
            I => \N__12329\
        );

    \I__1838\ : InMux
    port map (
            O => \N__12339\,
            I => \N__12329\
        );

    \I__1837\ : LocalMux
    port map (
            O => \N__12334\,
            I => \N__12326\
        );

    \I__1836\ : LocalMux
    port map (
            O => \N__12329\,
            I => \reset_module_System.reset6_14\
        );

    \I__1835\ : Odrv4
    port map (
            O => \N__12326\,
            I => \reset_module_System.reset6_14\
        );

    \I__1834\ : SRMux
    port map (
            O => \N__12321\,
            I => \N__12318\
        );

    \I__1833\ : LocalMux
    port map (
            O => \N__12318\,
            I => \N__12315\
        );

    \I__1832\ : Odrv12
    port map (
            O => \N__12315\,
            I => \uart.state_RNIAFHLZ0Z_3\
        );

    \I__1831\ : InMux
    port map (
            O => \N__12312\,
            I => \N__12306\
        );

    \I__1830\ : InMux
    port map (
            O => \N__12311\,
            I => \N__12303\
        );

    \I__1829\ : InMux
    port map (
            O => \N__12310\,
            I => \N__12300\
        );

    \I__1828\ : InMux
    port map (
            O => \N__12309\,
            I => \N__12297\
        );

    \I__1827\ : LocalMux
    port map (
            O => \N__12306\,
            I => \N__12292\
        );

    \I__1826\ : LocalMux
    port map (
            O => \N__12303\,
            I => \N__12292\
        );

    \I__1825\ : LocalMux
    port map (
            O => \N__12300\,
            I => \uart.N_153_0\
        );

    \I__1824\ : LocalMux
    port map (
            O => \N__12297\,
            I => \uart.N_153_0\
        );

    \I__1823\ : Odrv4
    port map (
            O => \N__12292\,
            I => \uart.N_153_0\
        );

    \I__1822\ : InMux
    port map (
            O => \N__12285\,
            I => \N__12281\
        );

    \I__1821\ : InMux
    port map (
            O => \N__12284\,
            I => \N__12278\
        );

    \I__1820\ : LocalMux
    port map (
            O => \N__12281\,
            I => \N__12267\
        );

    \I__1819\ : LocalMux
    port map (
            O => \N__12278\,
            I => \N__12267\
        );

    \I__1818\ : InMux
    port map (
            O => \N__12277\,
            I => \N__12264\
        );

    \I__1817\ : InMux
    port map (
            O => \N__12276\,
            I => \N__12261\
        );

    \I__1816\ : InMux
    port map (
            O => \N__12275\,
            I => \N__12258\
        );

    \I__1815\ : InMux
    port map (
            O => \N__12274\,
            I => \N__12255\
        );

    \I__1814\ : InMux
    port map (
            O => \N__12273\,
            I => \N__12250\
        );

    \I__1813\ : InMux
    port map (
            O => \N__12272\,
            I => \N__12250\
        );

    \I__1812\ : Odrv4
    port map (
            O => \N__12267\,
            I => \uart.stateZ0Z_3\
        );

    \I__1811\ : LocalMux
    port map (
            O => \N__12264\,
            I => \uart.stateZ0Z_3\
        );

    \I__1810\ : LocalMux
    port map (
            O => \N__12261\,
            I => \uart.stateZ0Z_3\
        );

    \I__1809\ : LocalMux
    port map (
            O => \N__12258\,
            I => \uart.stateZ0Z_3\
        );

    \I__1808\ : LocalMux
    port map (
            O => \N__12255\,
            I => \uart.stateZ0Z_3\
        );

    \I__1807\ : LocalMux
    port map (
            O => \N__12250\,
            I => \uart.stateZ0Z_3\
        );

    \I__1806\ : CascadeMux
    port map (
            O => \N__12237\,
            I => \N__12234\
        );

    \I__1805\ : InMux
    port map (
            O => \N__12234\,
            I => \N__12231\
        );

    \I__1804\ : LocalMux
    port map (
            O => \N__12231\,
            I => \N__12228\
        );

    \I__1803\ : Odrv4
    port map (
            O => \N__12228\,
            I => \uart.N_168_1\
        );

    \I__1802\ : InMux
    port map (
            O => \N__12225\,
            I => \N__12222\
        );

    \I__1801\ : LocalMux
    port map (
            O => \N__12222\,
            I => \N__12219\
        );

    \I__1800\ : Odrv4
    port map (
            O => \N__12219\,
            I => \uart.N_167\
        );

    \I__1799\ : CascadeMux
    port map (
            O => \N__12216\,
            I => \N__12210\
        );

    \I__1798\ : CascadeMux
    port map (
            O => \N__12215\,
            I => \N__12203\
        );

    \I__1797\ : InMux
    port map (
            O => \N__12214\,
            I => \N__12197\
        );

    \I__1796\ : InMux
    port map (
            O => \N__12213\,
            I => \N__12197\
        );

    \I__1795\ : InMux
    port map (
            O => \N__12210\,
            I => \N__12192\
        );

    \I__1794\ : InMux
    port map (
            O => \N__12209\,
            I => \N__12192\
        );

    \I__1793\ : InMux
    port map (
            O => \N__12208\,
            I => \N__12189\
        );

    \I__1792\ : InMux
    port map (
            O => \N__12207\,
            I => \N__12186\
        );

    \I__1791\ : InMux
    port map (
            O => \N__12206\,
            I => \N__12183\
        );

    \I__1790\ : InMux
    port map (
            O => \N__12203\,
            I => \N__12180\
        );

    \I__1789\ : InMux
    port map (
            O => \N__12202\,
            I => \N__12177\
        );

    \I__1788\ : LocalMux
    port map (
            O => \N__12197\,
            I => \N__12174\
        );

    \I__1787\ : LocalMux
    port map (
            O => \N__12192\,
            I => \N__12171\
        );

    \I__1786\ : LocalMux
    port map (
            O => \N__12189\,
            I => \uart.stateZ0Z_4\
        );

    \I__1785\ : LocalMux
    port map (
            O => \N__12186\,
            I => \uart.stateZ0Z_4\
        );

    \I__1784\ : LocalMux
    port map (
            O => \N__12183\,
            I => \uart.stateZ0Z_4\
        );

    \I__1783\ : LocalMux
    port map (
            O => \N__12180\,
            I => \uart.stateZ0Z_4\
        );

    \I__1782\ : LocalMux
    port map (
            O => \N__12177\,
            I => \uart.stateZ0Z_4\
        );

    \I__1781\ : Odrv4
    port map (
            O => \N__12174\,
            I => \uart.stateZ0Z_4\
        );

    \I__1780\ : Odrv4
    port map (
            O => \N__12171\,
            I => \uart.stateZ0Z_4\
        );

    \I__1779\ : CascadeMux
    port map (
            O => \N__12156\,
            I => \reset_module_System.count_1_1_cascade_\
        );

    \I__1778\ : CascadeMux
    port map (
            O => \N__12153\,
            I => \uart.N_153_0_cascade_\
        );

    \I__1777\ : CascadeMux
    port map (
            O => \N__12150\,
            I => \uart.state_srsts_i_a3_0_0_3_cascade_\
        );

    \I__1776\ : InMux
    port map (
            O => \N__12147\,
            I => \N__12144\
        );

    \I__1775\ : LocalMux
    port map (
            O => \N__12144\,
            I => \uart.N_170\
        );

    \I__1774\ : InMux
    port map (
            O => \N__12141\,
            I => \N__12138\
        );

    \I__1773\ : LocalMux
    port map (
            O => \N__12138\,
            I => \uart.un1_state_2_0_a3_2\
        );

    \I__1772\ : InMux
    port map (
            O => \N__12135\,
            I => \N__12132\
        );

    \I__1771\ : LocalMux
    port map (
            O => \N__12132\,
            I => \N__12128\
        );

    \I__1770\ : InMux
    port map (
            O => \N__12131\,
            I => \N__12125\
        );

    \I__1769\ : Odrv4
    port map (
            O => \N__12128\,
            I => \uart.N_146_0\
        );

    \I__1768\ : LocalMux
    port map (
            O => \N__12125\,
            I => \uart.N_146_0\
        );

    \I__1767\ : InMux
    port map (
            O => \N__12120\,
            I => \N__12096\
        );

    \I__1766\ : InMux
    port map (
            O => \N__12119\,
            I => \N__12096\
        );

    \I__1765\ : InMux
    port map (
            O => \N__12118\,
            I => \N__12096\
        );

    \I__1764\ : InMux
    port map (
            O => \N__12117\,
            I => \N__12096\
        );

    \I__1763\ : InMux
    port map (
            O => \N__12116\,
            I => \N__12096\
        );

    \I__1762\ : InMux
    port map (
            O => \N__12115\,
            I => \N__12096\
        );

    \I__1761\ : InMux
    port map (
            O => \N__12114\,
            I => \N__12096\
        );

    \I__1760\ : InMux
    port map (
            O => \N__12113\,
            I => \N__12096\
        );

    \I__1759\ : LocalMux
    port map (
            O => \N__12096\,
            I => \uart.un1_state_2_0\
        );

    \I__1758\ : InMux
    port map (
            O => \N__12093\,
            I => \N__12090\
        );

    \I__1757\ : LocalMux
    port map (
            O => \N__12090\,
            I => \uart.N_151\
        );

    \I__1756\ : InMux
    port map (
            O => \N__12087\,
            I => \N__12081\
        );

    \I__1755\ : InMux
    port map (
            O => \N__12086\,
            I => \N__12078\
        );

    \I__1754\ : InMux
    port map (
            O => \N__12085\,
            I => \N__12075\
        );

    \I__1753\ : InMux
    port map (
            O => \N__12084\,
            I => \N__12072\
        );

    \I__1752\ : LocalMux
    port map (
            O => \N__12081\,
            I => \uart.stateZ0Z_2\
        );

    \I__1751\ : LocalMux
    port map (
            O => \N__12078\,
            I => \uart.stateZ0Z_2\
        );

    \I__1750\ : LocalMux
    port map (
            O => \N__12075\,
            I => \uart.stateZ0Z_2\
        );

    \I__1749\ : LocalMux
    port map (
            O => \N__12072\,
            I => \uart.stateZ0Z_2\
        );

    \I__1748\ : InMux
    port map (
            O => \N__12063\,
            I => \N__12060\
        );

    \I__1747\ : LocalMux
    port map (
            O => \N__12060\,
            I => \uart.N_159\
        );

    \I__1746\ : CascadeMux
    port map (
            O => \N__12057\,
            I => \uart.timer_Count_0_sqmuxa_1_cascade_\
        );

    \I__1745\ : InMux
    port map (
            O => \N__12054\,
            I => \N__12048\
        );

    \I__1744\ : InMux
    port map (
            O => \N__12053\,
            I => \N__12048\
        );

    \I__1743\ : LocalMux
    port map (
            O => \N__12048\,
            I => \uart.N_180\
        );

    \I__1742\ : CascadeMux
    port map (
            O => \N__12045\,
            I => \uart.N_180_cascade_\
        );

    \I__1741\ : InMux
    port map (
            O => \N__12042\,
            I => \N__12033\
        );

    \I__1740\ : InMux
    port map (
            O => \N__12041\,
            I => \N__12033\
        );

    \I__1739\ : InMux
    port map (
            O => \N__12040\,
            I => \N__12033\
        );

    \I__1738\ : LocalMux
    port map (
            O => \N__12033\,
            I => \N__12029\
        );

    \I__1737\ : InMux
    port map (
            O => \N__12032\,
            I => \N__12026\
        );

    \I__1736\ : Odrv4
    port map (
            O => \N__12029\,
            I => \uart.un1_state_5_0\
        );

    \I__1735\ : LocalMux
    port map (
            O => \N__12026\,
            I => \uart.un1_state_5_0\
        );

    \I__1734\ : InMux
    port map (
            O => \N__12021\,
            I => \N__12017\
        );

    \I__1733\ : InMux
    port map (
            O => \N__12020\,
            I => \N__12014\
        );

    \I__1732\ : LocalMux
    port map (
            O => \N__12017\,
            I => \uart.N_143_0\
        );

    \I__1731\ : LocalMux
    port map (
            O => \N__12014\,
            I => \uart.N_143_0\
        );

    \I__1730\ : CascadeMux
    port map (
            O => \N__12009\,
            I => \N__12006\
        );

    \I__1729\ : InMux
    port map (
            O => \N__12006\,
            I => \N__12000\
        );

    \I__1728\ : InMux
    port map (
            O => \N__12005\,
            I => \N__12000\
        );

    \I__1727\ : LocalMux
    port map (
            O => \N__12000\,
            I => \scaler_1.un3_source_data_0_cry_6_c_RNI1HI11\
        );

    \I__1726\ : InMux
    port map (
            O => \N__11997\,
            I => \scaler_1.un2_source_data_0_cry_7\
        );

    \I__1725\ : InMux
    port map (
            O => \N__11994\,
            I => \N__11990\
        );

    \I__1724\ : InMux
    port map (
            O => \N__11993\,
            I => \N__11987\
        );

    \I__1723\ : LocalMux
    port map (
            O => \N__11990\,
            I => \scaler_1.un3_source_data_0_cry_7_c_RNI2JJ11\
        );

    \I__1722\ : LocalMux
    port map (
            O => \N__11987\,
            I => \scaler_1.un3_source_data_0_cry_7_c_RNI2JJ11\
        );

    \I__1721\ : CascadeMux
    port map (
            O => \N__11982\,
            I => \N__11979\
        );

    \I__1720\ : InMux
    port map (
            O => \N__11979\,
            I => \N__11976\
        );

    \I__1719\ : LocalMux
    port map (
            O => \N__11976\,
            I => \scaler_1.un3_source_data_0_cry_8_c_RNIPB6F\
        );

    \I__1718\ : InMux
    port map (
            O => \N__11973\,
            I => \bfn_3_29_0_\
        );

    \I__1717\ : InMux
    port map (
            O => \N__11970\,
            I => \scaler_1.un2_source_data_0_cry_9\
        );

    \I__1716\ : CEMux
    port map (
            O => \N__11967\,
            I => \N__11940\
        );

    \I__1715\ : CEMux
    port map (
            O => \N__11966\,
            I => \N__11940\
        );

    \I__1714\ : CEMux
    port map (
            O => \N__11965\,
            I => \N__11940\
        );

    \I__1713\ : CEMux
    port map (
            O => \N__11964\,
            I => \N__11940\
        );

    \I__1712\ : CEMux
    port map (
            O => \N__11963\,
            I => \N__11940\
        );

    \I__1711\ : CEMux
    port map (
            O => \N__11962\,
            I => \N__11940\
        );

    \I__1710\ : CEMux
    port map (
            O => \N__11961\,
            I => \N__11940\
        );

    \I__1709\ : CEMux
    port map (
            O => \N__11960\,
            I => \N__11940\
        );

    \I__1708\ : CEMux
    port map (
            O => \N__11959\,
            I => \N__11940\
        );

    \I__1707\ : GlobalMux
    port map (
            O => \N__11940\,
            I => \N__11937\
        );

    \I__1706\ : gio2CtrlBuf
    port map (
            O => \N__11937\,
            I => frame_decoder_dv_c_0_g
        );

    \I__1705\ : CascadeMux
    port map (
            O => \N__11934\,
            I => \N__11931\
        );

    \I__1704\ : InMux
    port map (
            O => \N__11931\,
            I => \N__11928\
        );

    \I__1703\ : LocalMux
    port map (
            O => \N__11928\,
            I => \N__11925\
        );

    \I__1702\ : Span4Mux_s3_h
    port map (
            O => \N__11925\,
            I => \N__11922\
        );

    \I__1701\ : Span4Mux_v
    port map (
            O => \N__11922\,
            I => \N__11919\
        );

    \I__1700\ : Odrv4
    port map (
            O => \N__11919\,
            I => \frame_decoder_OFF3data_1\
        );

    \I__1699\ : CEMux
    port map (
            O => \N__11916\,
            I => \N__11913\
        );

    \I__1698\ : LocalMux
    port map (
            O => \N__11913\,
            I => \N__11909\
        );

    \I__1697\ : CEMux
    port map (
            O => \N__11912\,
            I => \N__11906\
        );

    \I__1696\ : Span4Mux_v
    port map (
            O => \N__11909\,
            I => \N__11903\
        );

    \I__1695\ : LocalMux
    port map (
            O => \N__11906\,
            I => \N__11900\
        );

    \I__1694\ : Odrv4
    port map (
            O => \N__11903\,
            I => \uart_frame_decoder.source_offset3data_1_sqmuxa_0\
        );

    \I__1693\ : Odrv4
    port map (
            O => \N__11900\,
            I => \uart_frame_decoder.source_offset3data_1_sqmuxa_0\
        );

    \I__1692\ : InMux
    port map (
            O => \N__11895\,
            I => \N__11892\
        );

    \I__1691\ : LocalMux
    port map (
            O => \N__11892\,
            I => \uart_sync.aux_2__0_Z0Z_0\
        );

    \I__1690\ : InMux
    port map (
            O => \N__11889\,
            I => \N__11886\
        );

    \I__1689\ : LocalMux
    port map (
            O => \N__11886\,
            I => \N__11883\
        );

    \I__1688\ : Odrv12
    port map (
            O => \N__11883\,
            I => \uart_sync.aux_3__0_Z0Z_0\
        );

    \I__1687\ : InMux
    port map (
            O => \N__11880\,
            I => \N__11877\
        );

    \I__1686\ : LocalMux
    port map (
            O => \N__11877\,
            I => \N__11874\
        );

    \I__1685\ : Odrv4
    port map (
            O => \N__11874\,
            I => scaler_4_data_14
        );

    \I__1684\ : InMux
    port map (
            O => \N__11871\,
            I => \bfn_3_27_0_\
        );

    \I__1683\ : CascadeMux
    port map (
            O => \N__11868\,
            I => \N__11865\
        );

    \I__1682\ : InMux
    port map (
            O => \N__11865\,
            I => \N__11862\
        );

    \I__1681\ : LocalMux
    port map (
            O => \N__11862\,
            I => \scaler_1.un2_source_data_0_cry_1_c_RNOZ0\
        );

    \I__1680\ : InMux
    port map (
            O => \N__11859\,
            I => \N__11854\
        );

    \I__1679\ : CascadeMux
    port map (
            O => \N__11858\,
            I => \N__11851\
        );

    \I__1678\ : InMux
    port map (
            O => \N__11857\,
            I => \N__11847\
        );

    \I__1677\ : LocalMux
    port map (
            O => \N__11854\,
            I => \N__11844\
        );

    \I__1676\ : InMux
    port map (
            O => \N__11851\,
            I => \N__11839\
        );

    \I__1675\ : InMux
    port map (
            O => \N__11850\,
            I => \N__11839\
        );

    \I__1674\ : LocalMux
    port map (
            O => \N__11847\,
            I => \scaler_1.un2_source_data_0\
        );

    \I__1673\ : Odrv4
    port map (
            O => \N__11844\,
            I => \scaler_1.un2_source_data_0\
        );

    \I__1672\ : LocalMux
    port map (
            O => \N__11839\,
            I => \scaler_1.un2_source_data_0\
        );

    \I__1671\ : InMux
    port map (
            O => \N__11832\,
            I => \scaler_1.un2_source_data_0_cry_1\
        );

    \I__1670\ : CascadeMux
    port map (
            O => \N__11829\,
            I => \N__11826\
        );

    \I__1669\ : InMux
    port map (
            O => \N__11826\,
            I => \N__11820\
        );

    \I__1668\ : InMux
    port map (
            O => \N__11825\,
            I => \N__11820\
        );

    \I__1667\ : LocalMux
    port map (
            O => \N__11820\,
            I => \scaler_1.un3_source_data_0_cry_1_c_RNIISC11\
        );

    \I__1666\ : InMux
    port map (
            O => \N__11817\,
            I => \scaler_1.un2_source_data_0_cry_2\
        );

    \I__1665\ : CascadeMux
    port map (
            O => \N__11814\,
            I => \N__11811\
        );

    \I__1664\ : InMux
    port map (
            O => \N__11811\,
            I => \N__11805\
        );

    \I__1663\ : InMux
    port map (
            O => \N__11810\,
            I => \N__11805\
        );

    \I__1662\ : LocalMux
    port map (
            O => \N__11805\,
            I => \scaler_1.un3_source_data_0_cry_2_c_RNIL0E11\
        );

    \I__1661\ : InMux
    port map (
            O => \N__11802\,
            I => \scaler_1.un2_source_data_0_cry_3\
        );

    \I__1660\ : CascadeMux
    port map (
            O => \N__11799\,
            I => \N__11796\
        );

    \I__1659\ : InMux
    port map (
            O => \N__11796\,
            I => \N__11790\
        );

    \I__1658\ : InMux
    port map (
            O => \N__11795\,
            I => \N__11790\
        );

    \I__1657\ : LocalMux
    port map (
            O => \N__11790\,
            I => \scaler_1.un3_source_data_0_cry_3_c_RNIO4F11\
        );

    \I__1656\ : InMux
    port map (
            O => \N__11787\,
            I => \scaler_1.un2_source_data_0_cry_4\
        );

    \I__1655\ : CascadeMux
    port map (
            O => \N__11784\,
            I => \N__11781\
        );

    \I__1654\ : InMux
    port map (
            O => \N__11781\,
            I => \N__11775\
        );

    \I__1653\ : InMux
    port map (
            O => \N__11780\,
            I => \N__11775\
        );

    \I__1652\ : LocalMux
    port map (
            O => \N__11775\,
            I => \scaler_1.un3_source_data_0_cry_4_c_RNIR8G11\
        );

    \I__1651\ : InMux
    port map (
            O => \N__11772\,
            I => \scaler_1.un2_source_data_0_cry_5\
        );

    \I__1650\ : CascadeMux
    port map (
            O => \N__11769\,
            I => \N__11766\
        );

    \I__1649\ : InMux
    port map (
            O => \N__11766\,
            I => \N__11760\
        );

    \I__1648\ : InMux
    port map (
            O => \N__11765\,
            I => \N__11760\
        );

    \I__1647\ : LocalMux
    port map (
            O => \N__11760\,
            I => \scaler_1.un3_source_data_0_cry_5_c_RNIUCH11\
        );

    \I__1646\ : InMux
    port map (
            O => \N__11757\,
            I => \scaler_1.un2_source_data_0_cry_6\
        );

    \I__1645\ : InMux
    port map (
            O => \N__11754\,
            I => \N__11751\
        );

    \I__1644\ : LocalMux
    port map (
            O => \N__11751\,
            I => \N__11747\
        );

    \I__1643\ : InMux
    port map (
            O => \N__11750\,
            I => \N__11744\
        );

    \I__1642\ : Odrv4
    port map (
            O => \N__11747\,
            I => \frame_decoder_OFF1data_7\
        );

    \I__1641\ : LocalMux
    port map (
            O => \N__11744\,
            I => \frame_decoder_OFF1data_7\
        );

    \I__1640\ : InMux
    port map (
            O => \N__11739\,
            I => \N__11736\
        );

    \I__1639\ : LocalMux
    port map (
            O => \N__11736\,
            I => \N__11732\
        );

    \I__1638\ : InMux
    port map (
            O => \N__11735\,
            I => \N__11729\
        );

    \I__1637\ : Odrv4
    port map (
            O => \N__11732\,
            I => \frame_decoder_CH1data_7\
        );

    \I__1636\ : LocalMux
    port map (
            O => \N__11729\,
            I => \frame_decoder_CH1data_7\
        );

    \I__1635\ : CascadeMux
    port map (
            O => \N__11724\,
            I => \N__11721\
        );

    \I__1634\ : InMux
    port map (
            O => \N__11721\,
            I => \N__11718\
        );

    \I__1633\ : LocalMux
    port map (
            O => \N__11718\,
            I => \N__11715\
        );

    \I__1632\ : Odrv4
    port map (
            O => \N__11715\,
            I => \scaler_1.un3_source_data_0_axb_7\
        );

    \I__1631\ : InMux
    port map (
            O => \N__11712\,
            I => \ppm_encoder_1.un1_rudder_cry_6\
        );

    \I__1630\ : InMux
    port map (
            O => \N__11709\,
            I => \ppm_encoder_1.un1_rudder_cry_7\
        );

    \I__1629\ : InMux
    port map (
            O => \N__11706\,
            I => \ppm_encoder_1.un1_rudder_cry_8\
        );

    \I__1628\ : InMux
    port map (
            O => \N__11703\,
            I => \ppm_encoder_1.un1_rudder_cry_9\
        );

    \I__1627\ : InMux
    port map (
            O => \N__11700\,
            I => \ppm_encoder_1.un1_rudder_cry_10\
        );

    \I__1626\ : InMux
    port map (
            O => \N__11697\,
            I => \ppm_encoder_1.un1_rudder_cry_11\
        );

    \I__1625\ : InMux
    port map (
            O => \N__11694\,
            I => \ppm_encoder_1.un1_rudder_cry_12\
        );

    \I__1624\ : InMux
    port map (
            O => \N__11691\,
            I => \N__11687\
        );

    \I__1623\ : CascadeMux
    port map (
            O => \N__11690\,
            I => \N__11684\
        );

    \I__1622\ : LocalMux
    port map (
            O => \N__11687\,
            I => \N__11679\
        );

    \I__1621\ : InMux
    port map (
            O => \N__11684\,
            I => \N__11674\
        );

    \I__1620\ : InMux
    port map (
            O => \N__11683\,
            I => \N__11674\
        );

    \I__1619\ : InMux
    port map (
            O => \N__11682\,
            I => \N__11671\
        );

    \I__1618\ : Span4Mux_v
    port map (
            O => \N__11679\,
            I => \N__11668\
        );

    \I__1617\ : LocalMux
    port map (
            O => \N__11674\,
            I => \N__11665\
        );

    \I__1616\ : LocalMux
    port map (
            O => \N__11671\,
            I => \scaler_3.un2_source_data_0\
        );

    \I__1615\ : Odrv4
    port map (
            O => \N__11668\,
            I => \scaler_3.un2_source_data_0\
        );

    \I__1614\ : Odrv4
    port map (
            O => \N__11665\,
            I => \scaler_3.un2_source_data_0\
        );

    \I__1613\ : InMux
    port map (
            O => \N__11658\,
            I => \N__11655\
        );

    \I__1612\ : LocalMux
    port map (
            O => \N__11655\,
            I => \N__11651\
        );

    \I__1611\ : InMux
    port map (
            O => \N__11654\,
            I => \N__11648\
        );

    \I__1610\ : Span4Mux_h
    port map (
            O => \N__11651\,
            I => \N__11643\
        );

    \I__1609\ : LocalMux
    port map (
            O => \N__11648\,
            I => \N__11643\
        );

    \I__1608\ : Span4Mux_v
    port map (
            O => \N__11643\,
            I => \N__11640\
        );

    \I__1607\ : Odrv4
    port map (
            O => \N__11640\,
            I => \uart_frame_decoder.source_offset2data_1_sqmuxa\
        );

    \I__1606\ : CascadeMux
    port map (
            O => \N__11637\,
            I => \N__11633\
        );

    \I__1605\ : InMux
    port map (
            O => \N__11636\,
            I => \N__11630\
        );

    \I__1604\ : InMux
    port map (
            O => \N__11633\,
            I => \N__11627\
        );

    \I__1603\ : LocalMux
    port map (
            O => \N__11630\,
            I => \uart_frame_decoder.state_1Z0Z_8\
        );

    \I__1602\ : LocalMux
    port map (
            O => \N__11627\,
            I => \uart_frame_decoder.state_1Z0Z_8\
        );

    \I__1601\ : InMux
    port map (
            O => \N__11622\,
            I => \N__11619\
        );

    \I__1600\ : LocalMux
    port map (
            O => \N__11619\,
            I => \uart_frame_decoder.source_offset3data_1_sqmuxa\
        );

    \I__1599\ : CascadeMux
    port map (
            O => \N__11616\,
            I => \N__11613\
        );

    \I__1598\ : InMux
    port map (
            O => \N__11613\,
            I => \N__11607\
        );

    \I__1597\ : InMux
    port map (
            O => \N__11612\,
            I => \N__11607\
        );

    \I__1596\ : LocalMux
    port map (
            O => \N__11607\,
            I => \uart_frame_decoder.state_1Z0Z_9\
        );

    \I__1595\ : InMux
    port map (
            O => \N__11604\,
            I => \N__11600\
        );

    \I__1594\ : InMux
    port map (
            O => \N__11603\,
            I => \N__11597\
        );

    \I__1593\ : LocalMux
    port map (
            O => \N__11600\,
            I => \uart_frame_decoder.state_1Z0Z_5\
        );

    \I__1592\ : LocalMux
    port map (
            O => \N__11597\,
            I => \uart_frame_decoder.state_1Z0Z_5\
        );

    \I__1591\ : InMux
    port map (
            O => \N__11592\,
            I => \N__11589\
        );

    \I__1590\ : LocalMux
    port map (
            O => \N__11589\,
            I => \uart_frame_decoder.source_CH4data_1_sqmuxa\
        );

    \I__1589\ : InMux
    port map (
            O => \N__11586\,
            I => \N__11577\
        );

    \I__1588\ : InMux
    port map (
            O => \N__11585\,
            I => \N__11574\
        );

    \I__1587\ : InMux
    port map (
            O => \N__11584\,
            I => \N__11571\
        );

    \I__1586\ : InMux
    port map (
            O => \N__11583\,
            I => \N__11567\
        );

    \I__1585\ : InMux
    port map (
            O => \N__11582\,
            I => \N__11564\
        );

    \I__1584\ : InMux
    port map (
            O => \N__11581\,
            I => \N__11561\
        );

    \I__1583\ : InMux
    port map (
            O => \N__11580\,
            I => \N__11558\
        );

    \I__1582\ : LocalMux
    port map (
            O => \N__11577\,
            I => \N__11555\
        );

    \I__1581\ : LocalMux
    port map (
            O => \N__11574\,
            I => \N__11548\
        );

    \I__1580\ : LocalMux
    port map (
            O => \N__11571\,
            I => \N__11548\
        );

    \I__1579\ : CascadeMux
    port map (
            O => \N__11570\,
            I => \N__11545\
        );

    \I__1578\ : LocalMux
    port map (
            O => \N__11567\,
            I => \N__11533\
        );

    \I__1577\ : LocalMux
    port map (
            O => \N__11564\,
            I => \N__11533\
        );

    \I__1576\ : LocalMux
    port map (
            O => \N__11561\,
            I => \N__11533\
        );

    \I__1575\ : LocalMux
    port map (
            O => \N__11558\,
            I => \N__11533\
        );

    \I__1574\ : Span4Mux_s3_h
    port map (
            O => \N__11555\,
            I => \N__11533\
        );

    \I__1573\ : InMux
    port map (
            O => \N__11554\,
            I => \N__11530\
        );

    \I__1572\ : InMux
    port map (
            O => \N__11553\,
            I => \N__11527\
        );

    \I__1571\ : Span4Mux_v
    port map (
            O => \N__11548\,
            I => \N__11524\
        );

    \I__1570\ : InMux
    port map (
            O => \N__11545\,
            I => \N__11519\
        );

    \I__1569\ : InMux
    port map (
            O => \N__11544\,
            I => \N__11519\
        );

    \I__1568\ : Span4Mux_v
    port map (
            O => \N__11533\,
            I => \N__11514\
        );

    \I__1567\ : LocalMux
    port map (
            O => \N__11530\,
            I => \N__11514\
        );

    \I__1566\ : LocalMux
    port map (
            O => \N__11527\,
            I => uart_data_7
        );

    \I__1565\ : Odrv4
    port map (
            O => \N__11524\,
            I => uart_data_7
        );

    \I__1564\ : LocalMux
    port map (
            O => \N__11519\,
            I => uart_data_7
        );

    \I__1563\ : Odrv4
    port map (
            O => \N__11514\,
            I => uart_data_7
        );

    \I__1562\ : InMux
    port map (
            O => \N__11505\,
            I => \N__11502\
        );

    \I__1561\ : LocalMux
    port map (
            O => \N__11502\,
            I => \N__11499\
        );

    \I__1560\ : Span4Mux_s2_v
    port map (
            O => \N__11499\,
            I => \N__11495\
        );

    \I__1559\ : InMux
    port map (
            O => \N__11498\,
            I => \N__11492\
        );

    \I__1558\ : Span4Mux_v
    port map (
            O => \N__11495\,
            I => \N__11487\
        );

    \I__1557\ : LocalMux
    port map (
            O => \N__11492\,
            I => \N__11487\
        );

    \I__1556\ : Odrv4
    port map (
            O => \N__11487\,
            I => \frame_decoder_CH4data_7\
        );

    \I__1555\ : CEMux
    port map (
            O => \N__11484\,
            I => \N__11481\
        );

    \I__1554\ : LocalMux
    port map (
            O => \N__11481\,
            I => \N__11478\
        );

    \I__1553\ : Span4Mux_s3_v
    port map (
            O => \N__11478\,
            I => \N__11474\
        );

    \I__1552\ : CEMux
    port map (
            O => \N__11477\,
            I => \N__11471\
        );

    \I__1551\ : Span4Mux_v
    port map (
            O => \N__11474\,
            I => \N__11468\
        );

    \I__1550\ : LocalMux
    port map (
            O => \N__11471\,
            I => \uart_frame_decoder.source_CH4data_1_sqmuxa_0\
        );

    \I__1549\ : Odrv4
    port map (
            O => \N__11468\,
            I => \uart_frame_decoder.source_CH4data_1_sqmuxa_0\
        );

    \I__1548\ : InMux
    port map (
            O => \N__11463\,
            I => \N__11460\
        );

    \I__1547\ : LocalMux
    port map (
            O => \N__11460\,
            I => \N__11456\
        );

    \I__1546\ : InMux
    port map (
            O => \N__11459\,
            I => \N__11453\
        );

    \I__1545\ : Span4Mux_v
    port map (
            O => \N__11456\,
            I => \N__11448\
        );

    \I__1544\ : LocalMux
    port map (
            O => \N__11453\,
            I => \N__11448\
        );

    \I__1543\ : Odrv4
    port map (
            O => \N__11448\,
            I => \uart_frame_decoder.source_CH3data_1_sqmuxa\
        );

    \I__1542\ : CEMux
    port map (
            O => \N__11445\,
            I => \N__11442\
        );

    \I__1541\ : LocalMux
    port map (
            O => \N__11442\,
            I => \uart_frame_decoder.source_CH3data_1_sqmuxa_0\
        );

    \I__1540\ : InMux
    port map (
            O => \N__11439\,
            I => \N__11436\
        );

    \I__1539\ : LocalMux
    port map (
            O => \N__11436\,
            I => \N__11431\
        );

    \I__1538\ : InMux
    port map (
            O => \N__11435\,
            I => \N__11427\
        );

    \I__1537\ : CascadeMux
    port map (
            O => \N__11434\,
            I => \N__11424\
        );

    \I__1536\ : Span4Mux_v
    port map (
            O => \N__11431\,
            I => \N__11421\
        );

    \I__1535\ : InMux
    port map (
            O => \N__11430\,
            I => \N__11418\
        );

    \I__1534\ : LocalMux
    port map (
            O => \N__11427\,
            I => \N__11415\
        );

    \I__1533\ : InMux
    port map (
            O => \N__11424\,
            I => \N__11412\
        );

    \I__1532\ : Odrv4
    port map (
            O => \N__11421\,
            I => \frame_decoder_OFF1data_0\
        );

    \I__1531\ : LocalMux
    port map (
            O => \N__11418\,
            I => \frame_decoder_OFF1data_0\
        );

    \I__1530\ : Odrv4
    port map (
            O => \N__11415\,
            I => \frame_decoder_OFF1data_0\
        );

    \I__1529\ : LocalMux
    port map (
            O => \N__11412\,
            I => \frame_decoder_OFF1data_0\
        );

    \I__1528\ : InMux
    port map (
            O => \N__11403\,
            I => \N__11399\
        );

    \I__1527\ : InMux
    port map (
            O => \N__11402\,
            I => \N__11396\
        );

    \I__1526\ : LocalMux
    port map (
            O => \N__11399\,
            I => \N__11391\
        );

    \I__1525\ : LocalMux
    port map (
            O => \N__11396\,
            I => \N__11388\
        );

    \I__1524\ : InMux
    port map (
            O => \N__11395\,
            I => \N__11385\
        );

    \I__1523\ : InMux
    port map (
            O => \N__11394\,
            I => \N__11382\
        );

    \I__1522\ : Span4Mux_v
    port map (
            O => \N__11391\,
            I => \N__11375\
        );

    \I__1521\ : Span4Mux_s3_v
    port map (
            O => \N__11388\,
            I => \N__11375\
        );

    \I__1520\ : LocalMux
    port map (
            O => \N__11385\,
            I => \N__11375\
        );

    \I__1519\ : LocalMux
    port map (
            O => \N__11382\,
            I => \frame_decoder_CH1data_0\
        );

    \I__1518\ : Odrv4
    port map (
            O => \N__11375\,
            I => \frame_decoder_CH1data_0\
        );

    \I__1517\ : CascadeMux
    port map (
            O => \N__11370\,
            I => \N__11367\
        );

    \I__1516\ : InMux
    port map (
            O => \N__11367\,
            I => \N__11361\
        );

    \I__1515\ : InMux
    port map (
            O => \N__11366\,
            I => \N__11361\
        );

    \I__1514\ : LocalMux
    port map (
            O => \N__11361\,
            I => \scaler_2.un3_source_data_0_cry_1_c_RNILSPH\
        );

    \I__1513\ : InMux
    port map (
            O => \N__11358\,
            I => \scaler_2.un2_source_data_0_cry_2\
        );

    \I__1512\ : CascadeMux
    port map (
            O => \N__11355\,
            I => \N__11352\
        );

    \I__1511\ : InMux
    port map (
            O => \N__11352\,
            I => \N__11346\
        );

    \I__1510\ : InMux
    port map (
            O => \N__11351\,
            I => \N__11346\
        );

    \I__1509\ : LocalMux
    port map (
            O => \N__11346\,
            I => \scaler_2.un3_source_data_0_cry_2_c_RNIO0RH\
        );

    \I__1508\ : InMux
    port map (
            O => \N__11343\,
            I => \scaler_2.un2_source_data_0_cry_3\
        );

    \I__1507\ : CascadeMux
    port map (
            O => \N__11340\,
            I => \N__11337\
        );

    \I__1506\ : InMux
    port map (
            O => \N__11337\,
            I => \N__11331\
        );

    \I__1505\ : InMux
    port map (
            O => \N__11336\,
            I => \N__11331\
        );

    \I__1504\ : LocalMux
    port map (
            O => \N__11331\,
            I => \scaler_2.un3_source_data_0_cry_3_c_RNIR4SH\
        );

    \I__1503\ : InMux
    port map (
            O => \N__11328\,
            I => \scaler_2.un2_source_data_0_cry_4\
        );

    \I__1502\ : CascadeMux
    port map (
            O => \N__11325\,
            I => \N__11322\
        );

    \I__1501\ : InMux
    port map (
            O => \N__11322\,
            I => \N__11316\
        );

    \I__1500\ : InMux
    port map (
            O => \N__11321\,
            I => \N__11316\
        );

    \I__1499\ : LocalMux
    port map (
            O => \N__11316\,
            I => \scaler_2.un3_source_data_0_cry_4_c_RNIU8TH\
        );

    \I__1498\ : InMux
    port map (
            O => \N__11313\,
            I => \scaler_2.un2_source_data_0_cry_5\
        );

    \I__1497\ : CascadeMux
    port map (
            O => \N__11310\,
            I => \N__11307\
        );

    \I__1496\ : InMux
    port map (
            O => \N__11307\,
            I => \N__11301\
        );

    \I__1495\ : InMux
    port map (
            O => \N__11306\,
            I => \N__11301\
        );

    \I__1494\ : LocalMux
    port map (
            O => \N__11301\,
            I => \scaler_2.un3_source_data_0_cry_5_c_RNI1DUH\
        );

    \I__1493\ : InMux
    port map (
            O => \N__11298\,
            I => \scaler_2.un2_source_data_0_cry_6\
        );

    \I__1492\ : CascadeMux
    port map (
            O => \N__11295\,
            I => \N__11292\
        );

    \I__1491\ : InMux
    port map (
            O => \N__11292\,
            I => \N__11286\
        );

    \I__1490\ : InMux
    port map (
            O => \N__11291\,
            I => \N__11286\
        );

    \I__1489\ : LocalMux
    port map (
            O => \N__11286\,
            I => \scaler_2.un3_source_data_0_cry_6_c_RNI4HVH\
        );

    \I__1488\ : InMux
    port map (
            O => \N__11283\,
            I => \scaler_2.un2_source_data_0_cry_7\
        );

    \I__1487\ : InMux
    port map (
            O => \N__11280\,
            I => \N__11276\
        );

    \I__1486\ : InMux
    port map (
            O => \N__11279\,
            I => \N__11273\
        );

    \I__1485\ : LocalMux
    port map (
            O => \N__11276\,
            I => \scaler_2.un3_source_data_0_cry_7_c_RNI5J0I\
        );

    \I__1484\ : LocalMux
    port map (
            O => \N__11273\,
            I => \scaler_2.un3_source_data_0_cry_7_c_RNI5J0I\
        );

    \I__1483\ : CascadeMux
    port map (
            O => \N__11268\,
            I => \N__11265\
        );

    \I__1482\ : InMux
    port map (
            O => \N__11265\,
            I => \N__11262\
        );

    \I__1481\ : LocalMux
    port map (
            O => \N__11262\,
            I => \scaler_2.un3_source_data_0_cry_8_c_RNIQL42\
        );

    \I__1480\ : InMux
    port map (
            O => \N__11259\,
            I => \bfn_3_22_0_\
        );

    \I__1479\ : InMux
    port map (
            O => \N__11256\,
            I => \scaler_2.un2_source_data_0_cry_9\
        );

    \I__1478\ : InMux
    port map (
            O => \N__11253\,
            I => \N__11249\
        );

    \I__1477\ : InMux
    port map (
            O => \N__11252\,
            I => \N__11246\
        );

    \I__1476\ : LocalMux
    port map (
            O => \N__11249\,
            I => \N__11236\
        );

    \I__1475\ : LocalMux
    port map (
            O => \N__11246\,
            I => \N__11236\
        );

    \I__1474\ : InMux
    port map (
            O => \N__11245\,
            I => \N__11233\
        );

    \I__1473\ : InMux
    port map (
            O => \N__11244\,
            I => \N__11230\
        );

    \I__1472\ : InMux
    port map (
            O => \N__11243\,
            I => \N__11227\
        );

    \I__1471\ : InMux
    port map (
            O => \N__11242\,
            I => \N__11224\
        );

    \I__1470\ : InMux
    port map (
            O => \N__11241\,
            I => \N__11221\
        );

    \I__1469\ : Span4Mux_v
    port map (
            O => \N__11236\,
            I => \N__11217\
        );

    \I__1468\ : LocalMux
    port map (
            O => \N__11233\,
            I => \N__11214\
        );

    \I__1467\ : LocalMux
    port map (
            O => \N__11230\,
            I => \N__11204\
        );

    \I__1466\ : LocalMux
    port map (
            O => \N__11227\,
            I => \N__11204\
        );

    \I__1465\ : LocalMux
    port map (
            O => \N__11224\,
            I => \N__11204\
        );

    \I__1464\ : LocalMux
    port map (
            O => \N__11221\,
            I => \N__11201\
        );

    \I__1463\ : InMux
    port map (
            O => \N__11220\,
            I => \N__11198\
        );

    \I__1462\ : Span4Mux_v
    port map (
            O => \N__11217\,
            I => \N__11195\
        );

    \I__1461\ : Span4Mux_s3_h
    port map (
            O => \N__11214\,
            I => \N__11192\
        );

    \I__1460\ : InMux
    port map (
            O => \N__11213\,
            I => \N__11189\
        );

    \I__1459\ : InMux
    port map (
            O => \N__11212\,
            I => \N__11184\
        );

    \I__1458\ : InMux
    port map (
            O => \N__11211\,
            I => \N__11184\
        );

    \I__1457\ : Span4Mux_v
    port map (
            O => \N__11204\,
            I => \N__11177\
        );

    \I__1456\ : Span4Mux_s3_h
    port map (
            O => \N__11201\,
            I => \N__11177\
        );

    \I__1455\ : LocalMux
    port map (
            O => \N__11198\,
            I => \N__11177\
        );

    \I__1454\ : Odrv4
    port map (
            O => \N__11195\,
            I => uart_data_0
        );

    \I__1453\ : Odrv4
    port map (
            O => \N__11192\,
            I => uart_data_0
        );

    \I__1452\ : LocalMux
    port map (
            O => \N__11189\,
            I => uart_data_0
        );

    \I__1451\ : LocalMux
    port map (
            O => \N__11184\,
            I => uart_data_0
        );

    \I__1450\ : Odrv4
    port map (
            O => \N__11177\,
            I => uart_data_0
        );

    \I__1449\ : InMux
    port map (
            O => \N__11166\,
            I => \N__11162\
        );

    \I__1448\ : CascadeMux
    port map (
            O => \N__11165\,
            I => \N__11158\
        );

    \I__1447\ : LocalMux
    port map (
            O => \N__11162\,
            I => \N__11155\
        );

    \I__1446\ : CascadeMux
    port map (
            O => \N__11161\,
            I => \N__11152\
        );

    \I__1445\ : InMux
    port map (
            O => \N__11158\,
            I => \N__11147\
        );

    \I__1444\ : Span4Mux_h
    port map (
            O => \N__11155\,
            I => \N__11144\
        );

    \I__1443\ : InMux
    port map (
            O => \N__11152\,
            I => \N__11137\
        );

    \I__1442\ : InMux
    port map (
            O => \N__11151\,
            I => \N__11137\
        );

    \I__1441\ : InMux
    port map (
            O => \N__11150\,
            I => \N__11137\
        );

    \I__1440\ : LocalMux
    port map (
            O => \N__11147\,
            I => \uart_frame_decoder.state_1Z0Z_1\
        );

    \I__1439\ : Odrv4
    port map (
            O => \N__11144\,
            I => \uart_frame_decoder.state_1Z0Z_1\
        );

    \I__1438\ : LocalMux
    port map (
            O => \N__11137\,
            I => \uart_frame_decoder.state_1Z0Z_1\
        );

    \I__1437\ : CascadeMux
    port map (
            O => \N__11130\,
            I => \uart_frame_decoder.state_1_ns_0_i_a2_0_0_1Z0Z_2_cascade_\
        );

    \I__1436\ : InMux
    port map (
            O => \N__11127\,
            I => \N__11124\
        );

    \I__1435\ : LocalMux
    port map (
            O => \N__11124\,
            I => \N__11120\
        );

    \I__1434\ : InMux
    port map (
            O => \N__11123\,
            I => \N__11117\
        );

    \I__1433\ : Odrv4
    port map (
            O => \N__11120\,
            I => \uart_frame_decoder.state_1_ns_0_i_a2_0_2\
        );

    \I__1432\ : LocalMux
    port map (
            O => \N__11117\,
            I => \uart_frame_decoder.state_1_ns_0_i_a2_0_2\
        );

    \I__1431\ : InMux
    port map (
            O => \N__11112\,
            I => \N__11108\
        );

    \I__1430\ : CascadeMux
    port map (
            O => \N__11111\,
            I => \N__11105\
        );

    \I__1429\ : LocalMux
    port map (
            O => \N__11108\,
            I => \N__11102\
        );

    \I__1428\ : InMux
    port map (
            O => \N__11105\,
            I => \N__11099\
        );

    \I__1427\ : Odrv4
    port map (
            O => \N__11102\,
            I => \uart.data_AuxZ0Z_5\
        );

    \I__1426\ : LocalMux
    port map (
            O => \N__11099\,
            I => \uart.data_AuxZ0Z_5\
        );

    \I__1425\ : InMux
    port map (
            O => \N__11094\,
            I => \N__11090\
        );

    \I__1424\ : InMux
    port map (
            O => \N__11093\,
            I => \N__11087\
        );

    \I__1423\ : LocalMux
    port map (
            O => \N__11090\,
            I => \N__11076\
        );

    \I__1422\ : LocalMux
    port map (
            O => \N__11087\,
            I => \N__11076\
        );

    \I__1421\ : InMux
    port map (
            O => \N__11086\,
            I => \N__11073\
        );

    \I__1420\ : InMux
    port map (
            O => \N__11085\,
            I => \N__11070\
        );

    \I__1419\ : InMux
    port map (
            O => \N__11084\,
            I => \N__11067\
        );

    \I__1418\ : InMux
    port map (
            O => \N__11083\,
            I => \N__11064\
        );

    \I__1417\ : InMux
    port map (
            O => \N__11082\,
            I => \N__11061\
        );

    \I__1416\ : CascadeMux
    port map (
            O => \N__11081\,
            I => \N__11058\
        );

    \I__1415\ : Span4Mux_v
    port map (
            O => \N__11076\,
            I => \N__11051\
        );

    \I__1414\ : LocalMux
    port map (
            O => \N__11073\,
            I => \N__11051\
        );

    \I__1413\ : LocalMux
    port map (
            O => \N__11070\,
            I => \N__11051\
        );

    \I__1412\ : LocalMux
    port map (
            O => \N__11067\,
            I => \N__11048\
        );

    \I__1411\ : LocalMux
    port map (
            O => \N__11064\,
            I => \N__11040\
        );

    \I__1410\ : LocalMux
    port map (
            O => \N__11061\,
            I => \N__11040\
        );

    \I__1409\ : InMux
    port map (
            O => \N__11058\,
            I => \N__11037\
        );

    \I__1408\ : Span4Mux_v
    port map (
            O => \N__11051\,
            I => \N__11034\
        );

    \I__1407\ : Span4Mux_s3_h
    port map (
            O => \N__11048\,
            I => \N__11031\
        );

    \I__1406\ : InMux
    port map (
            O => \N__11047\,
            I => \N__11028\
        );

    \I__1405\ : InMux
    port map (
            O => \N__11046\,
            I => \N__11023\
        );

    \I__1404\ : InMux
    port map (
            O => \N__11045\,
            I => \N__11023\
        );

    \I__1403\ : Span4Mux_v
    port map (
            O => \N__11040\,
            I => \N__11018\
        );

    \I__1402\ : LocalMux
    port map (
            O => \N__11037\,
            I => \N__11018\
        );

    \I__1401\ : Odrv4
    port map (
            O => \N__11034\,
            I => uart_data_5
        );

    \I__1400\ : Odrv4
    port map (
            O => \N__11031\,
            I => uart_data_5
        );

    \I__1399\ : LocalMux
    port map (
            O => \N__11028\,
            I => uart_data_5
        );

    \I__1398\ : LocalMux
    port map (
            O => \N__11023\,
            I => uart_data_5
        );

    \I__1397\ : Odrv4
    port map (
            O => \N__11018\,
            I => uart_data_5
        );

    \I__1396\ : InMux
    port map (
            O => \N__11007\,
            I => \N__11004\
        );

    \I__1395\ : LocalMux
    port map (
            O => \N__11004\,
            I => \N__11000\
        );

    \I__1394\ : CascadeMux
    port map (
            O => \N__11003\,
            I => \N__10997\
        );

    \I__1393\ : Span4Mux_v
    port map (
            O => \N__11000\,
            I => \N__10994\
        );

    \I__1392\ : InMux
    port map (
            O => \N__10997\,
            I => \N__10991\
        );

    \I__1391\ : Odrv4
    port map (
            O => \N__10994\,
            I => \uart.data_AuxZ1Z_2\
        );

    \I__1390\ : LocalMux
    port map (
            O => \N__10991\,
            I => \uart.data_AuxZ1Z_2\
        );

    \I__1389\ : InMux
    port map (
            O => \N__10986\,
            I => \N__10982\
        );

    \I__1388\ : InMux
    port map (
            O => \N__10985\,
            I => \N__10979\
        );

    \I__1387\ : LocalMux
    port map (
            O => \N__10982\,
            I => \N__10969\
        );

    \I__1386\ : LocalMux
    port map (
            O => \N__10979\,
            I => \N__10969\
        );

    \I__1385\ : InMux
    port map (
            O => \N__10978\,
            I => \N__10966\
        );

    \I__1384\ : InMux
    port map (
            O => \N__10977\,
            I => \N__10963\
        );

    \I__1383\ : InMux
    port map (
            O => \N__10976\,
            I => \N__10960\
        );

    \I__1382\ : InMux
    port map (
            O => \N__10975\,
            I => \N__10957\
        );

    \I__1381\ : InMux
    port map (
            O => \N__10974\,
            I => \N__10954\
        );

    \I__1380\ : Span4Mux_v
    port map (
            O => \N__10969\,
            I => \N__10946\
        );

    \I__1379\ : LocalMux
    port map (
            O => \N__10966\,
            I => \N__10946\
        );

    \I__1378\ : LocalMux
    port map (
            O => \N__10963\,
            I => \N__10946\
        );

    \I__1377\ : LocalMux
    port map (
            O => \N__10960\,
            I => \N__10936\
        );

    \I__1376\ : LocalMux
    port map (
            O => \N__10957\,
            I => \N__10936\
        );

    \I__1375\ : LocalMux
    port map (
            O => \N__10954\,
            I => \N__10936\
        );

    \I__1374\ : InMux
    port map (
            O => \N__10953\,
            I => \N__10933\
        );

    \I__1373\ : Span4Mux_v
    port map (
            O => \N__10946\,
            I => \N__10930\
        );

    \I__1372\ : InMux
    port map (
            O => \N__10945\,
            I => \N__10927\
        );

    \I__1371\ : InMux
    port map (
            O => \N__10944\,
            I => \N__10922\
        );

    \I__1370\ : InMux
    port map (
            O => \N__10943\,
            I => \N__10922\
        );

    \I__1369\ : Span4Mux_v
    port map (
            O => \N__10936\,
            I => \N__10917\
        );

    \I__1368\ : LocalMux
    port map (
            O => \N__10933\,
            I => \N__10917\
        );

    \I__1367\ : Odrv4
    port map (
            O => \N__10930\,
            I => uart_data_2
        );

    \I__1366\ : LocalMux
    port map (
            O => \N__10927\,
            I => uart_data_2
        );

    \I__1365\ : LocalMux
    port map (
            O => \N__10922\,
            I => uart_data_2
        );

    \I__1364\ : Odrv4
    port map (
            O => \N__10917\,
            I => uart_data_2
        );

    \I__1363\ : InMux
    port map (
            O => \N__10908\,
            I => \N__10905\
        );

    \I__1362\ : LocalMux
    port map (
            O => \N__10905\,
            I => \N__10901\
        );

    \I__1361\ : InMux
    port map (
            O => \N__10904\,
            I => \N__10898\
        );

    \I__1360\ : Odrv4
    port map (
            O => \N__10901\,
            I => \uart.data_AuxZ0Z_7\
        );

    \I__1359\ : LocalMux
    port map (
            O => \N__10898\,
            I => \uart.data_AuxZ0Z_7\
        );

    \I__1358\ : InMux
    port map (
            O => \N__10893\,
            I => \N__10890\
        );

    \I__1357\ : LocalMux
    port map (
            O => \N__10890\,
            I => \N__10886\
        );

    \I__1356\ : InMux
    port map (
            O => \N__10889\,
            I => \N__10883\
        );

    \I__1355\ : Odrv12
    port map (
            O => \N__10886\,
            I => \uart.data_AuxZ1Z_1\
        );

    \I__1354\ : LocalMux
    port map (
            O => \N__10883\,
            I => \uart.data_AuxZ1Z_1\
        );

    \I__1353\ : InMux
    port map (
            O => \N__10878\,
            I => \scaler_2.un2_source_data_0_cry_1\
        );

    \I__1352\ : CascadeMux
    port map (
            O => \N__10875\,
            I => \N__10872\
        );

    \I__1351\ : InMux
    port map (
            O => \N__10872\,
            I => \N__10869\
        );

    \I__1350\ : LocalMux
    port map (
            O => \N__10869\,
            I => \N__10866\
        );

    \I__1349\ : Odrv12
    port map (
            O => \N__10866\,
            I => \uart.N_177\
        );

    \I__1348\ : CascadeMux
    port map (
            O => \N__10863\,
            I => \uart.state_srsts_0_0_0_cascade_\
        );

    \I__1347\ : InMux
    port map (
            O => \N__10860\,
            I => \N__10857\
        );

    \I__1346\ : LocalMux
    port map (
            O => \N__10857\,
            I => \N__10853\
        );

    \I__1345\ : InMux
    port map (
            O => \N__10856\,
            I => \N__10850\
        );

    \I__1344\ : Odrv4
    port map (
            O => \N__10853\,
            I => \uart_frame_decoder.state_1_RNI592GZ0Z_10\
        );

    \I__1343\ : LocalMux
    port map (
            O => \N__10850\,
            I => \uart_frame_decoder.state_1_RNI592GZ0Z_10\
        );

    \I__1342\ : InMux
    port map (
            O => \N__10845\,
            I => \N__10842\
        );

    \I__1341\ : LocalMux
    port map (
            O => \N__10842\,
            I => \uart_frame_decoder.state_1_RNO_3Z0Z_0\
        );

    \I__1340\ : InMux
    port map (
            O => \N__10839\,
            I => \N__10836\
        );

    \I__1339\ : LocalMux
    port map (
            O => \N__10836\,
            I => \uart_frame_decoder.N_168_i_1\
        );

    \I__1338\ : CascadeMux
    port map (
            O => \N__10833\,
            I => \N__10830\
        );

    \I__1337\ : InMux
    port map (
            O => \N__10830\,
            I => \N__10827\
        );

    \I__1336\ : LocalMux
    port map (
            O => \N__10827\,
            I => \uart_frame_decoder.state_1_RNO_2Z0Z_0\
        );

    \I__1335\ : InMux
    port map (
            O => \N__10824\,
            I => \N__10820\
        );

    \I__1334\ : InMux
    port map (
            O => \N__10823\,
            I => \N__10817\
        );

    \I__1333\ : LocalMux
    port map (
            O => \N__10820\,
            I => \N__10814\
        );

    \I__1332\ : LocalMux
    port map (
            O => \N__10817\,
            I => \uart_frame_decoder.state_1Z0Z_7\
        );

    \I__1331\ : Odrv4
    port map (
            O => \N__10814\,
            I => \uart_frame_decoder.state_1Z0Z_7\
        );

    \I__1330\ : InMux
    port map (
            O => \N__10809\,
            I => \N__10800\
        );

    \I__1329\ : InMux
    port map (
            O => \N__10808\,
            I => \N__10800\
        );

    \I__1328\ : InMux
    port map (
            O => \N__10807\,
            I => \N__10800\
        );

    \I__1327\ : LocalMux
    port map (
            O => \N__10800\,
            I => \N__10797\
        );

    \I__1326\ : Odrv4
    port map (
            O => \N__10797\,
            I => \uart_frame_decoder.state_1Z0Z_0\
        );

    \I__1325\ : InMux
    port map (
            O => \N__10794\,
            I => \N__10788\
        );

    \I__1324\ : InMux
    port map (
            O => \N__10793\,
            I => \N__10788\
        );

    \I__1323\ : LocalMux
    port map (
            O => \N__10788\,
            I => \N__10785\
        );

    \I__1322\ : Span4Mux_v
    port map (
            O => \N__10785\,
            I => \N__10782\
        );

    \I__1321\ : Odrv4
    port map (
            O => \N__10782\,
            I => \uart_frame_decoder.N_79_4\
        );

    \I__1320\ : InMux
    port map (
            O => \N__10779\,
            I => \N__10776\
        );

    \I__1319\ : LocalMux
    port map (
            O => \N__10776\,
            I => \uart_frame_decoder.state_1_ns_0_i_a2_0_0_1\
        );

    \I__1318\ : InMux
    port map (
            O => \N__10773\,
            I => \N__10769\
        );

    \I__1317\ : CascadeMux
    port map (
            O => \N__10772\,
            I => \N__10766\
        );

    \I__1316\ : LocalMux
    port map (
            O => \N__10769\,
            I => \N__10763\
        );

    \I__1315\ : InMux
    port map (
            O => \N__10766\,
            I => \N__10760\
        );

    \I__1314\ : Odrv4
    port map (
            O => \N__10763\,
            I => \uart.data_AuxZ1Z_0\
        );

    \I__1313\ : LocalMux
    port map (
            O => \N__10760\,
            I => \uart.data_AuxZ1Z_0\
        );

    \I__1312\ : InMux
    port map (
            O => \N__10755\,
            I => \N__10752\
        );

    \I__1311\ : LocalMux
    port map (
            O => \N__10752\,
            I => \N__10749\
        );

    \I__1310\ : Odrv4
    port map (
            O => \N__10749\,
            I => \uart.data_Auxce_0_0_0\
        );

    \I__1309\ : CascadeMux
    port map (
            O => \N__10746\,
            I => \N__10743\
        );

    \I__1308\ : InMux
    port map (
            O => \N__10743\,
            I => \N__10740\
        );

    \I__1307\ : LocalMux
    port map (
            O => \N__10740\,
            I => \N__10737\
        );

    \I__1306\ : Odrv4
    port map (
            O => \N__10737\,
            I => \uart.data_Auxce_0_1\
        );

    \I__1305\ : InMux
    port map (
            O => \N__10734\,
            I => \N__10731\
        );

    \I__1304\ : LocalMux
    port map (
            O => \N__10731\,
            I => \N__10728\
        );

    \I__1303\ : Odrv4
    port map (
            O => \N__10728\,
            I => \uart.data_Auxce_0_3\
        );

    \I__1302\ : InMux
    port map (
            O => \N__10725\,
            I => \N__10722\
        );

    \I__1301\ : LocalMux
    port map (
            O => \N__10722\,
            I => \N__10719\
        );

    \I__1300\ : Odrv4
    port map (
            O => \N__10719\,
            I => \uart.data_Auxce_0_5\
        );

    \I__1299\ : InMux
    port map (
            O => \N__10716\,
            I => \N__10713\
        );

    \I__1298\ : LocalMux
    port map (
            O => \N__10713\,
            I => \N__10710\
        );

    \I__1297\ : Odrv4
    port map (
            O => \N__10710\,
            I => \uart.data_Auxce_0_6\
        );

    \I__1296\ : InMux
    port map (
            O => \N__10707\,
            I => \N__10704\
        );

    \I__1295\ : LocalMux
    port map (
            O => \N__10704\,
            I => \uart.CO1\
        );

    \I__1294\ : CascadeMux
    port map (
            O => \N__10701\,
            I => \N__10697\
        );

    \I__1293\ : CascadeMux
    port map (
            O => \N__10700\,
            I => \N__10694\
        );

    \I__1292\ : InMux
    port map (
            O => \N__10697\,
            I => \N__10686\
        );

    \I__1291\ : InMux
    port map (
            O => \N__10694\,
            I => \N__10686\
        );

    \I__1290\ : InMux
    port map (
            O => \N__10693\,
            I => \N__10686\
        );

    \I__1289\ : LocalMux
    port map (
            O => \N__10686\,
            I => \uart.N_133_0\
        );

    \I__1288\ : CascadeMux
    port map (
            O => \N__10683\,
            I => \uart.N_177_cascade_\
        );

    \I__1287\ : InMux
    port map (
            O => \N__10680\,
            I => \N__10677\
        );

    \I__1286\ : LocalMux
    port map (
            O => \N__10677\,
            I => \uart.state_srsts_i_0_3\
        );

    \I__1285\ : CascadeMux
    port map (
            O => \N__10674\,
            I => \uart.N_168_1_cascade_\
        );

    \I__1284\ : InMux
    port map (
            O => \N__10671\,
            I => \N__10668\
        );

    \I__1283\ : LocalMux
    port map (
            O => \N__10668\,
            I => \uart.N_154_0\
        );

    \I__1282\ : CascadeMux
    port map (
            O => \N__10665\,
            I => \N__10662\
        );

    \I__1281\ : InMux
    port map (
            O => \N__10662\,
            I => \N__10656\
        );

    \I__1280\ : InMux
    port map (
            O => \N__10661\,
            I => \N__10656\
        );

    \I__1279\ : LocalMux
    port map (
            O => \N__10656\,
            I => \scaler_4.un3_source_data_0_cry_1_c_RNIRSJI\
        );

    \I__1278\ : InMux
    port map (
            O => \N__10653\,
            I => \scaler_4.un2_source_data_0_cry_2\
        );

    \I__1277\ : CascadeMux
    port map (
            O => \N__10650\,
            I => \N__10647\
        );

    \I__1276\ : InMux
    port map (
            O => \N__10647\,
            I => \N__10641\
        );

    \I__1275\ : InMux
    port map (
            O => \N__10646\,
            I => \N__10641\
        );

    \I__1274\ : LocalMux
    port map (
            O => \N__10641\,
            I => \scaler_4.un3_source_data_0_cry_2_c_RNIU0LI\
        );

    \I__1273\ : InMux
    port map (
            O => \N__10638\,
            I => \scaler_4.un2_source_data_0_cry_3\
        );

    \I__1272\ : CascadeMux
    port map (
            O => \N__10635\,
            I => \N__10632\
        );

    \I__1271\ : InMux
    port map (
            O => \N__10632\,
            I => \N__10626\
        );

    \I__1270\ : InMux
    port map (
            O => \N__10631\,
            I => \N__10626\
        );

    \I__1269\ : LocalMux
    port map (
            O => \N__10626\,
            I => \scaler_4.un3_source_data_0_cry_3_c_RNI15MI\
        );

    \I__1268\ : InMux
    port map (
            O => \N__10623\,
            I => \scaler_4.un2_source_data_0_cry_4\
        );

    \I__1267\ : CascadeMux
    port map (
            O => \N__10620\,
            I => \N__10617\
        );

    \I__1266\ : InMux
    port map (
            O => \N__10617\,
            I => \N__10611\
        );

    \I__1265\ : InMux
    port map (
            O => \N__10616\,
            I => \N__10611\
        );

    \I__1264\ : LocalMux
    port map (
            O => \N__10611\,
            I => \scaler_4.un3_source_data_0_cry_4_c_RNI49NI\
        );

    \I__1263\ : InMux
    port map (
            O => \N__10608\,
            I => \scaler_4.un2_source_data_0_cry_5\
        );

    \I__1262\ : CascadeMux
    port map (
            O => \N__10605\,
            I => \N__10602\
        );

    \I__1261\ : InMux
    port map (
            O => \N__10602\,
            I => \N__10596\
        );

    \I__1260\ : InMux
    port map (
            O => \N__10601\,
            I => \N__10596\
        );

    \I__1259\ : LocalMux
    port map (
            O => \N__10596\,
            I => \scaler_4.un3_source_data_0_cry_5_c_RNI7DOI\
        );

    \I__1258\ : InMux
    port map (
            O => \N__10593\,
            I => \scaler_4.un2_source_data_0_cry_6\
        );

    \I__1257\ : CascadeMux
    port map (
            O => \N__10590\,
            I => \N__10587\
        );

    \I__1256\ : InMux
    port map (
            O => \N__10587\,
            I => \N__10581\
        );

    \I__1255\ : InMux
    port map (
            O => \N__10586\,
            I => \N__10581\
        );

    \I__1254\ : LocalMux
    port map (
            O => \N__10581\,
            I => \scaler_4.un3_source_data_0_cry_6_c_RNIAHPI\
        );

    \I__1253\ : InMux
    port map (
            O => \N__10578\,
            I => \scaler_4.un2_source_data_0_cry_7\
        );

    \I__1252\ : InMux
    port map (
            O => \N__10575\,
            I => \N__10571\
        );

    \I__1251\ : InMux
    port map (
            O => \N__10574\,
            I => \N__10568\
        );

    \I__1250\ : LocalMux
    port map (
            O => \N__10571\,
            I => \scaler_4.un3_source_data_0_cry_7_c_RNIBJQI\
        );

    \I__1249\ : LocalMux
    port map (
            O => \N__10568\,
            I => \scaler_4.un3_source_data_0_cry_7_c_RNIBJQI\
        );

    \I__1248\ : CascadeMux
    port map (
            O => \N__10563\,
            I => \N__10560\
        );

    \I__1247\ : InMux
    port map (
            O => \N__10560\,
            I => \N__10557\
        );

    \I__1246\ : LocalMux
    port map (
            O => \N__10557\,
            I => \scaler_4.un3_source_data_0_cry_8_c_RNIS918\
        );

    \I__1245\ : InMux
    port map (
            O => \N__10554\,
            I => \bfn_2_30_0_\
        );

    \I__1244\ : InMux
    port map (
            O => \N__10551\,
            I => \scaler_4.un2_source_data_0_cry_9\
        );

    \I__1243\ : InMux
    port map (
            O => \N__10548\,
            I => \N__10545\
        );

    \I__1242\ : LocalMux
    port map (
            O => \N__10545\,
            I => \frame_decoder_OFF1data_6\
        );

    \I__1241\ : CascadeMux
    port map (
            O => \N__10542\,
            I => \N__10539\
        );

    \I__1240\ : InMux
    port map (
            O => \N__10539\,
            I => \N__10536\
        );

    \I__1239\ : LocalMux
    port map (
            O => \N__10536\,
            I => \N__10533\
        );

    \I__1238\ : Odrv4
    port map (
            O => \N__10533\,
            I => \frame_decoder_CH1data_6\
        );

    \I__1237\ : InMux
    port map (
            O => \N__10530\,
            I => \scaler_1.un3_source_data_0_cry_5\
        );

    \I__1236\ : InMux
    port map (
            O => \N__10527\,
            I => \scaler_1.un3_source_data_0_cry_6\
        );

    \I__1235\ : InMux
    port map (
            O => \N__10524\,
            I => \bfn_2_28_0_\
        );

    \I__1234\ : InMux
    port map (
            O => \N__10521\,
            I => \scaler_1.un3_source_data_0_cry_8\
        );

    \I__1233\ : InMux
    port map (
            O => \N__10518\,
            I => \N__10515\
        );

    \I__1232\ : LocalMux
    port map (
            O => \N__10515\,
            I => \scaler_1.N_771_i_l_ofxZ0\
        );

    \I__1231\ : InMux
    port map (
            O => \N__10512\,
            I => \N__10508\
        );

    \I__1230\ : InMux
    port map (
            O => \N__10511\,
            I => \N__10505\
        );

    \I__1229\ : LocalMux
    port map (
            O => \N__10508\,
            I => \N__10500\
        );

    \I__1228\ : LocalMux
    port map (
            O => \N__10505\,
            I => \N__10497\
        );

    \I__1227\ : InMux
    port map (
            O => \N__10504\,
            I => \N__10494\
        );

    \I__1226\ : InMux
    port map (
            O => \N__10503\,
            I => \N__10491\
        );

    \I__1225\ : Odrv4
    port map (
            O => \N__10500\,
            I => \frame_decoder_CH4data_0\
        );

    \I__1224\ : Odrv12
    port map (
            O => \N__10497\,
            I => \frame_decoder_CH4data_0\
        );

    \I__1223\ : LocalMux
    port map (
            O => \N__10494\,
            I => \frame_decoder_CH4data_0\
        );

    \I__1222\ : LocalMux
    port map (
            O => \N__10491\,
            I => \frame_decoder_CH4data_0\
        );

    \I__1221\ : CascadeMux
    port map (
            O => \N__10482\,
            I => \N__10478\
        );

    \I__1220\ : InMux
    port map (
            O => \N__10481\,
            I => \N__10475\
        );

    \I__1219\ : InMux
    port map (
            O => \N__10478\,
            I => \N__10470\
        );

    \I__1218\ : LocalMux
    port map (
            O => \N__10475\,
            I => \N__10467\
        );

    \I__1217\ : InMux
    port map (
            O => \N__10474\,
            I => \N__10464\
        );

    \I__1216\ : InMux
    port map (
            O => \N__10473\,
            I => \N__10461\
        );

    \I__1215\ : LocalMux
    port map (
            O => \N__10470\,
            I => \N__10458\
        );

    \I__1214\ : Odrv12
    port map (
            O => \N__10467\,
            I => \frame_decoder_OFF4data_0\
        );

    \I__1213\ : LocalMux
    port map (
            O => \N__10464\,
            I => \frame_decoder_OFF4data_0\
        );

    \I__1212\ : LocalMux
    port map (
            O => \N__10461\,
            I => \frame_decoder_OFF4data_0\
        );

    \I__1211\ : Odrv4
    port map (
            O => \N__10458\,
            I => \frame_decoder_OFF4data_0\
        );

    \I__1210\ : CascadeMux
    port map (
            O => \N__10449\,
            I => \N__10446\
        );

    \I__1209\ : InMux
    port map (
            O => \N__10446\,
            I => \N__10443\
        );

    \I__1208\ : LocalMux
    port map (
            O => \N__10443\,
            I => \scaler_4.un2_source_data_0_cry_1_c_RNO_2\
        );

    \I__1207\ : InMux
    port map (
            O => \N__10440\,
            I => \N__10435\
        );

    \I__1206\ : CascadeMux
    port map (
            O => \N__10439\,
            I => \N__10432\
        );

    \I__1205\ : InMux
    port map (
            O => \N__10438\,
            I => \N__10428\
        );

    \I__1204\ : LocalMux
    port map (
            O => \N__10435\,
            I => \N__10425\
        );

    \I__1203\ : InMux
    port map (
            O => \N__10432\,
            I => \N__10420\
        );

    \I__1202\ : InMux
    port map (
            O => \N__10431\,
            I => \N__10420\
        );

    \I__1201\ : LocalMux
    port map (
            O => \N__10428\,
            I => \scaler_4.un2_source_data_0\
        );

    \I__1200\ : Odrv4
    port map (
            O => \N__10425\,
            I => \scaler_4.un2_source_data_0\
        );

    \I__1199\ : LocalMux
    port map (
            O => \N__10420\,
            I => \scaler_4.un2_source_data_0\
        );

    \I__1198\ : InMux
    port map (
            O => \N__10413\,
            I => \scaler_4.un2_source_data_0_cry_1\
        );

    \I__1197\ : InMux
    port map (
            O => \N__10410\,
            I => \N__10407\
        );

    \I__1196\ : LocalMux
    port map (
            O => \N__10407\,
            I => \N__10404\
        );

    \I__1195\ : Odrv4
    port map (
            O => \N__10404\,
            I => \frame_decoder_CH1data_1\
        );

    \I__1194\ : CascadeMux
    port map (
            O => \N__10401\,
            I => \N__10398\
        );

    \I__1193\ : InMux
    port map (
            O => \N__10398\,
            I => \N__10395\
        );

    \I__1192\ : LocalMux
    port map (
            O => \N__10395\,
            I => \frame_decoder_OFF1data_1\
        );

    \I__1191\ : InMux
    port map (
            O => \N__10392\,
            I => \scaler_1.un3_source_data_0_cry_0\
        );

    \I__1190\ : InMux
    port map (
            O => \N__10389\,
            I => \N__10386\
        );

    \I__1189\ : LocalMux
    port map (
            O => \N__10386\,
            I => \N__10383\
        );

    \I__1188\ : Odrv4
    port map (
            O => \N__10383\,
            I => \frame_decoder_CH1data_2\
        );

    \I__1187\ : CascadeMux
    port map (
            O => \N__10380\,
            I => \N__10377\
        );

    \I__1186\ : InMux
    port map (
            O => \N__10377\,
            I => \N__10374\
        );

    \I__1185\ : LocalMux
    port map (
            O => \N__10374\,
            I => \frame_decoder_OFF1data_2\
        );

    \I__1184\ : InMux
    port map (
            O => \N__10371\,
            I => \scaler_1.un3_source_data_0_cry_1\
        );

    \I__1183\ : InMux
    port map (
            O => \N__10368\,
            I => \N__10365\
        );

    \I__1182\ : LocalMux
    port map (
            O => \N__10365\,
            I => \N__10362\
        );

    \I__1181\ : Odrv4
    port map (
            O => \N__10362\,
            I => \frame_decoder_CH1data_3\
        );

    \I__1180\ : CascadeMux
    port map (
            O => \N__10359\,
            I => \N__10356\
        );

    \I__1179\ : InMux
    port map (
            O => \N__10356\,
            I => \N__10353\
        );

    \I__1178\ : LocalMux
    port map (
            O => \N__10353\,
            I => \frame_decoder_OFF1data_3\
        );

    \I__1177\ : InMux
    port map (
            O => \N__10350\,
            I => \scaler_1.un3_source_data_0_cry_2\
        );

    \I__1176\ : CascadeMux
    port map (
            O => \N__10347\,
            I => \N__10344\
        );

    \I__1175\ : InMux
    port map (
            O => \N__10344\,
            I => \N__10341\
        );

    \I__1174\ : LocalMux
    port map (
            O => \N__10341\,
            I => \frame_decoder_OFF1data_4\
        );

    \I__1173\ : InMux
    port map (
            O => \N__10338\,
            I => \scaler_1.un3_source_data_0_cry_3\
        );

    \I__1172\ : InMux
    port map (
            O => \N__10335\,
            I => \N__10332\
        );

    \I__1171\ : LocalMux
    port map (
            O => \N__10332\,
            I => \N__10329\
        );

    \I__1170\ : Odrv4
    port map (
            O => \N__10329\,
            I => \frame_decoder_CH1data_5\
        );

    \I__1169\ : CascadeMux
    port map (
            O => \N__10326\,
            I => \N__10323\
        );

    \I__1168\ : InMux
    port map (
            O => \N__10323\,
            I => \N__10320\
        );

    \I__1167\ : LocalMux
    port map (
            O => \N__10320\,
            I => \frame_decoder_OFF1data_5\
        );

    \I__1166\ : InMux
    port map (
            O => \N__10317\,
            I => \scaler_1.un3_source_data_0_cry_4\
        );

    \I__1165\ : InMux
    port map (
            O => \N__10314\,
            I => \N__10311\
        );

    \I__1164\ : LocalMux
    port map (
            O => \N__10311\,
            I => \frame_decoder_CH3data_1\
        );

    \I__1163\ : InMux
    port map (
            O => \N__10308\,
            I => \N__10305\
        );

    \I__1162\ : LocalMux
    port map (
            O => \N__10305\,
            I => \frame_decoder_CH3data_2\
        );

    \I__1161\ : InMux
    port map (
            O => \N__10302\,
            I => \N__10299\
        );

    \I__1160\ : LocalMux
    port map (
            O => \N__10299\,
            I => \frame_decoder_CH3data_3\
        );

    \I__1159\ : InMux
    port map (
            O => \N__10296\,
            I => \N__10293\
        );

    \I__1158\ : LocalMux
    port map (
            O => \N__10293\,
            I => \frame_decoder_CH3data_4\
        );

    \I__1157\ : InMux
    port map (
            O => \N__10290\,
            I => \N__10287\
        );

    \I__1156\ : LocalMux
    port map (
            O => \N__10287\,
            I => \frame_decoder_CH3data_5\
        );

    \I__1155\ : InMux
    port map (
            O => \N__10284\,
            I => \N__10281\
        );

    \I__1154\ : LocalMux
    port map (
            O => \N__10281\,
            I => \frame_decoder_CH3data_6\
        );

    \I__1153\ : InMux
    port map (
            O => \N__10278\,
            I => \N__10274\
        );

    \I__1152\ : InMux
    port map (
            O => \N__10277\,
            I => \N__10271\
        );

    \I__1151\ : LocalMux
    port map (
            O => \N__10274\,
            I => \frame_decoder_CH3data_7\
        );

    \I__1150\ : LocalMux
    port map (
            O => \N__10271\,
            I => \frame_decoder_CH3data_7\
        );

    \I__1149\ : InMux
    port map (
            O => \N__10266\,
            I => \N__10260\
        );

    \I__1148\ : InMux
    port map (
            O => \N__10265\,
            I => \N__10260\
        );

    \I__1147\ : LocalMux
    port map (
            O => \N__10260\,
            I => \frame_decoder_CH2data_7\
        );

    \I__1146\ : CascadeMux
    port map (
            O => \N__10257\,
            I => \N__10254\
        );

    \I__1145\ : InMux
    port map (
            O => \N__10254\,
            I => \N__10248\
        );

    \I__1144\ : InMux
    port map (
            O => \N__10253\,
            I => \N__10248\
        );

    \I__1143\ : LocalMux
    port map (
            O => \N__10248\,
            I => \N__10245\
        );

    \I__1142\ : Odrv4
    port map (
            O => \N__10245\,
            I => \frame_decoder_OFF2data_7\
        );

    \I__1141\ : InMux
    port map (
            O => \N__10242\,
            I => \N__10239\
        );

    \I__1140\ : LocalMux
    port map (
            O => \N__10239\,
            I => \scaler_2.N_783_i_l_ofxZ0\
        );

    \I__1139\ : InMux
    port map (
            O => \N__10236\,
            I => \N__10232\
        );

    \I__1138\ : InMux
    port map (
            O => \N__10235\,
            I => \N__10229\
        );

    \I__1137\ : LocalMux
    port map (
            O => \N__10232\,
            I => \N__10226\
        );

    \I__1136\ : LocalMux
    port map (
            O => \N__10229\,
            I => \uart_frame_decoder.source_CH2data_1_sqmuxa\
        );

    \I__1135\ : Odrv12
    port map (
            O => \N__10226\,
            I => \uart_frame_decoder.source_CH2data_1_sqmuxa\
        );

    \I__1134\ : CEMux
    port map (
            O => \N__10221\,
            I => \N__10218\
        );

    \I__1133\ : LocalMux
    port map (
            O => \N__10218\,
            I => \N__10215\
        );

    \I__1132\ : Span4Mux_s3_h
    port map (
            O => \N__10215\,
            I => \N__10212\
        );

    \I__1131\ : Odrv4
    port map (
            O => \N__10212\,
            I => \uart_frame_decoder.source_CH2data_1_sqmuxa_0\
        );

    \I__1130\ : CascadeMux
    port map (
            O => \N__10209\,
            I => \uart_frame_decoder.source_CH4data_1_sqmuxa_cascade_\
        );

    \I__1129\ : InMux
    port map (
            O => \N__10206\,
            I => \N__10203\
        );

    \I__1128\ : LocalMux
    port map (
            O => \N__10203\,
            I => \N__10199\
        );

    \I__1127\ : InMux
    port map (
            O => \N__10202\,
            I => \N__10196\
        );

    \I__1126\ : Odrv4
    port map (
            O => \N__10199\,
            I => \frame_decoder_OFF3data_7\
        );

    \I__1125\ : LocalMux
    port map (
            O => \N__10196\,
            I => \frame_decoder_OFF3data_7\
        );

    \I__1124\ : InMux
    port map (
            O => \N__10191\,
            I => \N__10188\
        );

    \I__1123\ : LocalMux
    port map (
            O => \N__10188\,
            I => \scaler_3.un3_source_data_0_axb_7\
        );

    \I__1122\ : CascadeMux
    port map (
            O => \N__10185\,
            I => \uart_frame_decoder.source_offset3data_1_sqmuxa_cascade_\
        );

    \I__1121\ : CascadeMux
    port map (
            O => \N__10182\,
            I => \N__10179\
        );

    \I__1120\ : InMux
    port map (
            O => \N__10179\,
            I => \N__10176\
        );

    \I__1119\ : LocalMux
    port map (
            O => \N__10176\,
            I => \frame_decoder_OFF2data_4\
        );

    \I__1118\ : InMux
    port map (
            O => \N__10173\,
            I => \scaler_2.un3_source_data_0_cry_3\
        );

    \I__1117\ : InMux
    port map (
            O => \N__10170\,
            I => \N__10167\
        );

    \I__1116\ : LocalMux
    port map (
            O => \N__10167\,
            I => \frame_decoder_CH2data_5\
        );

    \I__1115\ : CascadeMux
    port map (
            O => \N__10164\,
            I => \N__10161\
        );

    \I__1114\ : InMux
    port map (
            O => \N__10161\,
            I => \N__10158\
        );

    \I__1113\ : LocalMux
    port map (
            O => \N__10158\,
            I => \frame_decoder_OFF2data_5\
        );

    \I__1112\ : InMux
    port map (
            O => \N__10155\,
            I => \scaler_2.un3_source_data_0_cry_4\
        );

    \I__1111\ : InMux
    port map (
            O => \N__10152\,
            I => \N__10149\
        );

    \I__1110\ : LocalMux
    port map (
            O => \N__10149\,
            I => \frame_decoder_CH2data_6\
        );

    \I__1109\ : CascadeMux
    port map (
            O => \N__10146\,
            I => \N__10143\
        );

    \I__1108\ : InMux
    port map (
            O => \N__10143\,
            I => \N__10140\
        );

    \I__1107\ : LocalMux
    port map (
            O => \N__10140\,
            I => \frame_decoder_OFF2data_6\
        );

    \I__1106\ : InMux
    port map (
            O => \N__10137\,
            I => \scaler_2.un3_source_data_0_cry_5\
        );

    \I__1105\ : InMux
    port map (
            O => \N__10134\,
            I => \scaler_2.un3_source_data_0_cry_6\
        );

    \I__1104\ : InMux
    port map (
            O => \N__10131\,
            I => \bfn_2_22_0_\
        );

    \I__1103\ : InMux
    port map (
            O => \N__10128\,
            I => \scaler_2.un3_source_data_0_cry_8\
        );

    \I__1102\ : InMux
    port map (
            O => \N__10125\,
            I => \N__10122\
        );

    \I__1101\ : LocalMux
    port map (
            O => \N__10122\,
            I => \scaler_2.un3_source_data_0_axb_7\
        );

    \I__1100\ : InMux
    port map (
            O => \N__10119\,
            I => \N__10115\
        );

    \I__1099\ : InMux
    port map (
            O => \N__10118\,
            I => \N__10112\
        );

    \I__1098\ : LocalMux
    port map (
            O => \N__10115\,
            I => \N__10109\
        );

    \I__1097\ : LocalMux
    port map (
            O => \N__10112\,
            I => \uart_frame_decoder.source_CH1data_1_sqmuxa\
        );

    \I__1096\ : Odrv12
    port map (
            O => \N__10109\,
            I => \uart_frame_decoder.source_CH1data_1_sqmuxa\
        );

    \I__1095\ : CEMux
    port map (
            O => \N__10104\,
            I => \N__10101\
        );

    \I__1094\ : LocalMux
    port map (
            O => \N__10101\,
            I => \N__10098\
        );

    \I__1093\ : Odrv4
    port map (
            O => \N__10098\,
            I => \uart_frame_decoder.source_offset2data_1_sqmuxa_0\
        );

    \I__1092\ : InMux
    port map (
            O => \N__10095\,
            I => \N__10092\
        );

    \I__1091\ : LocalMux
    port map (
            O => \N__10092\,
            I => \frame_decoder_CH2data_1\
        );

    \I__1090\ : CascadeMux
    port map (
            O => \N__10089\,
            I => \N__10086\
        );

    \I__1089\ : InMux
    port map (
            O => \N__10086\,
            I => \N__10083\
        );

    \I__1088\ : LocalMux
    port map (
            O => \N__10083\,
            I => \frame_decoder_OFF2data_1\
        );

    \I__1087\ : InMux
    port map (
            O => \N__10080\,
            I => \scaler_2.un3_source_data_0_cry_0\
        );

    \I__1086\ : InMux
    port map (
            O => \N__10077\,
            I => \N__10074\
        );

    \I__1085\ : LocalMux
    port map (
            O => \N__10074\,
            I => \frame_decoder_CH2data_2\
        );

    \I__1084\ : CascadeMux
    port map (
            O => \N__10071\,
            I => \N__10068\
        );

    \I__1083\ : InMux
    port map (
            O => \N__10068\,
            I => \N__10065\
        );

    \I__1082\ : LocalMux
    port map (
            O => \N__10065\,
            I => \N__10062\
        );

    \I__1081\ : Odrv4
    port map (
            O => \N__10062\,
            I => \frame_decoder_OFF2data_2\
        );

    \I__1080\ : InMux
    port map (
            O => \N__10059\,
            I => \scaler_2.un3_source_data_0_cry_1\
        );

    \I__1079\ : InMux
    port map (
            O => \N__10056\,
            I => \N__10053\
        );

    \I__1078\ : LocalMux
    port map (
            O => \N__10053\,
            I => \frame_decoder_CH2data_3\
        );

    \I__1077\ : CascadeMux
    port map (
            O => \N__10050\,
            I => \N__10047\
        );

    \I__1076\ : InMux
    port map (
            O => \N__10047\,
            I => \N__10044\
        );

    \I__1075\ : LocalMux
    port map (
            O => \N__10044\,
            I => \frame_decoder_OFF2data_3\
        );

    \I__1074\ : InMux
    port map (
            O => \N__10041\,
            I => \scaler_2.un3_source_data_0_cry_2\
        );

    \I__1073\ : InMux
    port map (
            O => \N__10038\,
            I => \N__10035\
        );

    \I__1072\ : LocalMux
    port map (
            O => \N__10035\,
            I => \frame_decoder_CH2data_4\
        );

    \I__1071\ : InMux
    port map (
            O => \N__10032\,
            I => \N__10028\
        );

    \I__1070\ : InMux
    port map (
            O => \N__10031\,
            I => \N__10025\
        );

    \I__1069\ : LocalMux
    port map (
            O => \N__10028\,
            I => \uart_frame_decoder.state_1Z0Z_2\
        );

    \I__1068\ : LocalMux
    port map (
            O => \N__10025\,
            I => \uart_frame_decoder.state_1Z0Z_2\
        );

    \I__1067\ : InMux
    port map (
            O => \N__10020\,
            I => \N__10017\
        );

    \I__1066\ : LocalMux
    port map (
            O => \N__10017\,
            I => \N__10013\
        );

    \I__1065\ : InMux
    port map (
            O => \N__10016\,
            I => \N__10010\
        );

    \I__1064\ : Span4Mux_v
    port map (
            O => \N__10013\,
            I => \N__10007\
        );

    \I__1063\ : LocalMux
    port map (
            O => \N__10010\,
            I => \uart_frame_decoder.state_1Z0Z_4\
        );

    \I__1062\ : Odrv4
    port map (
            O => \N__10007\,
            I => \uart_frame_decoder.state_1Z0Z_4\
        );

    \I__1061\ : CascadeMux
    port map (
            O => \N__10002\,
            I => \N__9998\
        );

    \I__1060\ : InMux
    port map (
            O => \N__10001\,
            I => \N__9994\
        );

    \I__1059\ : InMux
    port map (
            O => \N__9998\,
            I => \N__9989\
        );

    \I__1058\ : InMux
    port map (
            O => \N__9997\,
            I => \N__9989\
        );

    \I__1057\ : LocalMux
    port map (
            O => \N__9994\,
            I => \uart_frame_decoder.countZ0Z_2\
        );

    \I__1056\ : LocalMux
    port map (
            O => \N__9989\,
            I => \uart_frame_decoder.countZ0Z_2\
        );

    \I__1055\ : InMux
    port map (
            O => \N__9984\,
            I => \N__9978\
        );

    \I__1054\ : InMux
    port map (
            O => \N__9983\,
            I => \N__9971\
        );

    \I__1053\ : InMux
    port map (
            O => \N__9982\,
            I => \N__9971\
        );

    \I__1052\ : InMux
    port map (
            O => \N__9981\,
            I => \N__9971\
        );

    \I__1051\ : LocalMux
    port map (
            O => \N__9978\,
            I => \uart_frame_decoder.countZ0Z_1\
        );

    \I__1050\ : LocalMux
    port map (
            O => \N__9971\,
            I => \uart_frame_decoder.countZ0Z_1\
        );

    \I__1049\ : CascadeMux
    port map (
            O => \N__9966\,
            I => \N__9962\
        );

    \I__1048\ : InMux
    port map (
            O => \N__9965\,
            I => \N__9957\
        );

    \I__1047\ : InMux
    port map (
            O => \N__9962\,
            I => \N__9954\
        );

    \I__1046\ : InMux
    port map (
            O => \N__9961\,
            I => \N__9949\
        );

    \I__1045\ : InMux
    port map (
            O => \N__9960\,
            I => \N__9949\
        );

    \I__1044\ : LocalMux
    port map (
            O => \N__9957\,
            I => \uart_frame_decoder.count8_0\
        );

    \I__1043\ : LocalMux
    port map (
            O => \N__9954\,
            I => \uart_frame_decoder.count8_0\
        );

    \I__1042\ : LocalMux
    port map (
            O => \N__9949\,
            I => \uart_frame_decoder.count8_0\
        );

    \I__1041\ : CascadeMux
    port map (
            O => \N__9942\,
            I => \uart_frame_decoder.state_1_ns_i_i_0_0_cascade_\
        );

    \I__1040\ : InMux
    port map (
            O => \N__9939\,
            I => \N__9934\
        );

    \I__1039\ : InMux
    port map (
            O => \N__9938\,
            I => \N__9929\
        );

    \I__1038\ : InMux
    port map (
            O => \N__9937\,
            I => \N__9929\
        );

    \I__1037\ : LocalMux
    port map (
            O => \N__9934\,
            I => \uart_frame_decoder.WDTZ0Z_11\
        );

    \I__1036\ : LocalMux
    port map (
            O => \N__9929\,
            I => \uart_frame_decoder.WDTZ0Z_11\
        );

    \I__1035\ : InMux
    port map (
            O => \N__9924\,
            I => \N__9920\
        );

    \I__1034\ : InMux
    port map (
            O => \N__9923\,
            I => \N__9917\
        );

    \I__1033\ : LocalMux
    port map (
            O => \N__9920\,
            I => \uart_frame_decoder.WDTZ0Z_10\
        );

    \I__1032\ : LocalMux
    port map (
            O => \N__9917\,
            I => \uart_frame_decoder.WDTZ0Z_10\
        );

    \I__1031\ : CascadeMux
    port map (
            O => \N__9912\,
            I => \N__9908\
        );

    \I__1030\ : InMux
    port map (
            O => \N__9911\,
            I => \N__9905\
        );

    \I__1029\ : InMux
    port map (
            O => \N__9908\,
            I => \N__9902\
        );

    \I__1028\ : LocalMux
    port map (
            O => \N__9905\,
            I => \uart_frame_decoder.WDTZ0Z_13\
        );

    \I__1027\ : LocalMux
    port map (
            O => \N__9902\,
            I => \uart_frame_decoder.WDTZ0Z_13\
        );

    \I__1026\ : InMux
    port map (
            O => \N__9897\,
            I => \N__9892\
        );

    \I__1025\ : InMux
    port map (
            O => \N__9896\,
            I => \N__9887\
        );

    \I__1024\ : InMux
    port map (
            O => \N__9895\,
            I => \N__9887\
        );

    \I__1023\ : LocalMux
    port map (
            O => \N__9892\,
            I => \uart_frame_decoder.WDTZ0Z_12\
        );

    \I__1022\ : LocalMux
    port map (
            O => \N__9887\,
            I => \uart_frame_decoder.WDTZ0Z_12\
        );

    \I__1021\ : InMux
    port map (
            O => \N__9882\,
            I => \N__9878\
        );

    \I__1020\ : InMux
    port map (
            O => \N__9881\,
            I => \N__9875\
        );

    \I__1019\ : LocalMux
    port map (
            O => \N__9878\,
            I => \uart_frame_decoder.WDTZ0Z_9\
        );

    \I__1018\ : LocalMux
    port map (
            O => \N__9875\,
            I => \uart_frame_decoder.WDTZ0Z_9\
        );

    \I__1017\ : CascadeMux
    port map (
            O => \N__9870\,
            I => \uart_frame_decoder.WDT_RNIAGPBZ0Z_10_cascade_\
        );

    \I__1016\ : InMux
    port map (
            O => \N__9867\,
            I => \N__9864\
        );

    \I__1015\ : LocalMux
    port map (
            O => \N__9864\,
            I => \uart_frame_decoder.WDT8lto13_1\
        );

    \I__1014\ : CascadeMux
    port map (
            O => \N__9861\,
            I => \uart_frame_decoder.WDT8lt14_0_cascade_\
        );

    \I__1013\ : CascadeMux
    port map (
            O => \N__9858\,
            I => \N__9854\
        );

    \I__1012\ : InMux
    port map (
            O => \N__9857\,
            I => \N__9851\
        );

    \I__1011\ : InMux
    port map (
            O => \N__9854\,
            I => \N__9848\
        );

    \I__1010\ : LocalMux
    port map (
            O => \N__9851\,
            I => \uart_frame_decoder.WDT8_0_i\
        );

    \I__1009\ : LocalMux
    port map (
            O => \N__9848\,
            I => \uart_frame_decoder.WDT8_0_i\
        );

    \I__1008\ : InMux
    port map (
            O => \N__9843\,
            I => \N__9839\
        );

    \I__1007\ : InMux
    port map (
            O => \N__9842\,
            I => \N__9836\
        );

    \I__1006\ : LocalMux
    port map (
            O => \N__9839\,
            I => \uart_frame_decoder.WDTZ0Z_6\
        );

    \I__1005\ : LocalMux
    port map (
            O => \N__9836\,
            I => \uart_frame_decoder.WDTZ0Z_6\
        );

    \I__1004\ : InMux
    port map (
            O => \N__9831\,
            I => \N__9827\
        );

    \I__1003\ : InMux
    port map (
            O => \N__9830\,
            I => \N__9824\
        );

    \I__1002\ : LocalMux
    port map (
            O => \N__9827\,
            I => \uart_frame_decoder.WDTZ0Z_5\
        );

    \I__1001\ : LocalMux
    port map (
            O => \N__9824\,
            I => \uart_frame_decoder.WDTZ0Z_5\
        );

    \I__1000\ : CascadeMux
    port map (
            O => \N__9819\,
            I => \N__9815\
        );

    \I__999\ : InMux
    port map (
            O => \N__9818\,
            I => \N__9812\
        );

    \I__998\ : InMux
    port map (
            O => \N__9815\,
            I => \N__9809\
        );

    \I__997\ : LocalMux
    port map (
            O => \N__9812\,
            I => \uart_frame_decoder.WDTZ0Z_7\
        );

    \I__996\ : LocalMux
    port map (
            O => \N__9809\,
            I => \uart_frame_decoder.WDTZ0Z_7\
        );

    \I__995\ : InMux
    port map (
            O => \N__9804\,
            I => \N__9800\
        );

    \I__994\ : InMux
    port map (
            O => \N__9803\,
            I => \N__9797\
        );

    \I__993\ : LocalMux
    port map (
            O => \N__9800\,
            I => \uart_frame_decoder.WDTZ0Z_4\
        );

    \I__992\ : LocalMux
    port map (
            O => \N__9797\,
            I => \uart_frame_decoder.WDTZ0Z_4\
        );

    \I__991\ : InMux
    port map (
            O => \N__9792\,
            I => \N__9789\
        );

    \I__990\ : LocalMux
    port map (
            O => \N__9789\,
            I => \uart_frame_decoder.WDT_RNIM6B11Z0Z_4\
        );

    \I__989\ : InMux
    port map (
            O => \N__9786\,
            I => \N__9781\
        );

    \I__988\ : InMux
    port map (
            O => \N__9785\,
            I => \N__9778\
        );

    \I__987\ : InMux
    port map (
            O => \N__9784\,
            I => \N__9775\
        );

    \I__986\ : LocalMux
    port map (
            O => \N__9781\,
            I => \uart_frame_decoder.WDTZ0Z_15\
        );

    \I__985\ : LocalMux
    port map (
            O => \N__9778\,
            I => \uart_frame_decoder.WDTZ0Z_15\
        );

    \I__984\ : LocalMux
    port map (
            O => \N__9775\,
            I => \uart_frame_decoder.WDTZ0Z_15\
        );

    \I__983\ : CascadeMux
    port map (
            O => \N__9768\,
            I => \N__9764\
        );

    \I__982\ : InMux
    port map (
            O => \N__9767\,
            I => \N__9760\
        );

    \I__981\ : InMux
    port map (
            O => \N__9764\,
            I => \N__9757\
        );

    \I__980\ : InMux
    port map (
            O => \N__9763\,
            I => \N__9754\
        );

    \I__979\ : LocalMux
    port map (
            O => \N__9760\,
            I => \uart_frame_decoder.WDTZ0Z_14\
        );

    \I__978\ : LocalMux
    port map (
            O => \N__9757\,
            I => \uart_frame_decoder.WDTZ0Z_14\
        );

    \I__977\ : LocalMux
    port map (
            O => \N__9754\,
            I => \uart_frame_decoder.WDTZ0Z_14\
        );

    \I__976\ : InMux
    port map (
            O => \N__9747\,
            I => \N__9744\
        );

    \I__975\ : LocalMux
    port map (
            O => \N__9744\,
            I => \uart_frame_decoder.WDT8lt14_0\
        );

    \I__974\ : CascadeMux
    port map (
            O => \N__9741\,
            I => \uart_frame_decoder.WDT_RNIJUEI2Z0Z_15_cascade_\
        );

    \I__973\ : InMux
    port map (
            O => \N__9738\,
            I => \N__9732\
        );

    \I__972\ : InMux
    port map (
            O => \N__9737\,
            I => \N__9732\
        );

    \I__971\ : LocalMux
    port map (
            O => \N__9732\,
            I => \uart_frame_decoder.state_1Z0Z_3\
        );

    \I__970\ : InMux
    port map (
            O => \N__9729\,
            I => \N__9726\
        );

    \I__969\ : LocalMux
    port map (
            O => \N__9726\,
            I => \N__9723\
        );

    \I__968\ : Span4Mux_s3_v
    port map (
            O => \N__9723\,
            I => \N__9720\
        );

    \I__967\ : Odrv4
    port map (
            O => \N__9720\,
            I => \scaler_4.un3_source_data_0_axb_7\
        );

    \I__966\ : InMux
    port map (
            O => \N__9717\,
            I => \scaler_4.un3_source_data_0_cry_6\
        );

    \I__965\ : InMux
    port map (
            O => \N__9714\,
            I => \bfn_1_30_0_\
        );

    \I__964\ : InMux
    port map (
            O => \N__9711\,
            I => \scaler_4.un3_source_data_0_cry_8\
        );

    \I__963\ : InMux
    port map (
            O => \N__9708\,
            I => \N__9704\
        );

    \I__962\ : InMux
    port map (
            O => \N__9707\,
            I => \N__9701\
        );

    \I__961\ : LocalMux
    port map (
            O => \N__9704\,
            I => \N__9696\
        );

    \I__960\ : LocalMux
    port map (
            O => \N__9701\,
            I => \N__9696\
        );

    \I__959\ : Odrv12
    port map (
            O => \N__9696\,
            I => \frame_decoder_OFF4data_7\
        );

    \I__958\ : InMux
    port map (
            O => \N__9693\,
            I => \N__9690\
        );

    \I__957\ : LocalMux
    port map (
            O => \N__9690\,
            I => \scaler_4.N_807_i_l_ofxZ0\
        );

    \I__956\ : InMux
    port map (
            O => \N__9687\,
            I => \N__9683\
        );

    \I__955\ : InMux
    port map (
            O => \N__9686\,
            I => \N__9680\
        );

    \I__954\ : LocalMux
    port map (
            O => \N__9683\,
            I => \uart_frame_decoder.WDTZ0Z_8\
        );

    \I__953\ : LocalMux
    port map (
            O => \N__9680\,
            I => \uart_frame_decoder.WDTZ0Z_8\
        );

    \I__952\ : InMux
    port map (
            O => \N__9675\,
            I => \N__9672\
        );

    \I__951\ : LocalMux
    port map (
            O => \N__9672\,
            I => \frame_decoder_CH4data_1\
        );

    \I__950\ : CascadeMux
    port map (
            O => \N__9669\,
            I => \N__9666\
        );

    \I__949\ : InMux
    port map (
            O => \N__9666\,
            I => \N__9663\
        );

    \I__948\ : LocalMux
    port map (
            O => \N__9663\,
            I => \N__9660\
        );

    \I__947\ : Odrv4
    port map (
            O => \N__9660\,
            I => \frame_decoder_OFF4data_1\
        );

    \I__946\ : InMux
    port map (
            O => \N__9657\,
            I => \scaler_4.un3_source_data_0_cry_0\
        );

    \I__945\ : InMux
    port map (
            O => \N__9654\,
            I => \N__9651\
        );

    \I__944\ : LocalMux
    port map (
            O => \N__9651\,
            I => \frame_decoder_CH4data_2\
        );

    \I__943\ : CascadeMux
    port map (
            O => \N__9648\,
            I => \N__9645\
        );

    \I__942\ : InMux
    port map (
            O => \N__9645\,
            I => \N__9642\
        );

    \I__941\ : LocalMux
    port map (
            O => \N__9642\,
            I => \N__9639\
        );

    \I__940\ : Odrv4
    port map (
            O => \N__9639\,
            I => \frame_decoder_OFF4data_2\
        );

    \I__939\ : InMux
    port map (
            O => \N__9636\,
            I => \scaler_4.un3_source_data_0_cry_1\
        );

    \I__938\ : InMux
    port map (
            O => \N__9633\,
            I => \N__9630\
        );

    \I__937\ : LocalMux
    port map (
            O => \N__9630\,
            I => \frame_decoder_CH4data_3\
        );

    \I__936\ : CascadeMux
    port map (
            O => \N__9627\,
            I => \N__9624\
        );

    \I__935\ : InMux
    port map (
            O => \N__9624\,
            I => \N__9621\
        );

    \I__934\ : LocalMux
    port map (
            O => \N__9621\,
            I => \N__9618\
        );

    \I__933\ : Odrv4
    port map (
            O => \N__9618\,
            I => \frame_decoder_OFF4data_3\
        );

    \I__932\ : InMux
    port map (
            O => \N__9615\,
            I => \scaler_4.un3_source_data_0_cry_2\
        );

    \I__931\ : InMux
    port map (
            O => \N__9612\,
            I => \N__9609\
        );

    \I__930\ : LocalMux
    port map (
            O => \N__9609\,
            I => \frame_decoder_CH4data_4\
        );

    \I__929\ : CascadeMux
    port map (
            O => \N__9606\,
            I => \N__9603\
        );

    \I__928\ : InMux
    port map (
            O => \N__9603\,
            I => \N__9600\
        );

    \I__927\ : LocalMux
    port map (
            O => \N__9600\,
            I => \N__9597\
        );

    \I__926\ : Odrv4
    port map (
            O => \N__9597\,
            I => \frame_decoder_OFF4data_4\
        );

    \I__925\ : InMux
    port map (
            O => \N__9594\,
            I => \scaler_4.un3_source_data_0_cry_3\
        );

    \I__924\ : InMux
    port map (
            O => \N__9591\,
            I => \N__9588\
        );

    \I__923\ : LocalMux
    port map (
            O => \N__9588\,
            I => \N__9585\
        );

    \I__922\ : Odrv4
    port map (
            O => \N__9585\,
            I => \frame_decoder_OFF4data_5\
        );

    \I__921\ : CascadeMux
    port map (
            O => \N__9582\,
            I => \N__9579\
        );

    \I__920\ : InMux
    port map (
            O => \N__9579\,
            I => \N__9576\
        );

    \I__919\ : LocalMux
    port map (
            O => \N__9576\,
            I => \frame_decoder_CH4data_5\
        );

    \I__918\ : InMux
    port map (
            O => \N__9573\,
            I => \scaler_4.un3_source_data_0_cry_4\
        );

    \I__917\ : InMux
    port map (
            O => \N__9570\,
            I => \N__9567\
        );

    \I__916\ : LocalMux
    port map (
            O => \N__9567\,
            I => \frame_decoder_CH4data_6\
        );

    \I__915\ : CascadeMux
    port map (
            O => \N__9564\,
            I => \N__9561\
        );

    \I__914\ : InMux
    port map (
            O => \N__9561\,
            I => \N__9558\
        );

    \I__913\ : LocalMux
    port map (
            O => \N__9558\,
            I => \N__9555\
        );

    \I__912\ : Odrv4
    port map (
            O => \N__9555\,
            I => \frame_decoder_OFF4data_6\
        );

    \I__911\ : InMux
    port map (
            O => \N__9552\,
            I => \scaler_4.un3_source_data_0_cry_5\
        );

    \I__910\ : CEMux
    port map (
            O => \N__9549\,
            I => \N__9546\
        );

    \I__909\ : LocalMux
    port map (
            O => \N__9546\,
            I => \N__9543\
        );

    \I__908\ : Span4Mux_v
    port map (
            O => \N__9543\,
            I => \N__9540\
        );

    \I__907\ : Odrv4
    port map (
            O => \N__9540\,
            I => \uart_frame_decoder.source_offset4data_1_sqmuxa_0\
        );

    \I__906\ : CascadeMux
    port map (
            O => \N__9537\,
            I => \N__9534\
        );

    \I__905\ : InMux
    port map (
            O => \N__9534\,
            I => \N__9528\
        );

    \I__904\ : InMux
    port map (
            O => \N__9533\,
            I => \N__9528\
        );

    \I__903\ : LocalMux
    port map (
            O => \N__9528\,
            I => \N__9525\
        );

    \I__902\ : Odrv4
    port map (
            O => \N__9525\,
            I => \scaler_3.un3_source_data_0_cry_5_c_RNI4DBI\
        );

    \I__901\ : InMux
    port map (
            O => \N__9522\,
            I => \scaler_3.un2_source_data_0_cry_6\
        );

    \I__900\ : CascadeMux
    port map (
            O => \N__9519\,
            I => \N__9516\
        );

    \I__899\ : InMux
    port map (
            O => \N__9516\,
            I => \N__9510\
        );

    \I__898\ : InMux
    port map (
            O => \N__9515\,
            I => \N__9510\
        );

    \I__897\ : LocalMux
    port map (
            O => \N__9510\,
            I => \N__9507\
        );

    \I__896\ : Odrv4
    port map (
            O => \N__9507\,
            I => \scaler_3.un3_source_data_0_cry_6_c_RNI7HCI\
        );

    \I__895\ : InMux
    port map (
            O => \N__9504\,
            I => \scaler_3.un2_source_data_0_cry_7\
        );

    \I__894\ : InMux
    port map (
            O => \N__9501\,
            I => \N__9498\
        );

    \I__893\ : LocalMux
    port map (
            O => \N__9498\,
            I => \N__9494\
        );

    \I__892\ : InMux
    port map (
            O => \N__9497\,
            I => \N__9491\
        );

    \I__891\ : Odrv4
    port map (
            O => \N__9494\,
            I => \scaler_3.un3_source_data_0_cry_7_c_RNI8JDI\
        );

    \I__890\ : LocalMux
    port map (
            O => \N__9491\,
            I => \scaler_3.un3_source_data_0_cry_7_c_RNI8JDI\
        );

    \I__889\ : CascadeMux
    port map (
            O => \N__9486\,
            I => \N__9483\
        );

    \I__888\ : InMux
    port map (
            O => \N__9483\,
            I => \N__9480\
        );

    \I__887\ : LocalMux
    port map (
            O => \N__9480\,
            I => \N__9477\
        );

    \I__886\ : Odrv4
    port map (
            O => \N__9477\,
            I => \scaler_3.un3_source_data_0_cry_8_c_RNIRV25\
        );

    \I__885\ : InMux
    port map (
            O => \N__9474\,
            I => \bfn_1_26_0_\
        );

    \I__884\ : InMux
    port map (
            O => \N__9471\,
            I => \scaler_3.un2_source_data_0_cry_9\
        );

    \I__883\ : InMux
    port map (
            O => \N__9468\,
            I => \N__9465\
        );

    \I__882\ : LocalMux
    port map (
            O => \N__9465\,
            I => \scaler_3.N_795_i_l_ofxZ0\
        );

    \I__881\ : CascadeMux
    port map (
            O => \N__9462\,
            I => \N__9459\
        );

    \I__880\ : InMux
    port map (
            O => \N__9459\,
            I => \N__9456\
        );

    \I__879\ : LocalMux
    port map (
            O => \N__9456\,
            I => \scaler_3.un2_source_data_0_cry_1_c_RNO_1\
        );

    \I__878\ : InMux
    port map (
            O => \N__9453\,
            I => \scaler_3.un2_source_data_0_cry_1\
        );

    \I__877\ : CascadeMux
    port map (
            O => \N__9450\,
            I => \N__9447\
        );

    \I__876\ : InMux
    port map (
            O => \N__9447\,
            I => \N__9441\
        );

    \I__875\ : InMux
    port map (
            O => \N__9446\,
            I => \N__9441\
        );

    \I__874\ : LocalMux
    port map (
            O => \N__9441\,
            I => \N__9438\
        );

    \I__873\ : Odrv12
    port map (
            O => \N__9438\,
            I => \scaler_3.un3_source_data_0_cry_1_c_RNIOS6I\
        );

    \I__872\ : InMux
    port map (
            O => \N__9435\,
            I => \scaler_3.un2_source_data_0_cry_2\
        );

    \I__871\ : CascadeMux
    port map (
            O => \N__9432\,
            I => \N__9429\
        );

    \I__870\ : InMux
    port map (
            O => \N__9429\,
            I => \N__9423\
        );

    \I__869\ : InMux
    port map (
            O => \N__9428\,
            I => \N__9423\
        );

    \I__868\ : LocalMux
    port map (
            O => \N__9423\,
            I => \N__9420\
        );

    \I__867\ : Odrv4
    port map (
            O => \N__9420\,
            I => \scaler_3.un3_source_data_0_cry_2_c_RNIR08I\
        );

    \I__866\ : InMux
    port map (
            O => \N__9417\,
            I => \scaler_3.un2_source_data_0_cry_3\
        );

    \I__865\ : CascadeMux
    port map (
            O => \N__9414\,
            I => \N__9411\
        );

    \I__864\ : InMux
    port map (
            O => \N__9411\,
            I => \N__9405\
        );

    \I__863\ : InMux
    port map (
            O => \N__9410\,
            I => \N__9405\
        );

    \I__862\ : LocalMux
    port map (
            O => \N__9405\,
            I => \N__9402\
        );

    \I__861\ : Odrv4
    port map (
            O => \N__9402\,
            I => \scaler_3.un3_source_data_0_cry_3_c_RNIU49I\
        );

    \I__860\ : InMux
    port map (
            O => \N__9399\,
            I => \scaler_3.un2_source_data_0_cry_4\
        );

    \I__859\ : CascadeMux
    port map (
            O => \N__9396\,
            I => \N__9393\
        );

    \I__858\ : InMux
    port map (
            O => \N__9393\,
            I => \N__9387\
        );

    \I__857\ : InMux
    port map (
            O => \N__9392\,
            I => \N__9387\
        );

    \I__856\ : LocalMux
    port map (
            O => \N__9387\,
            I => \N__9384\
        );

    \I__855\ : Odrv4
    port map (
            O => \N__9384\,
            I => \scaler_3.un3_source_data_0_cry_4_c_RNI19AI\
        );

    \I__854\ : InMux
    port map (
            O => \N__9381\,
            I => \scaler_3.un2_source_data_0_cry_5\
        );

    \I__853\ : CascadeMux
    port map (
            O => \N__9378\,
            I => \N__9375\
        );

    \I__852\ : InMux
    port map (
            O => \N__9375\,
            I => \N__9372\
        );

    \I__851\ : LocalMux
    port map (
            O => \N__9372\,
            I => \frame_decoder_OFF3data_3\
        );

    \I__850\ : InMux
    port map (
            O => \N__9369\,
            I => \scaler_3.un3_source_data_0_cry_2\
        );

    \I__849\ : CascadeMux
    port map (
            O => \N__9366\,
            I => \N__9363\
        );

    \I__848\ : InMux
    port map (
            O => \N__9363\,
            I => \N__9360\
        );

    \I__847\ : LocalMux
    port map (
            O => \N__9360\,
            I => \frame_decoder_OFF3data_4\
        );

    \I__846\ : InMux
    port map (
            O => \N__9357\,
            I => \scaler_3.un3_source_data_0_cry_3\
        );

    \I__845\ : CascadeMux
    port map (
            O => \N__9354\,
            I => \N__9351\
        );

    \I__844\ : InMux
    port map (
            O => \N__9351\,
            I => \N__9348\
        );

    \I__843\ : LocalMux
    port map (
            O => \N__9348\,
            I => \frame_decoder_OFF3data_5\
        );

    \I__842\ : InMux
    port map (
            O => \N__9345\,
            I => \scaler_3.un3_source_data_0_cry_4\
        );

    \I__841\ : CascadeMux
    port map (
            O => \N__9342\,
            I => \N__9339\
        );

    \I__840\ : InMux
    port map (
            O => \N__9339\,
            I => \N__9336\
        );

    \I__839\ : LocalMux
    port map (
            O => \N__9336\,
            I => \frame_decoder_OFF3data_6\
        );

    \I__838\ : InMux
    port map (
            O => \N__9333\,
            I => \scaler_3.un3_source_data_0_cry_5\
        );

    \I__837\ : InMux
    port map (
            O => \N__9330\,
            I => \scaler_3.un3_source_data_0_cry_6\
        );

    \I__836\ : InMux
    port map (
            O => \N__9327\,
            I => \bfn_1_24_0_\
        );

    \I__835\ : InMux
    port map (
            O => \N__9324\,
            I => \scaler_3.un3_source_data_0_cry_8\
        );

    \I__834\ : InMux
    port map (
            O => \N__9321\,
            I => \scaler_3.un3_source_data_0_cry_0\
        );

    \I__833\ : CascadeMux
    port map (
            O => \N__9318\,
            I => \N__9315\
        );

    \I__832\ : InMux
    port map (
            O => \N__9315\,
            I => \N__9312\
        );

    \I__831\ : LocalMux
    port map (
            O => \N__9312\,
            I => \frame_decoder_OFF3data_2\
        );

    \I__830\ : InMux
    port map (
            O => \N__9309\,
            I => \scaler_3.un3_source_data_0_cry_1\
        );

    \I__829\ : InMux
    port map (
            O => \N__9306\,
            I => \N__9302\
        );

    \I__828\ : InMux
    port map (
            O => \N__9305\,
            I => \N__9299\
        );

    \I__827\ : LocalMux
    port map (
            O => \N__9302\,
            I => \uart_frame_decoder.count8_0_i\
        );

    \I__826\ : LocalMux
    port map (
            O => \N__9299\,
            I => \uart_frame_decoder.count8_0_i\
        );

    \I__825\ : InMux
    port map (
            O => \N__9294\,
            I => \N__9291\
        );

    \I__824\ : LocalMux
    port map (
            O => \N__9291\,
            I => \uart_frame_decoder.count_i_2\
        );

    \I__823\ : InMux
    port map (
            O => \N__9288\,
            I => \uart_frame_decoder.count8\
        );

    \I__822\ : InMux
    port map (
            O => \N__9285\,
            I => \N__9279\
        );

    \I__821\ : InMux
    port map (
            O => \N__9284\,
            I => \N__9279\
        );

    \I__820\ : LocalMux
    port map (
            O => \N__9279\,
            I => \uart_frame_decoder.count8_cry_2_c_RNICKSZ0Z21\
        );

    \I__819\ : CascadeMux
    port map (
            O => \N__9276\,
            I => \uart_frame_decoder.count8_cry_2_c_RNICKSZ0Z21_cascade_\
        );

    \I__818\ : CascadeMux
    port map (
            O => \N__9273\,
            I => \N__9269\
        );

    \I__817\ : InMux
    port map (
            O => \N__9272\,
            I => \N__9264\
        );

    \I__816\ : InMux
    port map (
            O => \N__9269\,
            I => \N__9264\
        );

    \I__815\ : LocalMux
    port map (
            O => \N__9264\,
            I => \uart_frame_decoder.count_RNIV5MSZ0Z_0\
        );

    \I__814\ : SRMux
    port map (
            O => \N__9261\,
            I => \N__9258\
        );

    \I__813\ : LocalMux
    port map (
            O => \N__9258\,
            I => \N__9254\
        );

    \I__812\ : SRMux
    port map (
            O => \N__9257\,
            I => \N__9251\
        );

    \I__811\ : Span4Mux_v
    port map (
            O => \N__9254\,
            I => \N__9246\
        );

    \I__810\ : LocalMux
    port map (
            O => \N__9251\,
            I => \N__9246\
        );

    \I__809\ : Odrv4
    port map (
            O => \N__9246\,
            I => \uart_frame_decoder.source_data_valid_2_sqmuxa_iZ0\
        );

    \I__808\ : InMux
    port map (
            O => \N__9243\,
            I => \uart_frame_decoder.un1_WDT_cry_8\
        );

    \I__807\ : InMux
    port map (
            O => \N__9240\,
            I => \uart_frame_decoder.un1_WDT_cry_9\
        );

    \I__806\ : InMux
    port map (
            O => \N__9237\,
            I => \uart_frame_decoder.un1_WDT_cry_10\
        );

    \I__805\ : InMux
    port map (
            O => \N__9234\,
            I => \uart_frame_decoder.un1_WDT_cry_11\
        );

    \I__804\ : InMux
    port map (
            O => \N__9231\,
            I => \uart_frame_decoder.un1_WDT_cry_12\
        );

    \I__803\ : InMux
    port map (
            O => \N__9228\,
            I => \uart_frame_decoder.un1_WDT_cry_13\
        );

    \I__802\ : InMux
    port map (
            O => \N__9225\,
            I => \uart_frame_decoder.un1_WDT_cry_14\
        );

    \I__801\ : InMux
    port map (
            O => \N__9222\,
            I => \N__9219\
        );

    \I__800\ : LocalMux
    port map (
            O => \N__9219\,
            I => \uart_frame_decoder.count8_axb_1\
        );

    \I__799\ : InMux
    port map (
            O => \N__9216\,
            I => \N__9213\
        );

    \I__798\ : LocalMux
    port map (
            O => \N__9213\,
            I => \uart_frame_decoder.WDTZ0Z_1\
        );

    \I__797\ : InMux
    port map (
            O => \N__9210\,
            I => \uart_frame_decoder.un1_WDT_cry_0\
        );

    \I__796\ : InMux
    port map (
            O => \N__9207\,
            I => \N__9204\
        );

    \I__795\ : LocalMux
    port map (
            O => \N__9204\,
            I => \uart_frame_decoder.WDTZ0Z_2\
        );

    \I__794\ : InMux
    port map (
            O => \N__9201\,
            I => \uart_frame_decoder.un1_WDT_cry_1\
        );

    \I__793\ : InMux
    port map (
            O => \N__9198\,
            I => \N__9195\
        );

    \I__792\ : LocalMux
    port map (
            O => \N__9195\,
            I => \uart_frame_decoder.WDTZ0Z_3\
        );

    \I__791\ : InMux
    port map (
            O => \N__9192\,
            I => \uart_frame_decoder.un1_WDT_cry_2\
        );

    \I__790\ : InMux
    port map (
            O => \N__9189\,
            I => \uart_frame_decoder.un1_WDT_cry_3\
        );

    \I__789\ : InMux
    port map (
            O => \N__9186\,
            I => \uart_frame_decoder.un1_WDT_cry_4\
        );

    \I__788\ : InMux
    port map (
            O => \N__9183\,
            I => \uart_frame_decoder.un1_WDT_cry_5\
        );

    \I__787\ : InMux
    port map (
            O => \N__9180\,
            I => \uart_frame_decoder.un1_WDT_cry_6\
        );

    \I__786\ : InMux
    port map (
            O => \N__9177\,
            I => \bfn_1_18_0_\
        );

    \I__785\ : InMux
    port map (
            O => \N__9174\,
            I => \N__9171\
        );

    \I__784\ : LocalMux
    port map (
            O => \N__9171\,
            I => \uart_frame_decoder.WDTZ0Z_0\
        );

    \IN_MUX_bfv_1_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_19_0_\
        );

    \IN_MUX_bfv_5_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_15_0_\
        );

    \IN_MUX_bfv_1_29_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_29_0_\
        );

    \IN_MUX_bfv_1_30_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \scaler_4.un3_source_data_0_cry_7\,
            carryinitout => \bfn_1_30_0_\
        );

    \IN_MUX_bfv_2_29_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_29_0_\
        );

    \IN_MUX_bfv_2_30_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \scaler_4.un2_source_data_0_cry_8\,
            carryinitout => \bfn_2_30_0_\
        );

    \IN_MUX_bfv_1_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_23_0_\
        );

    \IN_MUX_bfv_1_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \scaler_3.un3_source_data_0_cry_7\,
            carryinitout => \bfn_1_24_0_\
        );

    \IN_MUX_bfv_1_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_25_0_\
        );

    \IN_MUX_bfv_1_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \scaler_3.un2_source_data_0_cry_8\,
            carryinitout => \bfn_1_26_0_\
        );

    \IN_MUX_bfv_2_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_21_0_\
        );

    \IN_MUX_bfv_2_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \scaler_2.un3_source_data_0_cry_7\,
            carryinitout => \bfn_2_22_0_\
        );

    \IN_MUX_bfv_3_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_21_0_\
        );

    \IN_MUX_bfv_3_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \scaler_2.un2_source_data_0_cry_8\,
            carryinitout => \bfn_3_22_0_\
        );

    \IN_MUX_bfv_2_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_27_0_\
        );

    \IN_MUX_bfv_2_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \scaler_1.un3_source_data_0_cry_7\,
            carryinitout => \bfn_2_28_0_\
        );

    \IN_MUX_bfv_3_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_28_0_\
        );

    \IN_MUX_bfv_3_29_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \scaler_1.un2_source_data_0_cry_8\,
            carryinitout => \bfn_3_29_0_\
        );

    \IN_MUX_bfv_5_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_17_0_\
        );

    \IN_MUX_bfv_5_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \reset_module_System.count_1_cry_8\,
            carryinitout => \bfn_5_18_0_\
        );

    \IN_MUX_bfv_5_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \reset_module_System.count_1_cry_16\,
            carryinitout => \bfn_5_19_0_\
        );

    \IN_MUX_bfv_4_29_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_29_0_\
        );

    \IN_MUX_bfv_4_30_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ppm_encoder_1.un1_throttle_cry_13\,
            carryinitout => \bfn_4_30_0_\
        );

    \IN_MUX_bfv_3_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_26_0_\
        );

    \IN_MUX_bfv_3_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ppm_encoder_1.un1_rudder_cry_13\,
            carryinitout => \bfn_3_27_0_\
        );

    \IN_MUX_bfv_4_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_27_0_\
        );

    \IN_MUX_bfv_4_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ppm_encoder_1.un1_elevator_cry_13\,
            carryinitout => \bfn_4_28_0_\
        );

    \IN_MUX_bfv_4_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_24_0_\
        );

    \IN_MUX_bfv_4_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ppm_encoder_1.un1_aileron_cry_13\,
            carryinitout => \bfn_4_25_0_\
        );

    \IN_MUX_bfv_9_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_26_0_\
        );

    \IN_MUX_bfv_9_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ppm_encoder_1.un1_init_pulses_3_cry_7\,
            carryinitout => \bfn_9_27_0_\
        );

    \IN_MUX_bfv_9_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ppm_encoder_1.un1_init_pulses_3_cry_15\,
            carryinitout => \bfn_9_28_0_\
        );

    \IN_MUX_bfv_7_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_23_0_\
        );

    \IN_MUX_bfv_7_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ppm_encoder_1.un1_init_pulses_0_cry_7\,
            carryinitout => \bfn_7_24_0_\
        );

    \IN_MUX_bfv_7_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ppm_encoder_1.un1_init_pulses_0_cry_15\,
            carryinitout => \bfn_7_25_0_\
        );

    \IN_MUX_bfv_13_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_24_0_\
        );

    \IN_MUX_bfv_13_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ppm_encoder_1.counter24_0_data_tmp_7\,
            carryinitout => \bfn_13_25_0_\
        );

    \IN_MUX_bfv_1_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_17_0_\
        );

    \IN_MUX_bfv_1_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \uart_frame_decoder.un1_WDT_cry_7\,
            carryinitout => \bfn_1_18_0_\
        );

    \IN_MUX_bfv_11_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_24_0_\
        );

    \IN_MUX_bfv_11_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ppm_encoder_1.un1_counter_13_cry_7\,
            carryinitout => \bfn_11_25_0_\
        );

    \IN_MUX_bfv_11_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ppm_encoder_1.un1_counter_13_cry_15\,
            carryinitout => \bfn_11_26_0_\
        );

    \reset_module_System.reset_RNITC69\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__24524\,
            GLOBALBUFFEROUTPUT => reset_system_g
        );

    \frame_decoder_dv_c_0_g_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__14886\,
            GLOBALBUFFEROUTPUT => frame_decoder_dv_c_0_g
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \ppm_encoder_1.PPM_STATE_fast_RNI9VGK_0_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__20943\,
            GLOBALBUFFEROUTPUT => \ppm_encoder_1.N_238_i_0_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \ppm_encoder_1.counter24_0_I_57_c_RNIGCO83_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__24360\,
            GLOBALBUFFEROUTPUT => \ppm_encoder_1.N_512_g\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \uart_frame_decoder.WDT_0_LC_1_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9174\,
            in2 => \N__9858\,
            in3 => \N__9857\,
            lcout => \uart_frame_decoder.WDTZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_1_17_0_\,
            carryout => \uart_frame_decoder.un1_WDT_cry_0\,
            clk => \N__23875\,
            ce => 'H',
            sr => \N__9261\
        );

    \uart_frame_decoder.WDT_1_LC_1_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9216\,
            in2 => \_gnd_net_\,
            in3 => \N__9210\,
            lcout => \uart_frame_decoder.WDTZ0Z_1\,
            ltout => OPEN,
            carryin => \uart_frame_decoder.un1_WDT_cry_0\,
            carryout => \uart_frame_decoder.un1_WDT_cry_1\,
            clk => \N__23875\,
            ce => 'H',
            sr => \N__9261\
        );

    \uart_frame_decoder.WDT_2_LC_1_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9207\,
            in2 => \_gnd_net_\,
            in3 => \N__9201\,
            lcout => \uart_frame_decoder.WDTZ0Z_2\,
            ltout => OPEN,
            carryin => \uart_frame_decoder.un1_WDT_cry_1\,
            carryout => \uart_frame_decoder.un1_WDT_cry_2\,
            clk => \N__23875\,
            ce => 'H',
            sr => \N__9261\
        );

    \uart_frame_decoder.WDT_3_LC_1_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9198\,
            in2 => \_gnd_net_\,
            in3 => \N__9192\,
            lcout => \uart_frame_decoder.WDTZ0Z_3\,
            ltout => OPEN,
            carryin => \uart_frame_decoder.un1_WDT_cry_2\,
            carryout => \uart_frame_decoder.un1_WDT_cry_3\,
            clk => \N__23875\,
            ce => 'H',
            sr => \N__9261\
        );

    \uart_frame_decoder.WDT_4_LC_1_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9804\,
            in2 => \_gnd_net_\,
            in3 => \N__9189\,
            lcout => \uart_frame_decoder.WDTZ0Z_4\,
            ltout => OPEN,
            carryin => \uart_frame_decoder.un1_WDT_cry_3\,
            carryout => \uart_frame_decoder.un1_WDT_cry_4\,
            clk => \N__23875\,
            ce => 'H',
            sr => \N__9261\
        );

    \uart_frame_decoder.WDT_5_LC_1_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9831\,
            in2 => \_gnd_net_\,
            in3 => \N__9186\,
            lcout => \uart_frame_decoder.WDTZ0Z_5\,
            ltout => OPEN,
            carryin => \uart_frame_decoder.un1_WDT_cry_4\,
            carryout => \uart_frame_decoder.un1_WDT_cry_5\,
            clk => \N__23875\,
            ce => 'H',
            sr => \N__9261\
        );

    \uart_frame_decoder.WDT_6_LC_1_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9843\,
            in2 => \_gnd_net_\,
            in3 => \N__9183\,
            lcout => \uart_frame_decoder.WDTZ0Z_6\,
            ltout => OPEN,
            carryin => \uart_frame_decoder.un1_WDT_cry_5\,
            carryout => \uart_frame_decoder.un1_WDT_cry_6\,
            clk => \N__23875\,
            ce => 'H',
            sr => \N__9261\
        );

    \uart_frame_decoder.WDT_7_LC_1_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9818\,
            in2 => \_gnd_net_\,
            in3 => \N__9180\,
            lcout => \uart_frame_decoder.WDTZ0Z_7\,
            ltout => OPEN,
            carryin => \uart_frame_decoder.un1_WDT_cry_6\,
            carryout => \uart_frame_decoder.un1_WDT_cry_7\,
            clk => \N__23875\,
            ce => 'H',
            sr => \N__9261\
        );

    \uart_frame_decoder.WDT_8_LC_1_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9687\,
            in2 => \_gnd_net_\,
            in3 => \N__9177\,
            lcout => \uart_frame_decoder.WDTZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_1_18_0_\,
            carryout => \uart_frame_decoder.un1_WDT_cry_8\,
            clk => \N__23871\,
            ce => 'H',
            sr => \N__9257\
        );

    \uart_frame_decoder.WDT_9_LC_1_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9882\,
            in2 => \_gnd_net_\,
            in3 => \N__9243\,
            lcout => \uart_frame_decoder.WDTZ0Z_9\,
            ltout => OPEN,
            carryin => \uart_frame_decoder.un1_WDT_cry_8\,
            carryout => \uart_frame_decoder.un1_WDT_cry_9\,
            clk => \N__23871\,
            ce => 'H',
            sr => \N__9257\
        );

    \uart_frame_decoder.WDT_10_LC_1_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9924\,
            in2 => \_gnd_net_\,
            in3 => \N__9240\,
            lcout => \uart_frame_decoder.WDTZ0Z_10\,
            ltout => OPEN,
            carryin => \uart_frame_decoder.un1_WDT_cry_9\,
            carryout => \uart_frame_decoder.un1_WDT_cry_10\,
            clk => \N__23871\,
            ce => 'H',
            sr => \N__9257\
        );

    \uart_frame_decoder.WDT_11_LC_1_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9939\,
            in2 => \_gnd_net_\,
            in3 => \N__9237\,
            lcout => \uart_frame_decoder.WDTZ0Z_11\,
            ltout => OPEN,
            carryin => \uart_frame_decoder.un1_WDT_cry_10\,
            carryout => \uart_frame_decoder.un1_WDT_cry_11\,
            clk => \N__23871\,
            ce => 'H',
            sr => \N__9257\
        );

    \uart_frame_decoder.WDT_12_LC_1_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9897\,
            in2 => \_gnd_net_\,
            in3 => \N__9234\,
            lcout => \uart_frame_decoder.WDTZ0Z_12\,
            ltout => OPEN,
            carryin => \uart_frame_decoder.un1_WDT_cry_11\,
            carryout => \uart_frame_decoder.un1_WDT_cry_12\,
            clk => \N__23871\,
            ce => 'H',
            sr => \N__9257\
        );

    \uart_frame_decoder.WDT_13_LC_1_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9911\,
            in2 => \_gnd_net_\,
            in3 => \N__9231\,
            lcout => \uart_frame_decoder.WDTZ0Z_13\,
            ltout => OPEN,
            carryin => \uart_frame_decoder.un1_WDT_cry_12\,
            carryout => \uart_frame_decoder.un1_WDT_cry_13\,
            clk => \N__23871\,
            ce => 'H',
            sr => \N__9257\
        );

    \uart_frame_decoder.WDT_14_LC_1_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9767\,
            in2 => \_gnd_net_\,
            in3 => \N__9228\,
            lcout => \uart_frame_decoder.WDTZ0Z_14\,
            ltout => OPEN,
            carryin => \uart_frame_decoder.un1_WDT_cry_13\,
            carryout => \uart_frame_decoder.un1_WDT_cry_14\,
            clk => \N__23871\,
            ce => 'H',
            sr => \N__9257\
        );

    \uart_frame_decoder.WDT_15_LC_1_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9786\,
            in2 => \_gnd_net_\,
            in3 => \N__9225\,
            lcout => \uart_frame_decoder.WDTZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23871\,
            ce => 'H',
            sr => \N__9257\
        );

    \uart_frame_decoder.count8_cry_0_c_LC_1_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9305\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_19_0_\,
            carryout => \uart_frame_decoder.count8_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.count8_cry_1_c_inv_LC_1_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9222\,
            in2 => \_gnd_net_\,
            in3 => \N__9981\,
            lcout => \uart_frame_decoder.count8_axb_1\,
            ltout => OPEN,
            carryin => \uart_frame_decoder.count8_cry_0\,
            carryout => \uart_frame_decoder.count8_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.count8_cry_2_c_inv_LC_1_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9294\,
            in2 => \N__24690\,
            in3 => \N__9997\,
            lcout => \uart_frame_decoder.count_i_2\,
            ltout => OPEN,
            carryin => \uart_frame_decoder.count8_cry_1\,
            carryout => \uart_frame_decoder.count8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.count8_THRU_LUT4_0_LC_1_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9288\,
            lcout => \uart_frame_decoder.count8_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.count_1_LC_1_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010100101"
        )
    port map (
            in0 => \N__9982\,
            in1 => \_gnd_net_\,
            in2 => \N__9273\,
            in3 => \N__9284\,
            lcout => \uart_frame_decoder.countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23866\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.count_2_LC_1_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000101010000"
        )
    port map (
            in0 => \N__9285\,
            in1 => \N__9272\,
            in2 => \N__10002\,
            in3 => \N__9983\,
            lcout => \uart_frame_decoder.countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23866\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.count8_cry_2_c_RNICKS21_LC_1_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011101100"
        )
    port map (
            in0 => \N__13116\,
            in1 => \N__24507\,
            in2 => \N__13173\,
            in3 => \N__13004\,
            lcout => \uart_frame_decoder.count8_cry_2_c_RNICKSZ0Z21\,
            ltout => \uart_frame_decoder.count8_cry_2_c_RNICKSZ0Z21_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.count_0_LC_1_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110000000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10860\,
            in2 => \N__9276\,
            in3 => \N__9965\,
            lcout => \uart_frame_decoder.count8_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23866\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_1.source_data_1_4_LC_1_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010010111000"
        )
    port map (
            in0 => \N__11403\,
            in1 => \N__14946\,
            in2 => \N__16067\,
            in3 => \N__11439\,
            lcout => scaler_1_data_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23862\,
            ce => 'H',
            sr => \N__23358\
        );

    \scaler_4.source_data_1_4_LC_1_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001011011000"
        )
    port map (
            in0 => \N__14947\,
            in1 => \N__10481\,
            in2 => \N__16091\,
            in3 => \N__10511\,
            lcout => scaler_4_data_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23862\,
            ce => 'H',
            sr => \N__23358\
        );

    \uart_frame_decoder.count_RNIV5MS_0_LC_1_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111111111111"
        )
    port map (
            in0 => \N__13172\,
            in1 => \_gnd_net_\,
            in2 => \N__13119\,
            in3 => \N__9961\,
            lcout => \uart_frame_decoder.count_RNIV5MSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.source_data_valid_2_sqmuxa_i_LC_1_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13112\,
            in2 => \_gnd_net_\,
            in3 => \N__23496\,
            lcout => \uart_frame_decoder.source_data_valid_2_sqmuxa_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.count8_cry_0_c_inv_LC_1_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__9306\,
            in1 => \N__24716\,
            in2 => \_gnd_net_\,
            in3 => \N__9960\,
            lcout => \uart_frame_decoder.count8_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.source_CH2data_esr_0_LC_1_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11245\,
            lcout => \frame_decoder_CH2data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23857\,
            ce => \N__10221\,
            sr => \N__23362\
        );

    \uart_frame_decoder.source_CH2data_esr_1_LC_1_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12777\,
            lcout => \frame_decoder_CH2data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23857\,
            ce => \N__10221\,
            sr => \N__23362\
        );

    \uart_frame_decoder.source_CH2data_esr_2_LC_1_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10977\,
            lcout => \frame_decoder_CH2data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23857\,
            ce => \N__10221\,
            sr => \N__23362\
        );

    \uart_frame_decoder.source_CH2data_esr_3_LC_1_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12528\,
            lcout => \frame_decoder_CH2data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23857\,
            ce => \N__10221\,
            sr => \N__23362\
        );

    \uart_frame_decoder.source_CH2data_esr_4_LC_1_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15093\,
            lcout => \frame_decoder_CH2data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23857\,
            ce => \N__10221\,
            sr => \N__23362\
        );

    \uart_frame_decoder.source_CH2data_esr_5_LC_1_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11084\,
            lcout => \frame_decoder_CH2data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23857\,
            ce => \N__10221\,
            sr => \N__23362\
        );

    \uart_frame_decoder.source_CH2data_esr_6_LC_1_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12438\,
            lcout => \frame_decoder_CH2data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23857\,
            ce => \N__10221\,
            sr => \N__23362\
        );

    \uart_frame_decoder.source_CH2data_esr_7_LC_1_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11584\,
            lcout => \frame_decoder_CH2data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23857\,
            ce => \N__10221\,
            sr => \N__23362\
        );

    \uart_frame_decoder.source_offset3data_esr_0_LC_1_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11241\,
            lcout => \frame_decoder_OFF3data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23853\,
            ce => \N__11912\,
            sr => \N__23367\
        );

    \uart_frame_decoder.source_offset3data_esr_2_LC_1_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10978\,
            lcout => \frame_decoder_OFF3data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23853\,
            ce => \N__11912\,
            sr => \N__23367\
        );

    \uart_frame_decoder.source_offset3data_esr_3_LC_1_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12529\,
            lcout => \frame_decoder_OFF3data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23853\,
            ce => \N__11912\,
            sr => \N__23367\
        );

    \uart_frame_decoder.source_offset3data_esr_4_LC_1_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15094\,
            lcout => \frame_decoder_OFF3data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23853\,
            ce => \N__11912\,
            sr => \N__23367\
        );

    \uart_frame_decoder.source_offset3data_esr_5_LC_1_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11085\,
            lcout => \frame_decoder_OFF3data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23853\,
            ce => \N__11912\,
            sr => \N__23367\
        );

    \uart_frame_decoder.source_offset3data_esr_6_LC_1_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__12439\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \frame_decoder_OFF3data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23853\,
            ce => \N__11912\,
            sr => \N__23367\
        );

    \uart_frame_decoder.source_offset3data_esr_7_LC_1_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11585\,
            lcout => \frame_decoder_OFF3data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23853\,
            ce => \N__11912\,
            sr => \N__23367\
        );

    \scaler_3.un3_source_data_un3_source_data_0_cry_0_c_LC_1_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13459\,
            in2 => \N__13503\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_23_0_\,
            carryout => \scaler_3.un3_source_data_0_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_3.un3_source_data_un3_source_data_0_cry_0_c_RNILO5I_LC_1_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10314\,
            in2 => \N__11934\,
            in3 => \N__9321\,
            lcout => \scaler_3.un2_source_data_0\,
            ltout => OPEN,
            carryin => \scaler_3.un3_source_data_0_cry_0\,
            carryout => \scaler_3.un3_source_data_0_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_3.un3_source_data_un3_source_data_0_cry_1_c_RNIOS6I_LC_1_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10308\,
            in2 => \N__9318\,
            in3 => \N__9309\,
            lcout => \scaler_3.un3_source_data_0_cry_1_c_RNIOS6I\,
            ltout => OPEN,
            carryin => \scaler_3.un3_source_data_0_cry_1\,
            carryout => \scaler_3.un3_source_data_0_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_3.un3_source_data_un3_source_data_0_cry_2_c_RNIR08I_LC_1_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10302\,
            in2 => \N__9378\,
            in3 => \N__9369\,
            lcout => \scaler_3.un3_source_data_0_cry_2_c_RNIR08I\,
            ltout => OPEN,
            carryin => \scaler_3.un3_source_data_0_cry_2\,
            carryout => \scaler_3.un3_source_data_0_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_3.un3_source_data_un3_source_data_0_cry_3_c_RNIU49I_LC_1_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10296\,
            in2 => \N__9366\,
            in3 => \N__9357\,
            lcout => \scaler_3.un3_source_data_0_cry_3_c_RNIU49I\,
            ltout => OPEN,
            carryin => \scaler_3.un3_source_data_0_cry_3\,
            carryout => \scaler_3.un3_source_data_0_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_3.un3_source_data_un3_source_data_0_cry_4_c_RNI19AI_LC_1_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10290\,
            in2 => \N__9354\,
            in3 => \N__9345\,
            lcout => \scaler_3.un3_source_data_0_cry_4_c_RNI19AI\,
            ltout => OPEN,
            carryin => \scaler_3.un3_source_data_0_cry_4\,
            carryout => \scaler_3.un3_source_data_0_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_3.un3_source_data_un3_source_data_0_cry_5_c_RNI4DBI_LC_1_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10284\,
            in2 => \N__9342\,
            in3 => \N__9333\,
            lcout => \scaler_3.un3_source_data_0_cry_5_c_RNI4DBI\,
            ltout => OPEN,
            carryin => \scaler_3.un3_source_data_0_cry_5\,
            carryout => \scaler_3.un3_source_data_0_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_3.un3_source_data_un3_source_data_0_cry_6_c_RNI7HCI_LC_1_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10191\,
            in2 => \_gnd_net_\,
            in3 => \N__9330\,
            lcout => \scaler_3.un3_source_data_0_cry_6_c_RNI7HCI\,
            ltout => OPEN,
            carryin => \scaler_3.un3_source_data_0_cry_6\,
            carryout => \scaler_3.un3_source_data_0_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_3.un3_source_data_un3_source_data_0_cry_7_c_RNI8JDI_LC_1_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9468\,
            in2 => \N__24750\,
            in3 => \N__9327\,
            lcout => \scaler_3.un3_source_data_0_cry_7_c_RNI8JDI\,
            ltout => OPEN,
            carryin => \bfn_1_24_0_\,
            carryout => \scaler_3.un3_source_data_0_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_3.un3_source_data_un3_source_data_0_cry_8_c_RNIRV25_LC_1_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9324\,
            lcout => \scaler_3.un3_source_data_0_cry_8_c_RNIRV25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_RNIQ6GQ_9_LC_1_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13289\,
            in2 => \_gnd_net_\,
            in3 => \N__23501\,
            lcout => \uart_frame_decoder.source_offset4data_1_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_RNIOK9H_4_LC_1_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__10020\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13118\,
            lcout => \uart_frame_decoder.source_CH3data_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.un3_source_data_un3_source_data_0_axb_7_LC_1_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9707\,
            in2 => \_gnd_net_\,
            in3 => \N__11498\,
            lcout => \scaler_4.un3_source_data_0_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_3.un2_source_data_0_cry_1_c_RNO_LC_1_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__11682\,
            in1 => \N__13504\,
            in2 => \_gnd_net_\,
            in3 => \N__13460\,
            lcout => \scaler_3.un2_source_data_0_cry_1_c_RNO_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_3.N_795_i_l_ofx_LC_1_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10206\,
            in2 => \_gnd_net_\,
            in3 => \N__10278\,
            lcout => \scaler_3.N_795_i_l_ofxZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_3.un2_source_data_0_cry_1_c_LC_1_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11683\,
            in2 => \N__9462\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_25_0_\,
            carryout => \scaler_3.un2_source_data_0_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_3.source_data_1_esr_6_LC_1_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9446\,
            in2 => \N__11690\,
            in3 => \N__9453\,
            lcout => scaler_3_data_6,
            ltout => OPEN,
            carryin => \scaler_3.un2_source_data_0_cry_1\,
            carryout => \scaler_3.un2_source_data_0_cry_2\,
            clk => \N__23843\,
            ce => \N__11965\,
            sr => \N__23388\
        );

    \scaler_3.source_data_1_esr_7_LC_1_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9428\,
            in2 => \N__9450\,
            in3 => \N__9435\,
            lcout => scaler_3_data_7,
            ltout => OPEN,
            carryin => \scaler_3.un2_source_data_0_cry_2\,
            carryout => \scaler_3.un2_source_data_0_cry_3\,
            clk => \N__23843\,
            ce => \N__11965\,
            sr => \N__23388\
        );

    \scaler_3.source_data_1_esr_8_LC_1_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9410\,
            in2 => \N__9432\,
            in3 => \N__9417\,
            lcout => scaler_3_data_8,
            ltout => OPEN,
            carryin => \scaler_3.un2_source_data_0_cry_3\,
            carryout => \scaler_3.un2_source_data_0_cry_4\,
            clk => \N__23843\,
            ce => \N__11965\,
            sr => \N__23388\
        );

    \scaler_3.source_data_1_esr_9_LC_1_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9392\,
            in2 => \N__9414\,
            in3 => \N__9399\,
            lcout => scaler_3_data_9,
            ltout => OPEN,
            carryin => \scaler_3.un2_source_data_0_cry_4\,
            carryout => \scaler_3.un2_source_data_0_cry_5\,
            clk => \N__23843\,
            ce => \N__11965\,
            sr => \N__23388\
        );

    \scaler_3.source_data_1_esr_10_LC_1_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9533\,
            in2 => \N__9396\,
            in3 => \N__9381\,
            lcout => scaler_3_data_10,
            ltout => OPEN,
            carryin => \scaler_3.un2_source_data_0_cry_5\,
            carryout => \scaler_3.un2_source_data_0_cry_6\,
            clk => \N__23843\,
            ce => \N__11965\,
            sr => \N__23388\
        );

    \scaler_3.source_data_1_esr_11_LC_1_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9515\,
            in2 => \N__9537\,
            in3 => \N__9522\,
            lcout => scaler_3_data_11,
            ltout => OPEN,
            carryin => \scaler_3.un2_source_data_0_cry_6\,
            carryout => \scaler_3.un2_source_data_0_cry_7\,
            clk => \N__23843\,
            ce => \N__11965\,
            sr => \N__23388\
        );

    \scaler_3.source_data_1_esr_12_LC_1_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9497\,
            in2 => \N__9519\,
            in3 => \N__9504\,
            lcout => scaler_3_data_12,
            ltout => OPEN,
            carryin => \scaler_3.un2_source_data_0_cry_7\,
            carryout => \scaler_3.un2_source_data_0_cry_8\,
            clk => \N__23843\,
            ce => \N__11965\,
            sr => \N__23388\
        );

    \scaler_3.source_data_1_esr_13_LC_1_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9501\,
            in2 => \N__9486\,
            in3 => \N__9474\,
            lcout => scaler_3_data_13,
            ltout => OPEN,
            carryin => \bfn_1_26_0_\,
            carryout => \scaler_3.un2_source_data_0_cry_9\,
            clk => \N__23837\,
            ce => \N__11964\,
            sr => \N__23394\
        );

    \scaler_3.source_data_1_esr_14_LC_1_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9471\,
            lcout => scaler_3_data_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23837\,
            ce => \N__11964\,
            sr => \N__23394\
        );

    \scaler_4.source_data_1_esr_5_LC_1_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__10440\,
            in1 => \N__10474\,
            in2 => \_gnd_net_\,
            in3 => \N__10512\,
            lcout => scaler_4_data_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23837\,
            ce => \N__11964\,
            sr => \N__23394\
        );

    \uart_frame_decoder.source_offset4data_esr_0_LC_1_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11252\,
            lcout => \frame_decoder_OFF4data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23832\,
            ce => \N__9549\,
            sr => \N__23398\
        );

    \uart_frame_decoder.source_offset4data_esr_1_LC_1_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__12786\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \frame_decoder_OFF4data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23832\,
            ce => \N__9549\,
            sr => \N__23398\
        );

    \uart_frame_decoder.source_offset4data_esr_2_LC_1_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10985\,
            lcout => \frame_decoder_OFF4data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23832\,
            ce => \N__9549\,
            sr => \N__23398\
        );

    \uart_frame_decoder.source_offset4data_esr_3_LC_1_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12545\,
            lcout => \frame_decoder_OFF4data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23832\,
            ce => \N__9549\,
            sr => \N__23398\
        );

    \uart_frame_decoder.source_offset4data_esr_4_LC_1_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__15107\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \frame_decoder_OFF4data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23832\,
            ce => \N__9549\,
            sr => \N__23398\
        );

    \uart_frame_decoder.source_offset4data_esr_5_LC_1_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__11093\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \frame_decoder_OFF4data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23832\,
            ce => \N__9549\,
            sr => \N__23398\
        );

    \uart_frame_decoder.source_offset4data_esr_6_LC_1_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12456\,
            lcout => \frame_decoder_OFF4data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23832\,
            ce => \N__9549\,
            sr => \N__23398\
        );

    \uart_frame_decoder.source_offset4data_esr_7_LC_1_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11586\,
            lcout => \frame_decoder_OFF4data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23832\,
            ce => \N__9549\,
            sr => \N__23398\
        );

    \uart_frame_decoder.source_CH4data_esr_0_LC_1_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__11253\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \frame_decoder_CH4data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23828\,
            ce => \N__11484\,
            sr => \N__23402\
        );

    \uart_frame_decoder.source_CH4data_esr_2_LC_1_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10986\,
            lcout => \frame_decoder_CH4data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23828\,
            ce => \N__11484\,
            sr => \N__23402\
        );

    \uart_frame_decoder.source_CH4data_esr_3_LC_1_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12546\,
            lcout => \frame_decoder_CH4data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23828\,
            ce => \N__11484\,
            sr => \N__23402\
        );

    \uart_frame_decoder.source_CH4data_esr_4_LC_1_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15108\,
            lcout => \frame_decoder_CH4data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23828\,
            ce => \N__11484\,
            sr => \N__23402\
        );

    \uart_frame_decoder.source_CH4data_esr_5_LC_1_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__11094\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \frame_decoder_CH4data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23828\,
            ce => \N__11484\,
            sr => \N__23402\
        );

    \uart_frame_decoder.source_CH4data_esr_6_LC_1_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12457\,
            lcout => \frame_decoder_CH4data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23828\,
            ce => \N__11484\,
            sr => \N__23402\
        );

    \uart_frame_decoder.source_CH4data_esr_1_LC_1_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12787\,
            lcout => \frame_decoder_CH4data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23828\,
            ce => \N__11484\,
            sr => \N__23402\
        );

    \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_LC_1_29_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10503\,
            in2 => \N__10482\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_29_0_\,
            carryout => \scaler_4.un3_source_data_0_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_RNIOOII_LC_1_29_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9675\,
            in2 => \N__9669\,
            in3 => \N__9657\,
            lcout => \scaler_4.un2_source_data_0\,
            ltout => OPEN,
            carryin => \scaler_4.un3_source_data_0_cry_0\,
            carryout => \scaler_4.un3_source_data_0_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.un3_source_data_un3_source_data_0_cry_1_c_RNIRSJI_LC_1_29_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9654\,
            in2 => \N__9648\,
            in3 => \N__9636\,
            lcout => \scaler_4.un3_source_data_0_cry_1_c_RNIRSJI\,
            ltout => OPEN,
            carryin => \scaler_4.un3_source_data_0_cry_1\,
            carryout => \scaler_4.un3_source_data_0_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.un3_source_data_un3_source_data_0_cry_2_c_RNIU0LI_LC_1_29_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9633\,
            in2 => \N__9627\,
            in3 => \N__9615\,
            lcout => \scaler_4.un3_source_data_0_cry_2_c_RNIU0LI\,
            ltout => OPEN,
            carryin => \scaler_4.un3_source_data_0_cry_2\,
            carryout => \scaler_4.un3_source_data_0_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.un3_source_data_un3_source_data_0_cry_3_c_RNI15MI_LC_1_29_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9612\,
            in2 => \N__9606\,
            in3 => \N__9594\,
            lcout => \scaler_4.un3_source_data_0_cry_3_c_RNI15MI\,
            ltout => OPEN,
            carryin => \scaler_4.un3_source_data_0_cry_3\,
            carryout => \scaler_4.un3_source_data_0_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.un3_source_data_un3_source_data_0_cry_4_c_RNI49NI_LC_1_29_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9591\,
            in2 => \N__9582\,
            in3 => \N__9573\,
            lcout => \scaler_4.un3_source_data_0_cry_4_c_RNI49NI\,
            ltout => OPEN,
            carryin => \scaler_4.un3_source_data_0_cry_4\,
            carryout => \scaler_4.un3_source_data_0_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.un3_source_data_un3_source_data_0_cry_5_c_RNI7DOI_LC_1_29_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9570\,
            in2 => \N__9564\,
            in3 => \N__9552\,
            lcout => \scaler_4.un3_source_data_0_cry_5_c_RNI7DOI\,
            ltout => OPEN,
            carryin => \scaler_4.un3_source_data_0_cry_5\,
            carryout => \scaler_4.un3_source_data_0_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.un3_source_data_un3_source_data_0_cry_6_c_RNIAHPI_LC_1_29_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9729\,
            in2 => \_gnd_net_\,
            in3 => \N__9717\,
            lcout => \scaler_4.un3_source_data_0_cry_6_c_RNIAHPI\,
            ltout => OPEN,
            carryin => \scaler_4.un3_source_data_0_cry_6\,
            carryout => \scaler_4.un3_source_data_0_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.un3_source_data_un3_source_data_0_cry_7_c_RNIBJQI_LC_1_30_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9693\,
            in2 => \N__24768\,
            in3 => \N__9714\,
            lcout => \scaler_4.un3_source_data_0_cry_7_c_RNIBJQI\,
            ltout => OPEN,
            carryin => \bfn_1_30_0_\,
            carryout => \scaler_4.un3_source_data_0_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.un3_source_data_un3_source_data_0_cry_8_c_RNIS918_LC_1_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9711\,
            lcout => \scaler_4.un3_source_data_0_cry_8_c_RNIS918\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.N_807_i_l_ofx_LC_1_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__9708\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11505\,
            lcout => \scaler_4.N_807_i_l_ofxZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.bit_Count_0_LC_2_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011001100"
        )
    port map (
            in0 => \N__10693\,
            in1 => \N__12876\,
            in2 => \_gnd_net_\,
            in3 => \N__12040\,
            lcout => \uart.bit_CountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23878\,
            ce => 'H',
            sr => \N__23341\
        );

    \uart.bit_Count_2_LC_2_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000110100010"
        )
    port map (
            in0 => \N__12985\,
            in1 => \N__12042\,
            in2 => \N__10701\,
            in3 => \N__10707\,
            lcout => \uart.bit_CountZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23878\,
            ce => 'H',
            sr => \N__23341\
        );

    \uart.bit_Count_1_LC_2_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110000010101010"
        )
    port map (
            in0 => \N__12929\,
            in1 => \N__12877\,
            in2 => \N__10700\,
            in3 => \N__12041\,
            lcout => \uart.bit_CountZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23878\,
            ce => 'H',
            sr => \N__23341\
        );

    \uart.state_RNO_1_3_LC_2_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011101110"
        )
    port map (
            in0 => \N__10671\,
            in1 => \N__12277\,
            in2 => \_gnd_net_\,
            in3 => \N__24486\,
            lcout => \uart.state_srsts_i_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.data_Aux_RNO_0_1_LC_2_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__12981\,
            in1 => \N__12923\,
            in2 => \_gnd_net_\,
            in3 => \N__12862\,
            lcout => \uart.data_Auxce_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.WDT_RNIDK7E_8_LC_2_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__9895\,
            in1 => \N__9937\,
            in2 => \_gnd_net_\,
            in3 => \N__9686\,
            lcout => \uart_frame_decoder.WDT8lto13_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.WDT_RNIAGPB_10_LC_2_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100011111"
        )
    port map (
            in0 => \N__9938\,
            in1 => \N__9923\,
            in2 => \N__9912\,
            in3 => \N__9896\,
            lcout => OPEN,
            ltout => \uart_frame_decoder.WDT_RNIAGPBZ0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.WDT_RNIM8N32_9_LC_2_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101100001111"
        )
    port map (
            in0 => \N__9881\,
            in1 => \N__9792\,
            in2 => \N__9870\,
            in3 => \N__9867\,
            lcout => \uart_frame_decoder.WDT8lt14_0\,
            ltout => \uart_frame_decoder.WDT8lt14_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.WDT_RNI17K92_15_LC_2_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9784\,
            in2 => \N__9861\,
            in3 => \N__9763\,
            lcout => \uart_frame_decoder.WDT8_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.WDT_RNIM6B11_4_LC_2_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__9842\,
            in1 => \N__9830\,
            in2 => \N__9819\,
            in3 => \N__9803\,
            lcout => \uart_frame_decoder.WDT_RNIM6B11Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.WDT_RNIJUEI2_15_LC_2_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010011"
        )
    port map (
            in0 => \N__9785\,
            in1 => \N__13062\,
            in2 => \N__9768\,
            in3 => \N__9747\,
            lcout => \uart_frame_decoder.WDT_RNIJUEI2Z0Z_15\,
            ltout => \uart_frame_decoder.WDT_RNIJUEI2Z0Z_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_3_LC_2_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101010101010"
        )
    port map (
            in0 => \N__10118\,
            in1 => \_gnd_net_\,
            in2 => \N__9741\,
            in3 => \N__9738\,
            lcout => \uart_frame_decoder.state_1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23872\,
            ce => 'H',
            sr => \N__23343\
        );

    \uart_frame_decoder.state_1_RNINJ9H_3_LC_2_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__9737\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13061\,
            lcout => \uart_frame_decoder.source_CH2data_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_1_LC_2_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__10779\,
            in1 => \N__12704\,
            in2 => \N__11165\,
            in3 => \N__13234\,
            lcout => \uart_frame_decoder.state_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23867\,
            ce => 'H',
            sr => \N__23345\
        );

    \uart_frame_decoder.state_1_2_LC_2_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__13235\,
            in1 => \N__10032\,
            in2 => \N__12708\,
            in3 => \N__11127\,
            lcout => \uart_frame_decoder.state_1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23867\,
            ce => 'H',
            sr => \N__23345\
        );

    \uart_frame_decoder.state_1_RNIMI9H_2_LC_2_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10031\,
            in2 => \_gnd_net_\,
            in3 => \N__13089\,
            lcout => \uart_frame_decoder.source_CH1data_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_4_LC_2_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111010101010"
        )
    port map (
            in0 => \N__10235\,
            in1 => \N__10016\,
            in2 => \_gnd_net_\,
            in3 => \N__13236\,
            lcout => \uart_frame_decoder.state_1Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23867\,
            ce => 'H',
            sr => \N__23345\
        );

    \uart_frame_decoder.count_RNIM2UL1_2_LC_2_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010111"
        )
    port map (
            in0 => \N__10001\,
            in1 => \N__9984\,
            in2 => \N__9966\,
            in3 => \N__10856\,
            lcout => \uart_frame_decoder.state_1_ns_0_i_o2_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_RNO_1_0_LC_2_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111000"
        )
    port map (
            in0 => \N__11123\,
            in1 => \N__12698\,
            in2 => \N__10833\,
            in3 => \N__10845\,
            lcout => OPEN,
            ltout => \uart_frame_decoder.state_1_ns_i_i_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_0_LC_2_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000001000000011"
        )
    port map (
            in0 => \N__10839\,
            in1 => \N__13301\,
            in2 => \N__9942\,
            in3 => \N__13246\,
            lcout => \uart_frame_decoder.state_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23863\,
            ce => 'H',
            sr => \N__23348\
        );

    \uart_frame_decoder.source_offset2data_esr_0_LC_2_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11213\,
            lcout => \frame_decoder_OFF2data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23858\,
            ce => \N__10104\,
            sr => \N__23352\
        );

    \uart_frame_decoder.source_offset2data_esr_1_LC_2_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12741\,
            lcout => \frame_decoder_OFF2data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23858\,
            ce => \N__10104\,
            sr => \N__23352\
        );

    \uart_frame_decoder.source_offset2data_esr_2_LC_2_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10945\,
            lcout => \frame_decoder_OFF2data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23858\,
            ce => \N__10104\,
            sr => \N__23352\
        );

    \uart_frame_decoder.source_offset2data_esr_3_LC_2_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12509\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \frame_decoder_OFF2data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23858\,
            ce => \N__10104\,
            sr => \N__23352\
        );

    \uart_frame_decoder.source_offset2data_esr_4_LC_2_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15073\,
            lcout => \frame_decoder_OFF2data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23858\,
            ce => \N__10104\,
            sr => \N__23352\
        );

    \uart_frame_decoder.source_offset2data_esr_5_LC_2_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11047\,
            lcout => \frame_decoder_OFF2data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23858\,
            ce => \N__10104\,
            sr => \N__23352\
        );

    \uart_frame_decoder.source_offset2data_esr_6_LC_2_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12417\,
            lcout => \frame_decoder_OFF2data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23858\,
            ce => \N__10104\,
            sr => \N__23352\
        );

    \uart_frame_decoder.source_offset2data_esr_7_LC_2_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11553\,
            lcout => \frame_decoder_OFF2data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23858\,
            ce => \N__10104\,
            sr => \N__23352\
        );

    \scaler_2.un3_source_data_un3_source_data_0_cry_0_c_LC_2_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15174\,
            in2 => \N__15222\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_21_0_\,
            carryout => \scaler_2.un3_source_data_0_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_2.un3_source_data_un3_source_data_0_cry_0_c_RNIIOOH_LC_2_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10095\,
            in2 => \N__10089\,
            in3 => \N__10080\,
            lcout => \scaler_2.un2_source_data_0\,
            ltout => OPEN,
            carryin => \scaler_2.un3_source_data_0_cry_0\,
            carryout => \scaler_2.un3_source_data_0_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_2.un3_source_data_un3_source_data_0_cry_1_c_RNILSPH_LC_2_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10077\,
            in2 => \N__10071\,
            in3 => \N__10059\,
            lcout => \scaler_2.un3_source_data_0_cry_1_c_RNILSPH\,
            ltout => OPEN,
            carryin => \scaler_2.un3_source_data_0_cry_1\,
            carryout => \scaler_2.un3_source_data_0_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_2.un3_source_data_un3_source_data_0_cry_2_c_RNIO0RH_LC_2_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10056\,
            in2 => \N__10050\,
            in3 => \N__10041\,
            lcout => \scaler_2.un3_source_data_0_cry_2_c_RNIO0RH\,
            ltout => OPEN,
            carryin => \scaler_2.un3_source_data_0_cry_2\,
            carryout => \scaler_2.un3_source_data_0_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_2.un3_source_data_un3_source_data_0_cry_3_c_RNIR4SH_LC_2_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10038\,
            in2 => \N__10182\,
            in3 => \N__10173\,
            lcout => \scaler_2.un3_source_data_0_cry_3_c_RNIR4SH\,
            ltout => OPEN,
            carryin => \scaler_2.un3_source_data_0_cry_3\,
            carryout => \scaler_2.un3_source_data_0_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_2.un3_source_data_un3_source_data_0_cry_4_c_RNIU8TH_LC_2_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10170\,
            in2 => \N__10164\,
            in3 => \N__10155\,
            lcout => \scaler_2.un3_source_data_0_cry_4_c_RNIU8TH\,
            ltout => OPEN,
            carryin => \scaler_2.un3_source_data_0_cry_4\,
            carryout => \scaler_2.un3_source_data_0_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_2.un3_source_data_un3_source_data_0_cry_5_c_RNI1DUH_LC_2_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10152\,
            in2 => \N__10146\,
            in3 => \N__10137\,
            lcout => \scaler_2.un3_source_data_0_cry_5_c_RNI1DUH\,
            ltout => OPEN,
            carryin => \scaler_2.un3_source_data_0_cry_5\,
            carryout => \scaler_2.un3_source_data_0_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_2.un3_source_data_un3_source_data_0_cry_6_c_RNI4HVH_LC_2_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10125\,
            in2 => \_gnd_net_\,
            in3 => \N__10134\,
            lcout => \scaler_2.un3_source_data_0_cry_6_c_RNI4HVH\,
            ltout => OPEN,
            carryin => \scaler_2.un3_source_data_0_cry_6\,
            carryout => \scaler_2.un3_source_data_0_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_2.un3_source_data_un3_source_data_0_cry_7_c_RNI5J0I_LC_2_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10242\,
            in2 => \N__24749\,
            in3 => \N__10131\,
            lcout => \scaler_2.un3_source_data_0_cry_7_c_RNI5J0I\,
            ltout => OPEN,
            carryin => \bfn_2_22_0_\,
            carryout => \scaler_2.un3_source_data_0_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_2.un3_source_data_un3_source_data_0_cry_8_c_RNIQL42_LC_2_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10128\,
            lcout => \scaler_2.un3_source_data_0_cry_8_c_RNIQL42\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_2.un3_source_data_un3_source_data_0_axb_7_LC_2_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10253\,
            in2 => \_gnd_net_\,
            in3 => \N__10265\,
            lcout => \scaler_2.un3_source_data_0_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_RNIJVFQ_2_LC_2_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__10119\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23498\,
            lcout => \uart_frame_decoder.source_CH1data_1_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_RNIO4GQ_7_LC_2_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__23499\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11654\,
            lcout => \uart_frame_decoder.source_offset2data_1_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_ns_0_i_a2_0_4_1_LC_2_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__11220\,
            in1 => \N__11554\,
            in2 => \N__11081\,
            in3 => \N__10953\,
            lcout => \uart_frame_decoder.N_79_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_2.N_783_i_l_ofx_LC_2_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__10266\,
            in1 => \_gnd_net_\,
            in2 => \N__10257\,
            in3 => \_gnd_net_\,
            lcout => \scaler_2.N_783_i_l_ofxZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_RNIK0GQ_3_LC_2_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10236\,
            in2 => \_gnd_net_\,
            in3 => \N__23495\,
            lcout => \uart_frame_decoder.source_CH2data_1_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_RNIPL9H_5_LC_2_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11603\,
            in2 => \_gnd_net_\,
            in3 => \N__13110\,
            lcout => \uart_frame_decoder.source_CH4data_1_sqmuxa\,
            ltout => \uart_frame_decoder.source_CH4data_1_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_RNIM2GQ_5_LC_2_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10209\,
            in3 => \N__23493\,
            lcout => \uart_frame_decoder.source_CH4data_1_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_3.un3_source_data_un3_source_data_0_axb_7_LC_2_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10202\,
            in2 => \_gnd_net_\,
            in3 => \N__10277\,
            lcout => \scaler_3.un3_source_data_0_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_RNISO9H_8_LC_2_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__13111\,
            in1 => \_gnd_net_\,
            in2 => \N__11637\,
            in3 => \_gnd_net_\,
            lcout => \uart_frame_decoder.source_offset3data_1_sqmuxa\,
            ltout => \uart_frame_decoder.source_offset3data_1_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_RNIP5GQ_8_LC_2_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__23494\,
            in1 => \_gnd_net_\,
            in2 => \N__10185\,
            in3 => \_gnd_net_\,
            lcout => \uart_frame_decoder.source_offset3data_1_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.source_CH3data_esr_0_LC_2_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11242\,
            lcout => \frame_decoder_CH3data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23844\,
            ce => \N__11445\,
            sr => \N__23374\
        );

    \uart_frame_decoder.source_CH3data_esr_1_LC_2_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12778\,
            lcout => \frame_decoder_CH3data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23844\,
            ce => \N__11445\,
            sr => \N__23374\
        );

    \uart_frame_decoder.source_CH3data_esr_2_LC_2_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10974\,
            lcout => \frame_decoder_CH3data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23844\,
            ce => \N__11445\,
            sr => \N__23374\
        );

    \uart_frame_decoder.source_CH3data_esr_3_LC_2_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12530\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \frame_decoder_CH3data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23844\,
            ce => \N__11445\,
            sr => \N__23374\
        );

    \uart_frame_decoder.source_CH3data_esr_4_LC_2_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__15095\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \frame_decoder_CH3data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23844\,
            ce => \N__11445\,
            sr => \N__23374\
        );

    \uart_frame_decoder.source_CH3data_esr_5_LC_2_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11086\,
            lcout => \frame_decoder_CH3data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23844\,
            ce => \N__11445\,
            sr => \N__23374\
        );

    \uart_frame_decoder.source_CH3data_esr_6_LC_2_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12455\,
            lcout => \frame_decoder_CH3data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23844\,
            ce => \N__11445\,
            sr => \N__23374\
        );

    \uart_frame_decoder.source_CH3data_esr_7_LC_2_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11580\,
            lcout => \frame_decoder_CH3data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23844\,
            ce => \N__11445\,
            sr => \N__23374\
        );

    \uart_frame_decoder.source_CH1data_esr_0_LC_2_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__11243\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \frame_decoder_CH1data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23838\,
            ce => \N__15017\,
            sr => \N__23382\
        );

    \uart_frame_decoder.source_CH1data_esr_2_LC_2_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10975\,
            lcout => \frame_decoder_CH1data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23838\,
            ce => \N__15017\,
            sr => \N__23382\
        );

    \uart_frame_decoder.source_CH1data_esr_3_LC_2_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12543\,
            lcout => \frame_decoder_CH1data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23838\,
            ce => \N__15017\,
            sr => \N__23382\
        );

    \uart_frame_decoder.source_CH1data_esr_1_LC_2_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__12779\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \frame_decoder_CH1data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23838\,
            ce => \N__15017\,
            sr => \N__23382\
        );

    \uart_frame_decoder.source_CH1data_esr_5_LC_2_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11082\,
            lcout => \frame_decoder_CH1data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23838\,
            ce => \N__15017\,
            sr => \N__23382\
        );

    \uart_frame_decoder.source_CH1data_esr_6_LC_2_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12458\,
            lcout => \frame_decoder_CH1data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23838\,
            ce => \N__15017\,
            sr => \N__23382\
        );

    \uart_frame_decoder.source_CH1data_esr_7_LC_2_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11581\,
            lcout => \frame_decoder_CH1data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23838\,
            ce => \N__15017\,
            sr => \N__23382\
        );

    \uart_frame_decoder.source_offset1data_esr_0_LC_2_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__11244\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \frame_decoder_OFF1data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23833\,
            ce => \N__13401\,
            sr => \N__23389\
        );

    \uart_frame_decoder.source_offset1data_esr_1_LC_2_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12788\,
            lcout => \frame_decoder_OFF1data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23833\,
            ce => \N__13401\,
            sr => \N__23389\
        );

    \uart_frame_decoder.source_offset1data_esr_2_LC_2_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10976\,
            lcout => \frame_decoder_OFF1data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23833\,
            ce => \N__13401\,
            sr => \N__23389\
        );

    \uart_frame_decoder.source_offset1data_esr_3_LC_2_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12544\,
            lcout => \frame_decoder_OFF1data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23833\,
            ce => \N__13401\,
            sr => \N__23389\
        );

    \uart_frame_decoder.source_offset1data_esr_4_LC_2_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15106\,
            lcout => \frame_decoder_OFF1data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23833\,
            ce => \N__13401\,
            sr => \N__23389\
        );

    \uart_frame_decoder.source_offset1data_esr_5_LC_2_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11083\,
            lcout => \frame_decoder_OFF1data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23833\,
            ce => \N__13401\,
            sr => \N__23389\
        );

    \uart_frame_decoder.source_offset1data_esr_6_LC_2_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12459\,
            lcout => \frame_decoder_OFF1data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23833\,
            ce => \N__13401\,
            sr => \N__23389\
        );

    \uart_frame_decoder.source_offset1data_esr_7_LC_2_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11582\,
            lcout => \frame_decoder_OFF1data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23833\,
            ce => \N__13401\,
            sr => \N__23389\
        );

    \scaler_1.un3_source_data_un3_source_data_0_cry_0_c_LC_2_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11395\,
            in2 => \N__11434\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_27_0_\,
            carryout => \scaler_1.un3_source_data_0_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_1.un3_source_data_un3_source_data_0_cry_0_c_RNIFOB11_LC_2_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10410\,
            in2 => \N__10401\,
            in3 => \N__10392\,
            lcout => \scaler_1.un2_source_data_0\,
            ltout => OPEN,
            carryin => \scaler_1.un3_source_data_0_cry_0\,
            carryout => \scaler_1.un3_source_data_0_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_1.un3_source_data_un3_source_data_0_cry_1_c_RNIISC11_LC_2_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10389\,
            in2 => \N__10380\,
            in3 => \N__10371\,
            lcout => \scaler_1.un3_source_data_0_cry_1_c_RNIISC11\,
            ltout => OPEN,
            carryin => \scaler_1.un3_source_data_0_cry_1\,
            carryout => \scaler_1.un3_source_data_0_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_1.un3_source_data_un3_source_data_0_cry_2_c_RNIL0E11_LC_2_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10368\,
            in2 => \N__10359\,
            in3 => \N__10350\,
            lcout => \scaler_1.un3_source_data_0_cry_2_c_RNIL0E11\,
            ltout => OPEN,
            carryin => \scaler_1.un3_source_data_0_cry_2\,
            carryout => \scaler_1.un3_source_data_0_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_1.un3_source_data_un3_source_data_0_cry_3_c_RNIO4F11_LC_2_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15033\,
            in2 => \N__10347\,
            in3 => \N__10338\,
            lcout => \scaler_1.un3_source_data_0_cry_3_c_RNIO4F11\,
            ltout => OPEN,
            carryin => \scaler_1.un3_source_data_0_cry_3\,
            carryout => \scaler_1.un3_source_data_0_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_1.un3_source_data_un3_source_data_0_cry_4_c_RNIR8G11_LC_2_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10335\,
            in2 => \N__10326\,
            in3 => \N__10317\,
            lcout => \scaler_1.un3_source_data_0_cry_4_c_RNIR8G11\,
            ltout => OPEN,
            carryin => \scaler_1.un3_source_data_0_cry_4\,
            carryout => \scaler_1.un3_source_data_0_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_1.un3_source_data_un3_source_data_0_cry_5_c_RNIUCH11_LC_2_27_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10548\,
            in2 => \N__10542\,
            in3 => \N__10530\,
            lcout => \scaler_1.un3_source_data_0_cry_5_c_RNIUCH11\,
            ltout => OPEN,
            carryin => \scaler_1.un3_source_data_0_cry_5\,
            carryout => \scaler_1.un3_source_data_0_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_1.un3_source_data_un3_source_data_0_cry_6_c_RNI1HI11_LC_2_27_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__11724\,
            in3 => \N__10527\,
            lcout => \scaler_1.un3_source_data_0_cry_6_c_RNI1HI11\,
            ltout => OPEN,
            carryin => \scaler_1.un3_source_data_0_cry_6\,
            carryout => \scaler_1.un3_source_data_0_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_1.un3_source_data_un3_source_data_0_cry_7_c_RNI2JJ11_LC_2_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10518\,
            in2 => \N__24767\,
            in3 => \N__10524\,
            lcout => \scaler_1.un3_source_data_0_cry_7_c_RNI2JJ11\,
            ltout => OPEN,
            carryin => \bfn_2_28_0_\,
            carryout => \scaler_1.un3_source_data_0_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_1.un3_source_data_un3_source_data_0_cry_8_c_RNIPB6F_LC_2_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10521\,
            lcout => \scaler_1.un3_source_data_0_cry_8_c_RNIPB6F\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_1.N_771_i_l_ofx_LC_2_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11754\,
            in2 => \_gnd_net_\,
            in3 => \N__11739\,
            lcout => \scaler_1.N_771_i_l_ofxZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_1.un2_source_data_0_cry_1_c_RNO_LC_2_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__11435\,
            in1 => \N__11857\,
            in2 => \_gnd_net_\,
            in3 => \N__11402\,
            lcout => \scaler_1.un2_source_data_0_cry_1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.un2_source_data_0_cry_1_c_RNO_LC_2_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__10438\,
            in1 => \N__10504\,
            in2 => \_gnd_net_\,
            in3 => \N__10473\,
            lcout => \scaler_4.un2_source_data_0_cry_1_c_RNO_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.un2_source_data_0_cry_1_c_LC_2_29_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10431\,
            in2 => \N__10449\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_29_0_\,
            carryout => \scaler_4.un2_source_data_0_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.source_data_1_esr_6_LC_2_29_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10661\,
            in2 => \N__10439\,
            in3 => \N__10413\,
            lcout => scaler_4_data_6,
            ltout => OPEN,
            carryin => \scaler_4.un2_source_data_0_cry_1\,
            carryout => \scaler_4.un2_source_data_0_cry_2\,
            clk => \N__23818\,
            ce => \N__11961\,
            sr => \N__23403\
        );

    \scaler_4.source_data_1_esr_7_LC_2_29_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10646\,
            in2 => \N__10665\,
            in3 => \N__10653\,
            lcout => scaler_4_data_7,
            ltout => OPEN,
            carryin => \scaler_4.un2_source_data_0_cry_2\,
            carryout => \scaler_4.un2_source_data_0_cry_3\,
            clk => \N__23818\,
            ce => \N__11961\,
            sr => \N__23403\
        );

    \scaler_4.source_data_1_esr_8_LC_2_29_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10631\,
            in2 => \N__10650\,
            in3 => \N__10638\,
            lcout => scaler_4_data_8,
            ltout => OPEN,
            carryin => \scaler_4.un2_source_data_0_cry_3\,
            carryout => \scaler_4.un2_source_data_0_cry_4\,
            clk => \N__23818\,
            ce => \N__11961\,
            sr => \N__23403\
        );

    \scaler_4.source_data_1_esr_9_LC_2_29_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10616\,
            in2 => \N__10635\,
            in3 => \N__10623\,
            lcout => scaler_4_data_9,
            ltout => OPEN,
            carryin => \scaler_4.un2_source_data_0_cry_4\,
            carryout => \scaler_4.un2_source_data_0_cry_5\,
            clk => \N__23818\,
            ce => \N__11961\,
            sr => \N__23403\
        );

    \scaler_4.source_data_1_esr_10_LC_2_29_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10601\,
            in2 => \N__10620\,
            in3 => \N__10608\,
            lcout => scaler_4_data_10,
            ltout => OPEN,
            carryin => \scaler_4.un2_source_data_0_cry_5\,
            carryout => \scaler_4.un2_source_data_0_cry_6\,
            clk => \N__23818\,
            ce => \N__11961\,
            sr => \N__23403\
        );

    \scaler_4.source_data_1_esr_11_LC_2_29_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10586\,
            in2 => \N__10605\,
            in3 => \N__10593\,
            lcout => scaler_4_data_11,
            ltout => OPEN,
            carryin => \scaler_4.un2_source_data_0_cry_6\,
            carryout => \scaler_4.un2_source_data_0_cry_7\,
            clk => \N__23818\,
            ce => \N__11961\,
            sr => \N__23403\
        );

    \scaler_4.source_data_1_esr_12_LC_2_29_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10574\,
            in2 => \N__10590\,
            in3 => \N__10578\,
            lcout => scaler_4_data_12,
            ltout => OPEN,
            carryin => \scaler_4.un2_source_data_0_cry_7\,
            carryout => \scaler_4.un2_source_data_0_cry_8\,
            clk => \N__23818\,
            ce => \N__11961\,
            sr => \N__23403\
        );

    \scaler_4.source_data_1_esr_13_LC_2_30_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10575\,
            in2 => \N__10563\,
            in3 => \N__10554\,
            lcout => scaler_4_data_13,
            ltout => OPEN,
            carryin => \bfn_2_30_0_\,
            carryout => \scaler_4.un2_source_data_0_cry_9\,
            clk => \N__23812\,
            ce => \N__11959\,
            sr => \N__23405\
        );

    \scaler_4.source_data_1_esr_14_LC_2_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10551\,
            lcout => scaler_4_data_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23812\,
            ce => \N__11959\,
            sr => \N__23405\
        );

    \uart.bit_Count_RNO_0_2_LC_3_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__12921\,
            in1 => \N__12860\,
            in2 => \_gnd_net_\,
            in3 => \N__12032\,
            lcout => \uart.CO1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.state_RNI4ENK_3_LC_3_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__12922\,
            in1 => \N__12861\,
            in2 => \N__12986\,
            in3 => \N__12275\,
            lcout => \uart.N_133_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.bit_Count_RNIETHE_2_LC_3_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__12973\,
            in1 => \N__12918\,
            in2 => \_gnd_net_\,
            in3 => \N__12855\,
            lcout => \uart.N_177\,
            ltout => \uart.N_177_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.timer_Count_RNIBAKE2_6_LC_3_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__14248\,
            in1 => \N__14298\,
            in2 => \N__10683\,
            in3 => \N__12021\,
            lcout => \uart.N_168_1\,
            ltout => \uart.N_168_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.state_3_LC_3_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010001100"
        )
    port map (
            in0 => \N__12087\,
            in1 => \N__10680\,
            in2 => \N__10674\,
            in3 => \N__12147\,
            lcout => \uart.stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23873\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.data_Aux_RNO_0_5_LC_3_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__12858\,
            in1 => \N__12976\,
            in2 => \_gnd_net_\,
            in3 => \N__12925\,
            lcout => \uart.data_Auxce_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.data_Aux_RNO_0_6_LC_3_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__12977\,
            in1 => \N__12920\,
            in2 => \_gnd_net_\,
            in3 => \N__12859\,
            lcout => \uart.data_Auxce_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.data_Aux_RNO_0_0_LC_3_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__12856\,
            in1 => \N__12974\,
            in2 => \_gnd_net_\,
            in3 => \N__12924\,
            lcout => \uart.data_Auxce_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.data_Aux_RNO_0_3_LC_3_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__12975\,
            in1 => \N__12919\,
            in2 => \_gnd_net_\,
            in3 => \N__12857\,
            lcout => \uart.data_Auxce_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.state_RNO_3_3_LC_3_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__12084\,
            in1 => \N__14247\,
            in2 => \_gnd_net_\,
            in3 => \N__14297\,
            lcout => \uart.N_154_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_7_LC_3_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111010101010"
        )
    port map (
            in0 => \N__13416\,
            in1 => \N__10823\,
            in2 => \_gnd_net_\,
            in3 => \N__13237\,
            lcout => \uart_frame_decoder.state_1Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23868\,
            ce => 'H',
            sr => \N__23342\
        );

    \uart.data_rdy_LC_3_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010000000"
        )
    port map (
            in0 => \N__12207\,
            in1 => \N__14250\,
            in2 => \N__12638\,
            in3 => \N__12310\,
            lcout => uart_data_rdy,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23868\,
            ce => 'H',
            sr => \N__23342\
        );

    \uart.data_Aux_0_LC_3_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010111000"
        )
    port map (
            in0 => \N__12627\,
            in1 => \N__10755\,
            in2 => \N__10772\,
            in3 => \N__12113\,
            lcout => \uart.data_AuxZ1Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23864\,
            ce => 'H',
            sr => \N__12321\
        );

    \uart.data_Aux_1_LC_3_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111101000000"
        )
    port map (
            in0 => \N__12114\,
            in1 => \N__12630\,
            in2 => \N__10746\,
            in3 => \N__10889\,
            lcout => \uart.data_AuxZ1Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23864\,
            ce => 'H',
            sr => \N__12321\
        );

    \uart.data_Aux_2_LC_3_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010111000"
        )
    port map (
            in0 => \N__12628\,
            in1 => \N__12822\,
            in2 => \N__11003\,
            in3 => \N__12115\,
            lcout => \uart.data_AuxZ1Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23864\,
            ce => 'H',
            sr => \N__12321\
        );

    \uart.data_Aux_3_LC_3_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011110000"
        )
    port map (
            in0 => \N__12116\,
            in1 => \N__12631\,
            in2 => \N__12563\,
            in3 => \N__10734\,
            lcout => \uart.data_AuxZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23864\,
            ce => 'H',
            sr => \N__12321\
        );

    \uart.data_Aux_4_LC_3_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010111000"
        )
    port map (
            in0 => \N__12629\,
            in1 => \N__12348\,
            in2 => \N__13346\,
            in3 => \N__12117\,
            lcout => \uart.data_AuxZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23864\,
            ce => 'H',
            sr => \N__12321\
        );

    \uart.data_Aux_5_LC_3_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011110000"
        )
    port map (
            in0 => \N__12118\,
            in1 => \N__12632\,
            in2 => \N__11111\,
            in3 => \N__10725\,
            lcout => \uart.data_AuxZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23864\,
            ce => 'H',
            sr => \N__12321\
        );

    \uart.data_Aux_6_LC_3_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011100100"
        )
    port map (
            in0 => \N__10716\,
            in1 => \N__12470\,
            in2 => \N__12639\,
            in3 => \N__12119\,
            lcout => \uart.data_AuxZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23864\,
            ce => 'H',
            sr => \N__12321\
        );

    \uart.data_Aux_7_LC_3_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111101000000"
        )
    port map (
            in0 => \N__12120\,
            in1 => \N__12633\,
            in2 => \N__10875\,
            in3 => \N__10904\,
            lcout => \uart.data_AuxZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23864\,
            ce => 'H',
            sr => \N__12321\
        );

    \uart.state_RNO_0_0_LC_3_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011011101"
        )
    port map (
            in0 => \N__12681\,
            in1 => \N__12626\,
            in2 => \_gnd_net_\,
            in3 => \N__23503\,
            lcout => OPEN,
            ltout => \uart.state_srsts_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.state_0_LC_3_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110001111"
        )
    port map (
            in0 => \N__12208\,
            in1 => \N__14249\,
            in2 => \N__10863\,
            in3 => \N__12312\,
            lcout => \uart.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23859\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_RNI592G_10_LC_3_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13156\,
            in2 => \_gnd_net_\,
            in3 => \N__13090\,
            lcout => \uart_frame_decoder.state_1_RNI592GZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_RNO_3_0_LC_3_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__13157\,
            in1 => \N__11151\,
            in2 => \_gnd_net_\,
            in3 => \N__10793\,
            lcout => \uart_frame_decoder.state_1_RNO_3Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_RNO_0_0_LC_3_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001010"
        )
    port map (
            in0 => \N__10808\,
            in1 => \_gnd_net_\,
            in2 => \N__11161\,
            in3 => \N__13161\,
            lcout => \uart_frame_decoder.N_168_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_RNO_2_0_LC_3_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__13092\,
            in1 => \N__11150\,
            in2 => \N__13168\,
            in3 => \N__10807\,
            lcout => \uart_frame_decoder.state_1_RNO_2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_RNIRN9H_7_LC_3_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10824\,
            in2 => \_gnd_net_\,
            in3 => \N__13091\,
            lcout => \uart_frame_decoder.source_offset2data_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_RNO_0_1_LC_3_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10809\,
            in2 => \_gnd_net_\,
            in3 => \N__10794\,
            lcout => \uart_frame_decoder.state_1_ns_0_i_a2_0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.data_0_LC_3_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__11212\,
            in1 => \N__10773\,
            in2 => \_gnd_net_\,
            in3 => \N__13382\,
            lcout => uart_data_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23854\,
            ce => 'H',
            sr => \N__13329\
        );

    \uart_frame_decoder.state_1_ns_0_i_a2_0_0_1_2_LC_3_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11045\,
            in2 => \_gnd_net_\,
            in3 => \N__11211\,
            lcout => OPEN,
            ltout => \uart_frame_decoder.state_1_ns_0_i_a2_0_0_1Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_RNI12LB1_1_LC_3_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__11166\,
            in1 => \N__11544\,
            in2 => \N__11130\,
            in3 => \N__10943\,
            lcout => \uart_frame_decoder.state_1_ns_0_i_a2_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.data_5_LC_3_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__13385\,
            in1 => \N__11112\,
            in2 => \_gnd_net_\,
            in3 => \N__11046\,
            lcout => uart_data_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23854\,
            ce => 'H',
            sr => \N__13329\
        );

    \uart.data_2_LC_3_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__11007\,
            in1 => \N__10944\,
            in2 => \_gnd_net_\,
            in3 => \N__13384\,
            lcout => uart_data_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23854\,
            ce => 'H',
            sr => \N__13329\
        );

    \uart.data_7_LC_3_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__13386\,
            in1 => \_gnd_net_\,
            in2 => \N__11570\,
            in3 => \N__10908\,
            lcout => uart_data_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23854\,
            ce => 'H',
            sr => \N__13329\
        );

    \uart.data_1_LC_3_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__10893\,
            in1 => \N__12740\,
            in2 => \_gnd_net_\,
            in3 => \N__13383\,
            lcout => uart_data_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23854\,
            ce => 'H',
            sr => \N__13329\
        );

    \scaler_2.un2_source_data_0_cry_1_c_LC_3_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14598\,
            in2 => \N__14580\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_3_21_0_\,
            carryout => \scaler_2.un2_source_data_0_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_2.source_data_1_esr_6_LC_3_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11366\,
            in2 => \N__14606\,
            in3 => \N__10878\,
            lcout => scaler_2_data_6,
            ltout => OPEN,
            carryin => \scaler_2.un2_source_data_0_cry_1\,
            carryout => \scaler_2.un2_source_data_0_cry_2\,
            clk => \N__23850\,
            ce => \N__11967\,
            sr => \N__23353\
        );

    \scaler_2.source_data_1_esr_7_LC_3_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11351\,
            in2 => \N__11370\,
            in3 => \N__11358\,
            lcout => scaler_2_data_7,
            ltout => OPEN,
            carryin => \scaler_2.un2_source_data_0_cry_2\,
            carryout => \scaler_2.un2_source_data_0_cry_3\,
            clk => \N__23850\,
            ce => \N__11967\,
            sr => \N__23353\
        );

    \scaler_2.source_data_1_esr_8_LC_3_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11336\,
            in2 => \N__11355\,
            in3 => \N__11343\,
            lcout => scaler_2_data_8,
            ltout => OPEN,
            carryin => \scaler_2.un2_source_data_0_cry_3\,
            carryout => \scaler_2.un2_source_data_0_cry_4\,
            clk => \N__23850\,
            ce => \N__11967\,
            sr => \N__23353\
        );

    \scaler_2.source_data_1_esr_9_LC_3_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11321\,
            in2 => \N__11340\,
            in3 => \N__11328\,
            lcout => scaler_2_data_9,
            ltout => OPEN,
            carryin => \scaler_2.un2_source_data_0_cry_4\,
            carryout => \scaler_2.un2_source_data_0_cry_5\,
            clk => \N__23850\,
            ce => \N__11967\,
            sr => \N__23353\
        );

    \scaler_2.source_data_1_esr_10_LC_3_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11306\,
            in2 => \N__11325\,
            in3 => \N__11313\,
            lcout => scaler_2_data_10,
            ltout => OPEN,
            carryin => \scaler_2.un2_source_data_0_cry_5\,
            carryout => \scaler_2.un2_source_data_0_cry_6\,
            clk => \N__23850\,
            ce => \N__11967\,
            sr => \N__23353\
        );

    \scaler_2.source_data_1_esr_11_LC_3_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11291\,
            in2 => \N__11310\,
            in3 => \N__11298\,
            lcout => scaler_2_data_11,
            ltout => OPEN,
            carryin => \scaler_2.un2_source_data_0_cry_6\,
            carryout => \scaler_2.un2_source_data_0_cry_7\,
            clk => \N__23850\,
            ce => \N__11967\,
            sr => \N__23353\
        );

    \scaler_2.source_data_1_esr_12_LC_3_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11279\,
            in2 => \N__11295\,
            in3 => \N__11283\,
            lcout => scaler_2_data_12,
            ltout => OPEN,
            carryin => \scaler_2.un2_source_data_0_cry_7\,
            carryout => \scaler_2.un2_source_data_0_cry_8\,
            clk => \N__23850\,
            ce => \N__11967\,
            sr => \N__23353\
        );

    \scaler_2.source_data_1_esr_13_LC_3_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11280\,
            in2 => \N__11268\,
            in3 => \N__11259\,
            lcout => scaler_2_data_13,
            ltout => OPEN,
            carryin => \bfn_3_22_0_\,
            carryout => \scaler_2.un2_source_data_0_cry_9\,
            clk => \N__23848\,
            ce => \N__11966\,
            sr => \N__23359\
        );

    \scaler_2.source_data_1_esr_14_LC_3_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11256\,
            lcout => scaler_2_data_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23848\,
            ce => \N__11966\,
            sr => \N__23359\
        );

    \scaler_2.source_data_1_esr_5_LC_3_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__15229\,
            in1 => \N__14602\,
            in2 => \_gnd_net_\,
            in3 => \N__15194\,
            lcout => scaler_2_data_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23848\,
            ce => \N__11966\,
            sr => \N__23359\
        );

    \scaler_3.source_data_1_esr_5_LC_3_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__13505\,
            in1 => \N__11691\,
            in2 => \_gnd_net_\,
            in3 => \N__13473\,
            lcout => scaler_3_data_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23848\,
            ce => \N__11966\,
            sr => \N__23359\
        );

    \uart_frame_decoder.state_1_8_LC_3_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__11636\,
            in1 => \N__11658\,
            in2 => \_gnd_net_\,
            in3 => \N__13265\,
            lcout => \uart_frame_decoder.state_1Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23845\,
            ce => 'H',
            sr => \N__23363\
        );

    \uart_frame_decoder.state_1_9_LC_3_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110100000"
        )
    port map (
            in0 => \N__13266\,
            in1 => \_gnd_net_\,
            in2 => \N__11616\,
            in3 => \N__11622\,
            lcout => \uart_frame_decoder.state_1Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23845\,
            ce => 'H',
            sr => \N__23363\
        );

    \uart_frame_decoder.state_1_RNITP9H_9_LC_3_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11612\,
            in2 => \_gnd_net_\,
            in3 => \N__13106\,
            lcout => \uart_frame_decoder.source_offset4data_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_5_LC_3_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__11604\,
            in1 => \N__11463\,
            in2 => \_gnd_net_\,
            in3 => \N__13263\,
            lcout => \uart_frame_decoder.state_1Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23845\,
            ce => 'H',
            sr => \N__23363\
        );

    \uart_frame_decoder.state_1_6_LC_3_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__13264\,
            in1 => \N__11592\,
            in2 => \_gnd_net_\,
            in3 => \N__13430\,
            lcout => \uart_frame_decoder.state_1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23845\,
            ce => 'H',
            sr => \N__23363\
        );

    \uart_frame_decoder.source_CH4data_esr_7_LC_3_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11583\,
            lcout => \frame_decoder_CH4data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23839\,
            ce => \N__11477\,
            sr => \N__23368\
        );

    \uart_frame_decoder.state_1_RNIL1GQ_4_LC_3_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11459\,
            in2 => \_gnd_net_\,
            in3 => \N__23502\,
            lcout => \uart_frame_decoder.source_CH3data_1_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_1.source_data_1_esr_5_LC_3_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__11859\,
            in1 => \N__11430\,
            in2 => \_gnd_net_\,
            in3 => \N__11394\,
            lcout => scaler_1_data_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23834\,
            ce => \N__11963\,
            sr => \N__23375\
        );

    \scaler_1.un3_source_data_un3_source_data_0_axb_7_LC_3_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11750\,
            in2 => \_gnd_net_\,
            in3 => \N__11735\,
            lcout => \scaler_1.un3_source_data_0_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_rudder_cry_6_c_LC_3_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13526\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_3_26_0_\,
            carryout => \ppm_encoder_1.un1_rudder_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_rudder_cry_6_THRU_LUT4_0_LC_3_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16613\,
            in2 => \_gnd_net_\,
            in3 => \N__11712\,
            lcout => \ppm_encoder_1.un1_rudder_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_rudder_cry_6\,
            carryout => \ppm_encoder_1.un1_rudder_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_rudder_cry_7_THRU_LUT4_0_LC_3_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16688\,
            in2 => \_gnd_net_\,
            in3 => \N__11709\,
            lcout => \ppm_encoder_1.un1_rudder_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_rudder_cry_7\,
            carryout => \ppm_encoder_1.un1_rudder_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_rudder_cry_8_THRU_LUT4_0_LC_3_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15284\,
            in2 => \_gnd_net_\,
            in3 => \N__11706\,
            lcout => \ppm_encoder_1.un1_rudder_cry_8_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_rudder_cry_8\,
            carryout => \ppm_encoder_1.un1_rudder_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_rudder_cry_9_THRU_LUT4_0_LC_3_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13616\,
            in3 => \N__11703\,
            lcout => \ppm_encoder_1.un1_rudder_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_rudder_cry_9\,
            carryout => \ppm_encoder_1.un1_rudder_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_rudder_cry_10_THRU_LUT4_0_LC_3_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13208\,
            in2 => \_gnd_net_\,
            in3 => \N__11700\,
            lcout => \ppm_encoder_1.un1_rudder_cry_10_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_rudder_cry_10\,
            carryout => \ppm_encoder_1.un1_rudder_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_rudder_cry_11_THRU_LUT4_0_LC_3_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15134\,
            in2 => \_gnd_net_\,
            in3 => \N__11697\,
            lcout => \ppm_encoder_1.un1_rudder_cry_11_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_rudder_cry_11\,
            carryout => \ppm_encoder_1.un1_rudder_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_rudder_cry_12_THRU_LUT4_0_LC_3_26_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13559\,
            in2 => \N__24771\,
            in3 => \N__11694\,
            lcout => \ppm_encoder_1.un1_rudder_cry_12_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_rudder_cry_12\,
            carryout => \ppm_encoder_1.un1_rudder_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.rudder_esr_14_LC_3_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11880\,
            in2 => \_gnd_net_\,
            in3 => \N__11871\,
            lcout => \ppm_encoder_1.rudderZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23823\,
            ce => \N__16261\,
            sr => \N__23390\
        );

    \scaler_1.un2_source_data_0_cry_1_c_LC_3_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11850\,
            in2 => \N__11868\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_3_28_0_\,
            carryout => \scaler_1.un2_source_data_0_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_1.source_data_1_esr_6_LC_3_28_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11825\,
            in2 => \N__11858\,
            in3 => \N__11832\,
            lcout => scaler_1_data_6,
            ltout => OPEN,
            carryin => \scaler_1.un2_source_data_0_cry_1\,
            carryout => \scaler_1.un2_source_data_0_cry_2\,
            clk => \N__23819\,
            ce => \N__11962\,
            sr => \N__23395\
        );

    \scaler_1.source_data_1_esr_7_LC_3_28_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11810\,
            in2 => \N__11829\,
            in3 => \N__11817\,
            lcout => scaler_1_data_7,
            ltout => OPEN,
            carryin => \scaler_1.un2_source_data_0_cry_2\,
            carryout => \scaler_1.un2_source_data_0_cry_3\,
            clk => \N__23819\,
            ce => \N__11962\,
            sr => \N__23395\
        );

    \scaler_1.source_data_1_esr_8_LC_3_28_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11795\,
            in2 => \N__11814\,
            in3 => \N__11802\,
            lcout => scaler_1_data_8,
            ltout => OPEN,
            carryin => \scaler_1.un2_source_data_0_cry_3\,
            carryout => \scaler_1.un2_source_data_0_cry_4\,
            clk => \N__23819\,
            ce => \N__11962\,
            sr => \N__23395\
        );

    \scaler_1.source_data_1_esr_9_LC_3_28_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11780\,
            in2 => \N__11799\,
            in3 => \N__11787\,
            lcout => scaler_1_data_9,
            ltout => OPEN,
            carryin => \scaler_1.un2_source_data_0_cry_4\,
            carryout => \scaler_1.un2_source_data_0_cry_5\,
            clk => \N__23819\,
            ce => \N__11962\,
            sr => \N__23395\
        );

    \scaler_1.source_data_1_esr_10_LC_3_28_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11765\,
            in2 => \N__11784\,
            in3 => \N__11772\,
            lcout => scaler_1_data_10,
            ltout => OPEN,
            carryin => \scaler_1.un2_source_data_0_cry_5\,
            carryout => \scaler_1.un2_source_data_0_cry_6\,
            clk => \N__23819\,
            ce => \N__11962\,
            sr => \N__23395\
        );

    \scaler_1.source_data_1_esr_11_LC_3_28_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12005\,
            in2 => \N__11769\,
            in3 => \N__11757\,
            lcout => scaler_1_data_11,
            ltout => OPEN,
            carryin => \scaler_1.un2_source_data_0_cry_6\,
            carryout => \scaler_1.un2_source_data_0_cry_7\,
            clk => \N__23819\,
            ce => \N__11962\,
            sr => \N__23395\
        );

    \scaler_1.source_data_1_esr_12_LC_3_28_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11993\,
            in2 => \N__12009\,
            in3 => \N__11997\,
            lcout => scaler_1_data_12,
            ltout => OPEN,
            carryin => \scaler_1.un2_source_data_0_cry_7\,
            carryout => \scaler_1.un2_source_data_0_cry_8\,
            clk => \N__23819\,
            ce => \N__11962\,
            sr => \N__23395\
        );

    \scaler_1.source_data_1_esr_13_LC_3_29_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11994\,
            in2 => \N__11982\,
            in3 => \N__11973\,
            lcout => scaler_1_data_13,
            ltout => OPEN,
            carryin => \bfn_3_29_0_\,
            carryout => \scaler_1.un2_source_data_0_cry_9\,
            clk => \N__23813\,
            ce => \N__11960\,
            sr => \N__23399\
        );

    \scaler_1.source_data_1_esr_14_LC_3_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11970\,
            lcout => scaler_1_data_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23813\,
            ce => \N__11960\,
            sr => \N__23399\
        );

    \uart_frame_decoder.source_offset3data_esr_1_LC_3_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12792\,
            lcout => \frame_decoder_OFF3data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23808\,
            ce => \N__11916\,
            sr => \N__23404\
        );

    \uart_sync.aux_2__0__0_LC_4_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13980\,
            lcout => \uart_sync.aux_2__0_Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23881\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_sync.aux_3__0__0_LC_4_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11895\,
            lcout => \uart_sync.aux_3__0_Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23880\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.timer_Count_1_LC_4_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14143\,
            in2 => \_gnd_net_\,
            in3 => \N__13972\,
            lcout => \uart.timer_CountZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23879\,
            ce => 'H',
            sr => \N__14183\
        );

    \uart.state_RNO_0_2_LC_4_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010111011"
        )
    port map (
            in0 => \N__12595\,
            in1 => \N__12659\,
            in2 => \_gnd_net_\,
            in3 => \N__12086\,
            lcout => \uart.N_151\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_sync.Q_0__0_LC_4_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11889\,
            lcout => uart_input_sync,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23876\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.state_RNIB0BC_2_LC_4_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12085\,
            in2 => \_gnd_net_\,
            in3 => \N__12273\,
            lcout => \uart.N_159\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.state_2_LC_4_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001010001"
        )
    port map (
            in0 => \N__12093\,
            in1 => \N__12054\,
            in2 => \N__12666\,
            in3 => \N__24463\,
            lcout => \uart.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23874\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.state_RNIGITG2_0_4_LC_4_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010000"
        )
    port map (
            in0 => \N__14218\,
            in1 => \_gnd_net_\,
            in2 => \N__12216\,
            in3 => \N__12309\,
            lcout => OPEN,
            ltout => \uart.timer_Count_0_sqmuxa_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.state_RNILCH65_2_LC_4_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001110"
        )
    port map (
            in0 => \N__12063\,
            in1 => \N__12053\,
            in2 => \N__12057\,
            in3 => \N__24462\,
            lcout => \uart.timer_Count_1_sqmuxa_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.timer_Count_RNITC202_6_LC_4_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__14217\,
            in1 => \N__14279\,
            in2 => \_gnd_net_\,
            in3 => \N__12020\,
            lcout => \uart.N_180\,
            ltout => \uart.N_180_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.state_RNIAFDC2_3_LC_4_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110101"
        )
    port map (
            in0 => \N__12272\,
            in1 => \_gnd_net_\,
            in2 => \N__12045\,
            in3 => \N__12209\,
            lcout => \uart.un1_state_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.timer_Count_RNINU001_1_LC_4_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__13948\,
            in1 => \_gnd_net_\,
            in2 => \N__13926\,
            in3 => \N__13973\,
            lcout => \uart.N_146_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.timer_Count_RNIQPMA1_2_LC_4_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100001111"
        )
    port map (
            in0 => \N__14114\,
            in1 => \N__13920\,
            in2 => \N__14328\,
            in3 => \N__13947\,
            lcout => \uart.N_143_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_RNO_0_1_LC_4_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14081\,
            in2 => \_gnd_net_\,
            in3 => \N__14056\,
            lcout => OPEN,
            ltout => \reset_module_System.count_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_1_LC_4_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__12365\,
            in1 => \N__14647\,
            in2 => \N__12156\,
            in3 => \N__12342\,
            lcout => \reset_module_System.countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23869\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.timer_Count_RNIICSG1_5_LC_4_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__14326\,
            in1 => \N__12213\,
            in2 => \N__14291\,
            in3 => \N__14091\,
            lcout => \uart.un1_state_2_0_a3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.reset_LC_4_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__12364\,
            in1 => \N__14646\,
            in2 => \_gnd_net_\,
            in3 => \N__12341\,
            lcout => reset_system,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23869\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.timer_Count_RNIN6202_4_LC_4_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010000000"
        )
    port map (
            in0 => \N__14324\,
            in1 => \N__12131\,
            in2 => \N__14290\,
            in3 => \N__14115\,
            lcout => \uart.N_153_0\,
            ltout => \uart.N_153_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.state_RNO_0_4_LC_4_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__12214\,
            in1 => \N__24467\,
            in2 => \N__12153\,
            in3 => \N__14227\,
            lcout => \uart.N_167\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.state_RNO_2_3_LC_4_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__14325\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12274\,
            lcout => OPEN,
            ltout => \uart.state_srsts_i_a3_0_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.state_RNO_0_3_LC_4_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__14116\,
            in1 => \N__13925\,
            in2 => \N__12150\,
            in3 => \N__13950\,
            lcout => \uart.N_170\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.state_RNIMD8T2_3_LC_4_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001011111010"
        )
    port map (
            in0 => \N__12276\,
            in1 => \N__12141\,
            in2 => \N__12215\,
            in3 => \N__12135\,
            lcout => \uart.un1_state_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_2_LC_4_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010101010101010"
        )
    port map (
            in0 => \N__14022\,
            in1 => \N__12340\,
            in2 => \N__14652\,
            in3 => \N__12366\,
            lcout => \reset_module_System.countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23865\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_RNI97FD_5_LC_4_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__14408\,
            in1 => \N__14423\,
            in2 => \N__14394\,
            in3 => \N__14453\,
            lcout => \reset_module_System.reset6_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_RNI9O1P_2_LC_4_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__14012\,
            in1 => \N__14438\,
            in2 => \N__14490\,
            in3 => \N__14033\,
            lcout => OPEN,
            ltout => \reset_module_System.reset6_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_RNIN3HK3_12_LC_4_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__14346\,
            in1 => \N__14080\,
            in2 => \N__12369\,
            in3 => \N__12801\,
            lcout => \reset_module_System.reset6_19\,
            ltout => \reset_module_System.reset6_19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_0_LC_4_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011001100110011"
        )
    port map (
            in0 => \N__14648\,
            in1 => \N__14085\,
            in2 => \N__12351\,
            in3 => \N__12339\,
            lcout => \reset_module_System.countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23865\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_RNIP8RT_10_LC_4_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__14375\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14360\,
            lcout => \reset_module_System.reset6_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.data_Aux_RNO_0_4_LC_4_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000000"
        )
    port map (
            in0 => \N__12879\,
            in1 => \_gnd_net_\,
            in2 => \N__12939\,
            in3 => \N__12993\,
            lcout => \uart.data_Auxce_0_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_RNI10J41_1_LC_4_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__14469\,
            in1 => \N__14547\,
            in2 => \N__14514\,
            in3 => \N__14058\,
            lcout => \reset_module_System.reset6_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.state_RNIAFHL_3_LC_4_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100010001"
        )
    port map (
            in0 => \N__12206\,
            in1 => \N__12284\,
            in2 => \_gnd_net_\,
            in3 => \N__23500\,
            lcout => \uart.state_RNIAFHLZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.state_RNIGITG2_4_LC_4_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__12202\,
            in1 => \N__14240\,
            in2 => \_gnd_net_\,
            in3 => \N__12311\,
            lcout => \uart.data_rdyc_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.state_4_LC_4_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100100000"
        )
    port map (
            in0 => \N__12285\,
            in1 => \N__24487\,
            in2 => \N__12237\,
            in3 => \N__12225\,
            lcout => \uart.stateZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23860\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.data_Aux_RNO_0_2_LC_4_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__12992\,
            in1 => \N__12935\,
            in2 => \_gnd_net_\,
            in3 => \N__12878\,
            lcout => \uart.data_Auxce_0_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_RNI53692_14_LC_4_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__14564\,
            in1 => \N__12816\,
            in2 => \N__14532\,
            in3 => \N__12807\,
            lcout => \reset_module_System.reset6_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_ns_0_i_a2_1_1_2_LC_4_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__12495\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12397\,
            lcout => OPEN,
            ltout => \uart_frame_decoder.state_1_ns_0_i_a2_1_1Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_ns_0_i_a2_1_2_LC_4_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__15056\,
            in1 => \N__12739\,
            in2 => \N__12711\,
            in3 => \N__13099\,
            lcout => \uart_frame_decoder.state_1_ns_0_i_a2_1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.state_1_LC_4_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100000"
        )
    port map (
            in0 => \N__12680\,
            in1 => \N__12658\,
            in2 => \N__12637\,
            in3 => \N__23530\,
            lcout => \uart.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23855\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.state_RNIQABT2_4_LC_4_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111001100"
        )
    port map (
            in0 => \N__12599\,
            in1 => \N__24500\,
            in2 => \_gnd_net_\,
            in3 => \N__13360\,
            lcout => \uart.state_RNIQABT2Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.data_3_LC_4_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__12564\,
            in1 => \N__12496\,
            in2 => \_gnd_net_\,
            in3 => \N__13379\,
            lcout => uart_data_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23851\,
            ce => 'H',
            sr => \N__13325\
        );

    \uart.data_6_LC_4_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__12477\,
            in1 => \N__12398\,
            in2 => \_gnd_net_\,
            in3 => \N__13381\,
            lcout => uart_data_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23851\,
            ce => 'H',
            sr => \N__13325\
        );

    \uart_frame_decoder.state_1_RNIQM9H_6_LC_4_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__13434\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13093\,
            lcout => \uart_frame_decoder.source_offset1data_1_sqmuxa\,
            ltout => \uart_frame_decoder.source_offset1data_1_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_frame_decoder.state_1_RNIN3GQ_6_LC_4_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13404\,
            in3 => \N__23497\,
            lcout => \uart_frame_decoder.source_offset1data_1_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.data_4_LC_4_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__13380\,
            in1 => \N__13347\,
            in2 => \_gnd_net_\,
            in3 => \N__15057\,
            lcout => uart_data_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23851\,
            ce => 'H',
            sr => \N__13325\
        );

    \scaler_1.source_data_valid_LC_4_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__14916\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => scaler_1_dv,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23849\,
            ce => 'H',
            sr => \N__23349\
        );

    \uart_frame_decoder.state_1_10_LC_4_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__13154\,
            in1 => \N__13308\,
            in2 => \N__13290\,
            in3 => \N__13253\,
            lcout => \uart_frame_decoder.state_1Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23849\,
            ce => 'H',
            sr => \N__23349\
        );

    \ppm_encoder_1.rudder_11_LC_4_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__13209\,
            in1 => \N__13185\,
            in2 => \N__17460\,
            in3 => \N__18406\,
            lcout => \ppm_encoder_1.rudderZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23849\,
            ce => 'H',
            sr => \N__23349\
        );

    \uart_frame_decoder.source_data_valid_LC_4_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000011001000"
        )
    port map (
            in0 => \N__13155\,
            in1 => \N__13117\,
            in2 => \N__14932\,
            in3 => \N__13011\,
            lcout => frame_decoder_dv_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23849\,
            ce => 'H',
            sr => \N__23349\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_9_LC_4_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110001000100"
        )
    port map (
            in0 => \N__15315\,
            in1 => \N__20256\,
            in2 => \N__14865\,
            in3 => \N__20151\,
            lcout => \ppm_encoder_1.N_325\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_7_LC_4_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__13749\,
            in1 => \N__13728\,
            in2 => \N__17461\,
            in3 => \N__17147\,
            lcout => \ppm_encoder_1.elevatorZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23846\,
            ce => 'H',
            sr => \N__23354\
        );

    \ppm_encoder_1.aileron_11_LC_4_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0111001011011000"
        )
    port map (
            in0 => \N__17435\,
            in1 => \N__13656\,
            in2 => \N__19405\,
            in3 => \N__13674\,
            lcout => \ppm_encoder_1.aileronZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23840\,
            ce => 'H',
            sr => \N__23360\
        );

    \ppm_encoder_1.throttle_6_LC_4_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0111011100100010"
        )
    port map (
            in0 => \N__17434\,
            in1 => \N__13848\,
            in2 => \_gnd_net_\,
            in3 => \N__15371\,
            lcout => \ppm_encoder_1.throttleZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23840\,
            ce => 'H',
            sr => \N__23360\
        );

    \ppm_encoder_1.rudder_6_LC_4_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0111011100100010"
        )
    port map (
            in0 => \N__17433\,
            in1 => \N__13533\,
            in2 => \_gnd_net_\,
            in3 => \N__19235\,
            lcout => \ppm_encoder_1.rudderZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23840\,
            ce => 'H',
            sr => \N__23360\
        );

    \scaler_3.source_data_1_4_LC_4_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001011011000"
        )
    port map (
            in0 => \N__14933\,
            in1 => \N__13509\,
            in2 => \N__14624\,
            in3 => \N__13472\,
            lcout => scaler_3_data_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23840\,
            ce => 'H',
            sr => \N__23360\
        );

    \ppm_encoder_1.elevator_6_LC_4_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0111011100100010"
        )
    port map (
            in0 => \N__17432\,
            in1 => \N__13770\,
            in2 => \_gnd_net_\,
            in3 => \N__14735\,
            lcout => \ppm_encoder_1.elevatorZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23840\,
            ce => 'H',
            sr => \N__23360\
        );

    \ppm_encoder_1.un1_aileron_cry_6_c_LC_4_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14765\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_24_0_\,
            carryout => \ppm_encoder_1.un1_aileron_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_aileron_cry_6_THRU_LUT4_0_LC_4_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17105\,
            in2 => \_gnd_net_\,
            in3 => \N__13443\,
            lcout => \ppm_encoder_1.un1_aileron_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_aileron_cry_6\,
            carryout => \ppm_encoder_1.un1_aileron_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_aileron_cry_7_THRU_LUT4_0_LC_4_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15929\,
            in2 => \_gnd_net_\,
            in3 => \N__13440\,
            lcout => \ppm_encoder_1.un1_aileron_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_aileron_cry_7\,
            carryout => \ppm_encoder_1.un1_aileron_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_aileron_cry_8_THRU_LUT4_0_LC_4_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14810\,
            in2 => \_gnd_net_\,
            in3 => \N__13437\,
            lcout => \ppm_encoder_1.un1_aileron_cry_8_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_aileron_cry_8\,
            carryout => \ppm_encoder_1.un1_aileron_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_aileron_cry_9_THRU_LUT4_0_LC_4_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13589\,
            in2 => \_gnd_net_\,
            in3 => \N__13677\,
            lcout => \ppm_encoder_1.un1_aileron_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_aileron_cry_9\,
            carryout => \ppm_encoder_1.un1_aileron_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_aileron_cry_10_THRU_LUT4_0_LC_4_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13673\,
            in2 => \_gnd_net_\,
            in3 => \N__13650\,
            lcout => \ppm_encoder_1.un1_aileron_cry_10_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_aileron_cry_10\,
            carryout => \ppm_encoder_1.un1_aileron_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_aileron_cry_11_THRU_LUT4_0_LC_4_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__15992\,
            in3 => \N__13647\,
            lcout => \ppm_encoder_1.un1_aileron_cry_11_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_aileron_cry_11\,
            carryout => \ppm_encoder_1.un1_aileron_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_aileron_cry_12_THRU_LUT4_0_LC_4_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15839\,
            in2 => \N__24757\,
            in3 => \N__13644\,
            lcout => \ppm_encoder_1.un1_aileron_cry_12_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_aileron_cry_12\,
            carryout => \ppm_encoder_1.un1_aileron_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_esr_14_LC_4_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13641\,
            in2 => \_gnd_net_\,
            in3 => \N__13629\,
            lcout => \ppm_encoder_1.aileronZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23829\,
            ce => \N__16253\,
            sr => \N__23369\
        );

    \ppm_encoder_1.throttle_10_LC_4_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011110000"
        )
    port map (
            in0 => \N__13782\,
            in1 => \N__13797\,
            in2 => \N__19958\,
            in3 => \N__17486\,
            lcout => \ppm_encoder_1.throttleZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23824\,
            ce => 'H',
            sr => \N__23376\
        );

    \ppm_encoder_1.rudder_10_LC_4_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011110000"
        )
    port map (
            in0 => \N__13626\,
            in1 => \N__13620\,
            in2 => \N__19931\,
            in3 => \N__17484\,
            lcout => \ppm_encoder_1.rudderZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23824\,
            ce => 'H',
            sr => \N__23376\
        );

    \ppm_encoder_1.aileron_10_LC_4_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__13593\,
            in1 => \N__13572\,
            in2 => \N__17529\,
            in3 => \N__15649\,
            lcout => \ppm_encoder_1.aileronZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23824\,
            ce => 'H',
            sr => \N__23376\
        );

    \ppm_encoder_1.rudder_13_LC_4_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1001100111110000"
        )
    port map (
            in0 => \N__13563\,
            in1 => \N__13539\,
            in2 => \N__20663\,
            in3 => \N__17485\,
            lcout => \ppm_encoder_1.rudderZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23824\,
            ce => 'H',
            sr => \N__23376\
        );

    \ppm_encoder_1.elevator_12_LC_4_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__13875\,
            in1 => \N__13899\,
            in2 => \N__17530\,
            in3 => \N__19036\,
            lcout => \ppm_encoder_1.elevatorZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23824\,
            ce => 'H',
            sr => \N__23376\
        );

    \ppm_encoder_1.elevator_9_LC_4_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011110000"
        )
    port map (
            in0 => \N__13692\,
            in1 => \N__13713\,
            in2 => \N__14864\,
            in3 => \N__17483\,
            lcout => \ppm_encoder_1.elevatorZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23824\,
            ce => 'H',
            sr => \N__23376\
        );

    \ppm_encoder_1.throttle_9_LC_4_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001011011000"
        )
    port map (
            in0 => \N__17476\,
            in1 => \N__13824\,
            in2 => \N__19010\,
            in3 => \N__13809\,
            lcout => \ppm_encoder_1.throttleZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23824\,
            ce => 'H',
            sr => \N__23376\
        );

    \ppm_encoder_1.un1_elevator_cry_6_c_LC_4_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13769\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_27_0_\,
            carryout => \ppm_encoder_1.un1_elevator_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_elevator_cry_6_THRU_LUT4_0_LC_4_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13748\,
            in2 => \_gnd_net_\,
            in3 => \N__13719\,
            lcout => \ppm_encoder_1.un1_elevator_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_elevator_cry_6\,
            carryout => \ppm_encoder_1.un1_elevator_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_elevator_cry_7_THRU_LUT4_0_LC_4_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16133\,
            in2 => \_gnd_net_\,
            in3 => \N__13716\,
            lcout => \ppm_encoder_1.un1_elevator_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_elevator_cry_7\,
            carryout => \ppm_encoder_1.un1_elevator_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_elevator_cry_8_THRU_LUT4_0_LC_4_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13709\,
            in2 => \_gnd_net_\,
            in3 => \N__13686\,
            lcout => \ppm_encoder_1.un1_elevator_cry_8_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_elevator_cry_8\,
            carryout => \ppm_encoder_1.un1_elevator_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_elevator_cry_9_THRU_LUT4_0_LC_4_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15266\,
            in2 => \_gnd_net_\,
            in3 => \N__13683\,
            lcout => \ppm_encoder_1.un1_elevator_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_elevator_cry_9\,
            carryout => \ppm_encoder_1.un1_elevator_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_elevator_cry_10_THRU_LUT4_0_LC_4_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15716\,
            in2 => \_gnd_net_\,
            in3 => \N__13680\,
            lcout => \ppm_encoder_1.un1_elevator_cry_10_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_elevator_cry_10\,
            carryout => \ppm_encoder_1.un1_elevator_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_elevator_cry_11_THRU_LUT4_0_LC_4_27_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13898\,
            in2 => \_gnd_net_\,
            in3 => \N__13869\,
            lcout => \ppm_encoder_1.un1_elevator_cry_11_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_elevator_cry_11\,
            carryout => \ppm_encoder_1.un1_elevator_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_elevator_cry_12_THRU_LUT4_0_LC_4_27_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15776\,
            in2 => \N__24769\,
            in3 => \N__13866\,
            lcout => \ppm_encoder_1.un1_elevator_cry_12_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_elevator_cry_12\,
            carryout => \ppm_encoder_1.un1_elevator_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_esr_14_LC_4_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13863\,
            in2 => \_gnd_net_\,
            in3 => \N__13851\,
            lcout => \ppm_encoder_1.elevatorZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23814\,
            ce => \N__16266\,
            sr => \N__23391\
        );

    \ppm_encoder_1.un1_throttle_cry_6_c_LC_4_29_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13841\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_29_0_\,
            carryout => \ppm_encoder_1.un1_throttle_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_throttle_cry_6_THRU_LUT4_0_LC_4_29_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16649\,
            in2 => \_gnd_net_\,
            in3 => \N__13830\,
            lcout => \ppm_encoder_1.un1_throttle_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_throttle_cry_6\,
            carryout => \ppm_encoder_1.un1_throttle_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_throttle_cry_7_THRU_LUT4_0_LC_4_29_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15878\,
            in2 => \_gnd_net_\,
            in3 => \N__13827\,
            lcout => \ppm_encoder_1.un1_throttle_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_throttle_cry_7\,
            carryout => \ppm_encoder_1.un1_throttle_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_throttle_cry_8_THRU_LUT4_0_LC_4_29_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13820\,
            in2 => \_gnd_net_\,
            in3 => \N__13800\,
            lcout => \ppm_encoder_1.un1_throttle_cry_8_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_throttle_cry_8\,
            carryout => \ppm_encoder_1.un1_throttle_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_throttle_cry_9_THRU_LUT4_0_LC_4_29_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13793\,
            in2 => \_gnd_net_\,
            in3 => \N__13773\,
            lcout => \ppm_encoder_1.un1_throttle_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_throttle_cry_9\,
            carryout => \ppm_encoder_1.un1_throttle_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_throttle_cry_10_THRU_LUT4_0_LC_4_29_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16016\,
            in2 => \_gnd_net_\,
            in3 => \N__13998\,
            lcout => \ppm_encoder_1.un1_throttle_cry_10_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_throttle_cry_10\,
            carryout => \ppm_encoder_1.un1_throttle_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_throttle_cry_11_THRU_LUT4_0_LC_4_29_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14990\,
            in2 => \_gnd_net_\,
            in3 => \N__13995\,
            lcout => \ppm_encoder_1.un1_throttle_cry_11_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_throttle_cry_11\,
            carryout => \ppm_encoder_1.un1_throttle_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_throttle_cry_12_THRU_LUT4_0_LC_4_29_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14972\,
            in2 => \N__24770\,
            in3 => \N__13992\,
            lcout => \ppm_encoder_1.un1_throttle_cry_12_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_throttle_cry_12\,
            carryout => \ppm_encoder_1.un1_throttle_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_esr_14_LC_4_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13989\,
            in2 => \_gnd_net_\,
            in3 => \N__13983\,
            lcout => \ppm_encoder_1.throttleZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23802\,
            ce => \N__16262\,
            sr => \N__23400\
        );

    \uart_sync.aux_1__0__0_LC_5_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15387\,
            lcout => \uart_sync.aux_1__0_Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23882\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.timer_Count_0_LC_5_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14142\,
            lcout => \uart.timer_CountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23877\,
            ce => 'H',
            sr => \N__14184\
        );

    \uart.un4_timer_Count_1_cry_1_c_LC_5_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13974\,
            in2 => \N__14148\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_15_0_\,
            carryout => \uart.un4_timer_Count_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart.timer_Count_2_LC_5_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13949\,
            in2 => \_gnd_net_\,
            in3 => \N__13929\,
            lcout => \uart.timer_CountZ0Z_2\,
            ltout => OPEN,
            carryin => \uart.un4_timer_Count_1_cry_1\,
            carryout => \uart.un4_timer_Count_1_cry_2\,
            clk => \N__23870\,
            ce => 'H',
            sr => \N__14176\
        );

    \uart.timer_Count_3_LC_5_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13924\,
            in2 => \_gnd_net_\,
            in3 => \N__13902\,
            lcout => \uart.timer_CountZ0Z_3\,
            ltout => OPEN,
            carryin => \uart.un4_timer_Count_1_cry_2\,
            carryout => \uart.un4_timer_Count_1_cry_3\,
            clk => \N__23870\,
            ce => 'H',
            sr => \N__14176\
        );

    \uart.timer_Count_4_LC_5_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14118\,
            in2 => \_gnd_net_\,
            in3 => \N__14331\,
            lcout => \uart.timer_CountZ0Z_4\,
            ltout => OPEN,
            carryin => \uart.un4_timer_Count_1_cry_3\,
            carryout => \uart.un4_timer_Count_1_cry_4\,
            clk => \N__23870\,
            ce => 'H',
            sr => \N__14176\
        );

    \uart.timer_Count_5_LC_5_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14327\,
            in2 => \_gnd_net_\,
            in3 => \N__14301\,
            lcout => \uart.timer_CountZ0Z_5\,
            ltout => OPEN,
            carryin => \uart.un4_timer_Count_1_cry_4\,
            carryout => \uart.un4_timer_Count_1_cry_5\,
            clk => \N__23870\,
            ce => 'H',
            sr => \N__14176\
        );

    \uart.timer_Count_6_LC_5_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14289\,
            in2 => \_gnd_net_\,
            in3 => \N__14256\,
            lcout => \uart.timer_CountZ0Z_6\,
            ltout => OPEN,
            carryin => \uart.un4_timer_Count_1_cry_5\,
            carryout => \uart.un4_timer_Count_1_cry_6\,
            clk => \N__23870\,
            ce => 'H',
            sr => \N__14176\
        );

    \uart.timer_Count_7_LC_5_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14233\,
            in2 => \_gnd_net_\,
            in3 => \N__14253\,
            lcout => \uart.timer_CountZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23870\,
            ce => 'H',
            sr => \N__14176\
        );

    \uart.timer_Count_RNIQ9BL_0_LC_5_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14144\,
            in2 => \_gnd_net_\,
            in3 => \N__14117\,
            lcout => \uart.un1_state_2_0_a3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_1_cry_1_c_LC_5_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14079\,
            in2 => \N__14057\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_17_0_\,
            carryout => \reset_module_System.count_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_RNO_0_2_LC_5_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14034\,
            in2 => \_gnd_net_\,
            in3 => \N__14016\,
            lcout => \reset_module_System.count_1_2\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_1\,
            carryout => \reset_module_System.count_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_3_LC_5_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14013\,
            in2 => \_gnd_net_\,
            in3 => \N__14001\,
            lcout => \reset_module_System.countZ0Z_3\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_2\,
            carryout => \reset_module_System.count_1_cry_3\,
            clk => \N__23861\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_4_LC_5_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14468\,
            in2 => \_gnd_net_\,
            in3 => \N__14457\,
            lcout => \reset_module_System.countZ0Z_4\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_3\,
            carryout => \reset_module_System.count_1_cry_4\,
            clk => \N__23861\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_5_LC_5_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14454\,
            in2 => \_gnd_net_\,
            in3 => \N__14442\,
            lcout => \reset_module_System.countZ0Z_5\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_4\,
            carryout => \reset_module_System.count_1_cry_5\,
            clk => \N__23861\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_6_LC_5_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14439\,
            in2 => \_gnd_net_\,
            in3 => \N__14427\,
            lcout => \reset_module_System.countZ0Z_6\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_5\,
            carryout => \reset_module_System.count_1_cry_6\,
            clk => \N__23861\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_7_LC_5_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14424\,
            in2 => \_gnd_net_\,
            in3 => \N__14412\,
            lcout => \reset_module_System.countZ0Z_7\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_6\,
            carryout => \reset_module_System.count_1_cry_7\,
            clk => \N__23861\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_8_LC_5_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14409\,
            in2 => \_gnd_net_\,
            in3 => \N__14397\,
            lcout => \reset_module_System.countZ0Z_8\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_7\,
            carryout => \reset_module_System.count_1_cry_8\,
            clk => \N__23861\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_9_LC_5_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14393\,
            in2 => \_gnd_net_\,
            in3 => \N__14379\,
            lcout => \reset_module_System.countZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_5_18_0_\,
            carryout => \reset_module_System.count_1_cry_9\,
            clk => \N__23856\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_10_LC_5_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14376\,
            in2 => \_gnd_net_\,
            in3 => \N__14364\,
            lcout => \reset_module_System.countZ0Z_10\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_9\,
            carryout => \reset_module_System.count_1_cry_10\,
            clk => \N__23856\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_11_LC_5_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14361\,
            in2 => \_gnd_net_\,
            in3 => \N__14349\,
            lcout => \reset_module_System.countZ0Z_11\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_10\,
            carryout => \reset_module_System.count_1_cry_11\,
            clk => \N__23856\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_12_LC_5_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14345\,
            in2 => \_gnd_net_\,
            in3 => \N__14334\,
            lcout => \reset_module_System.countZ0Z_12\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_11\,
            carryout => \reset_module_System.count_1_cry_12\,
            clk => \N__23856\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_13_LC_5_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14663\,
            in2 => \_gnd_net_\,
            in3 => \N__14568\,
            lcout => \reset_module_System.countZ0Z_13\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_12\,
            carryout => \reset_module_System.count_1_cry_13\,
            clk => \N__23856\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_14_LC_5_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14565\,
            in2 => \_gnd_net_\,
            in3 => \N__14553\,
            lcout => \reset_module_System.countZ0Z_14\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_13\,
            carryout => \reset_module_System.count_1_cry_14\,
            clk => \N__23856\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_15_LC_5_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14687\,
            in2 => \_gnd_net_\,
            in3 => \N__14550\,
            lcout => \reset_module_System.countZ0Z_15\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_14\,
            carryout => \reset_module_System.count_1_cry_15\,
            clk => \N__23856\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_16_LC_5_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14546\,
            in2 => \_gnd_net_\,
            in3 => \N__14535\,
            lcout => \reset_module_System.countZ0Z_16\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_15\,
            carryout => \reset_module_System.count_1_cry_16\,
            clk => \N__23856\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_17_LC_5_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14531\,
            in2 => \_gnd_net_\,
            in3 => \N__14517\,
            lcout => \reset_module_System.countZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_5_19_0_\,
            carryout => \reset_module_System.count_1_cry_17\,
            clk => \N__23852\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_18_LC_5_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14510\,
            in2 => \_gnd_net_\,
            in3 => \N__14496\,
            lcout => \reset_module_System.countZ0Z_18\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_17\,
            carryout => \reset_module_System.count_1_cry_18\,
            clk => \N__23852\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_19_LC_5_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14697\,
            in2 => \_gnd_net_\,
            in3 => \N__14493\,
            lcout => \reset_module_System.countZ0Z_19\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_18\,
            carryout => \reset_module_System.count_1_cry_19\,
            clk => \N__23852\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_20_LC_5_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14486\,
            in2 => \_gnd_net_\,
            in3 => \N__14472\,
            lcout => \reset_module_System.countZ0Z_20\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_19\,
            carryout => \reset_module_System.count_1_cry_20\,
            clk => \N__23852\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_21_LC_5_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14675\,
            in2 => \_gnd_net_\,
            in3 => \N__14700\,
            lcout => \reset_module_System.countZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23852\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_RNI34OR1_21_LC_5_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__14696\,
            in1 => \N__14688\,
            in2 => \N__14676\,
            in3 => \N__14664\,
            lcout => \reset_module_System.reset6_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_esr_RNIJL8F_4_LC_5_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__14792\,
            in1 => \N__14780\,
            in2 => \_gnd_net_\,
            in3 => \N__18826\,
            lcout => \ppm_encoder_1.N_462\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_esr_4_LC_5_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15153\,
            lcout => \ppm_encoder_1.aileronZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23847\,
            ce => \N__16244\,
            sr => \N__23346\
        );

    \ppm_encoder_1.elevator_esr_4_LC_5_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14628\,
            lcout => \ppm_encoder_1.elevatorZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23847\,
            ce => \N__16244\,
            sr => \N__23346\
        );

    \scaler_2.un2_source_data_0_cry_1_c_RNO_LC_5_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__15184\,
            in1 => \N__14607\,
            in2 => \_gnd_net_\,
            in3 => \N__15230\,
            lcout => \scaler_2.un2_source_data_0_cry_1_c_RNO_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_LC_5_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111010101111"
        )
    port map (
            in0 => \N__23504\,
            in1 => \N__18854\,
            in2 => \N__16374\,
            in3 => \N__21210\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23841\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_1_LC_5_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000111110"
        )
    port map (
            in0 => \N__17310\,
            in1 => \N__22132\,
            in2 => \N__24090\,
            in3 => \N__21967\,
            lcout => \ppm_encoder_1.pulses2count_9_0_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNINGL11_6_LC_5_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010101010"
        )
    port map (
            in0 => \N__15367\,
            in1 => \N__19230\,
            in2 => \_gnd_net_\,
            in3 => \N__19538\,
            lcout => \ppm_encoder_1.un2_throttle_iv_0_rn_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_4_LC_5_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000001110000"
        )
    port map (
            in0 => \N__20150\,
            in1 => \N__14793\,
            in2 => \N__22134\,
            in3 => \N__14781\,
            lcout => \ppm_encoder_1.N_369\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_LC_5_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010001010000"
        )
    port map (
            in0 => \N__23505\,
            in1 => \N__19539\,
            in2 => \N__18294\,
            in3 => \N__21209\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23841\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_6_LC_5_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0111011101000100"
        )
    port map (
            in0 => \N__14769\,
            in1 => \N__17487\,
            in2 => \_gnd_net_\,
            in3 => \N__14748\,
            lcout => \ppm_encoder_1.aileronZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23835\,
            ce => 'H',
            sr => \N__23355\
        );

    \ppm_encoder_1.elevator_RNIDJ141_6_LC_5_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000000000"
        )
    port map (
            in0 => \N__14747\,
            in1 => \N__17193\,
            in2 => \N__14739\,
            in3 => \N__17883\,
            lcout => \ppm_encoder_1.pulses2count_9_0_o2_0_6\,
            ltout => \ppm_encoder_1.pulses2count_9_0_o2_0_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNI0LED3_6_LC_5_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14706\,
            in2 => \N__14721\,
            in3 => \N__14718\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un2_throttle_0_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNID1DC5_6_LC_5_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001101001"
        )
    port map (
            in0 => \N__17718\,
            in1 => \N__19187\,
            in2 => \N__14712\,
            in3 => \N__17051\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un1_init_pulses_0_axb_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNI6UPC6_6_LC_5_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__14709\,
            in3 => \N__17933\,
            lcout => \ppm_encoder_1.init_pulses_RNI6UPC6Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.rudder_RNISGN71_6_LC_5_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001110101111"
        )
    port map (
            in0 => \N__18763\,
            in1 => \N__19231\,
            in2 => \N__18881\,
            in3 => \N__19540\,
            lcout => \ppm_encoder_1.un2_throttle_iv_0_sn_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNI31EQ5_9_LC_5_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17216\,
            in2 => \_gnd_net_\,
            in3 => \N__14826\,
            lcout => \ppm_encoder_1.init_pulses_RNI31EQ5Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNICBGI_10_LC_5_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__19954\,
            in1 => \N__18876\,
            in2 => \_gnd_net_\,
            in3 => \N__18782\,
            lcout => \ppm_encoder_1.N_415\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNI55NT_10_LC_5_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010100000"
        )
    port map (
            in0 => \N__18783\,
            in1 => \N__15674\,
            in2 => \N__15650\,
            in3 => \N__18877\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.N_414_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.rudder_RNI5GRA2_10_LC_5_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__19927\,
            in1 => \N__14880\,
            in2 => \N__14874\,
            in3 => \N__19625\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un2_throttle_iv_0_1_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNITDM64_10_LC_5_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001101001"
        )
    port map (
            in0 => \N__22526\,
            in1 => \N__17713\,
            in2 => \N__14871\,
            in3 => \N__17060\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un1_init_pulses_0_axb_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIJ2JB5_10_LC_5_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__14868\,
            in3 => \N__17834\,
            lcout => \ppm_encoder_1.init_pulses_RNIJ2JB5Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNI4MTK_9_LC_5_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__19000\,
            in1 => \N__18776\,
            in2 => \_gnd_net_\,
            in3 => \N__18897\,
            lcout => \ppm_encoder_1.N_412\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNILQ941_9_LC_5_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000010000000"
        )
    port map (
            in0 => \N__18898\,
            in1 => \N__14854\,
            in2 => \N__18788\,
            in3 => \N__15310\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.N_411_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.rudder_RNI5BFJ2_9_LC_5_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__18955\,
            in1 => \N__14838\,
            in2 => \N__14832\,
            in3 => \N__19624\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un2_throttle_iv_0_1_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNILQDI4_9_LC_5_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001101001"
        )
    port map (
            in0 => \N__24161\,
            in1 => \N__17717\,
            in2 => \N__14829\,
            in3 => \N__17059\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_axb_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_9_LC_5_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__14820\,
            in1 => \N__14814\,
            in2 => \N__17540\,
            in3 => \N__15311\,
            lcout => \ppm_encoder_1.aileronZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23825\,
            ce => 'H',
            sr => \N__23364\
        );

    \ppm_encoder_1.rudder_9_LC_5_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011110000"
        )
    port map (
            in0 => \N__15297\,
            in1 => \N__15288\,
            in2 => \N__18965\,
            in3 => \N__17508\,
            lcout => \ppm_encoder_1.rudderZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23820\,
            ce => 'H',
            sr => \N__23370\
        );

    \ppm_encoder_1.elevator_10_LC_5_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__15267\,
            in1 => \N__15243\,
            in2 => \N__17541\,
            in3 => \N__15673\,
            lcout => \ppm_encoder_1.elevatorZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23820\,
            ce => 'H',
            sr => \N__23370\
        );

    \scaler_2.source_data_1_4_LC_5_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001011011000"
        )
    port map (
            in0 => \N__14948\,
            in1 => \N__15237\,
            in2 => \N__15152\,
            in3 => \N__15195\,
            lcout => scaler_2_data_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23820\,
            ce => 'H',
            sr => \N__23370\
        );

    \ppm_encoder_1.rudder_12_LC_5_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0110011011110000"
        )
    port map (
            in0 => \N__15135\,
            in1 => \N__15117\,
            in2 => \N__18493\,
            in3 => \N__17507\,
            lcout => \ppm_encoder_1.rudderZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23820\,
            ce => 'H',
            sr => \N__23370\
        );

    \uart_frame_decoder.source_CH1data_esr_4_LC_5_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15105\,
            lcout => \frame_decoder_CH1data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23815\,
            ce => \N__15024\,
            sr => \N__23377\
        );

    \ppm_encoder_1.throttle_12_LC_5_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__15000\,
            in1 => \N__14994\,
            in2 => \N__17560\,
            in3 => \N__19360\,
            lcout => \ppm_encoder_1.throttleZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23809\,
            ce => 'H',
            sr => \N__23383\
        );

    \ppm_encoder_1.throttle_13_LC_5_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1001100111110000"
        )
    port map (
            in0 => \N__14979\,
            in1 => \N__14961\,
            in2 => \N__15867\,
            in3 => \N__17539\,
            lcout => \ppm_encoder_1.throttleZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23809\,
            ce => 'H',
            sr => \N__23383\
        );

    \scaler_1.source_data_1_esr_ctle_14_LC_5_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14939\,
            in2 => \_gnd_net_\,
            in3 => \N__23492\,
            lcout => frame_decoder_dv_c_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_sync.aux_0__0__0_LC_7_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15414\,
            lcout => \uart_sync.aux_0__0_Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23883\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.rudder_esr_ctle_14_LC_7_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17462\,
            in2 => \_gnd_net_\,
            in3 => \N__23491\,
            lcout => \ppm_encoder_1.scaler_1_dv_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_6_LC_7_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011110000"
        )
    port map (
            in0 => \N__18780\,
            in1 => \N__15375\,
            in2 => \N__15351\,
            in3 => \N__18893\,
            lcout => \ppm_encoder_1.N_301\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNI7JM64_11_LC_7_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001110010110"
        )
    port map (
            in0 => \N__15333\,
            in1 => \N__17712\,
            in2 => \N__20043\,
            in3 => \N__17050\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un1_init_pulses_0_axb_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIV8JB5_11_LC_7_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__15336\,
            in3 => \N__19262\,
            lcout => \ppm_encoder_1.init_pulses_RNIV8JB5Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.rudder_RNIEKRA2_11_LC_7_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001110"
        )
    port map (
            in0 => \N__20397\,
            in1 => \N__15729\,
            in2 => \N__18413\,
            in3 => \N__15564\,
            lcout => \ppm_encoder_1.un2_throttle_iv_0_2_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNI0O131_0_17_LC_7_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001111000"
        )
    port map (
            in0 => \N__24056\,
            in1 => \N__21785\,
            in2 => \N__20931\,
            in3 => \N__21223\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_axb_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_esr_RNII84K_4_LC_7_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__17192\,
            in1 => \N__19877\,
            in2 => \_gnd_net_\,
            in3 => \N__20675\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un2_throttle_iv_i_i_1_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_1_rep2_RNIGT971_LC_7_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20242\,
            in2 => \N__15327\,
            in3 => \N__15324\,
            lcout => \ppm_encoder_1.un2_throttle_iv_i_i_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNI81081_0_4_LC_7_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001101100"
        )
    port map (
            in0 => \N__19587\,
            in1 => \N__22632\,
            in2 => \N__17817\,
            in3 => \N__21207\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_0_LC_7_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010011001"
        )
    port map (
            in0 => \N__21208\,
            in1 => \N__20458\,
            in2 => \_gnd_net_\,
            in3 => \N__17737\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un1_init_pulses_11_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_0_LC_7_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000000011010001"
        )
    port map (
            in0 => \N__20459\,
            in1 => \N__16918\,
            in2 => \N__15429\,
            in3 => \N__16793\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23830\,
            ce => 'H',
            sr => \N__23350\
        );

    \ppm_encoder_1.init_pulses_4_LC_7_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__16792\,
            in1 => \N__17973\,
            in2 => \N__16923\,
            in3 => \N__15471\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23830\,
            ce => 'H',
            sr => \N__23350\
        );

    \ppm_encoder_1.init_pulses_RNIR7863_4_LC_7_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001101001"
        )
    port map (
            in0 => \N__17710\,
            in1 => \N__15426\,
            in2 => \N__22640\,
            in3 => \N__17044\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un1_init_pulses_0_axb_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNI398E4_4_LC_7_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__15420\,
            in3 => \N__16449\,
            lcout => \ppm_encoder_1.init_pulses_RNI398E4Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNI83R42_0_LC_7_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__17735\,
            in1 => \N__20460\,
            in2 => \_gnd_net_\,
            in3 => \N__21205\,
            lcout => \ppm_encoder_1.init_pulses_RNI83R42Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIR0RR1_13_LC_7_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001110010110"
        )
    port map (
            in0 => \N__21206\,
            in1 => \N__17709\,
            in2 => \N__21351\,
            in3 => \N__17736\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIMR0V_0_0_LC_7_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20449\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_23_0_\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_1_LC_7_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17076\,
            in2 => \N__17283\,
            in3 => \N__15417\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_1\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_0\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_2_LC_7_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16323\,
            in2 => \N__18054\,
            in3 => \N__15483\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_2\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_1\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_3_LC_7_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16956\,
            in2 => \N__17265\,
            in3 => \N__15480\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_3\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_2\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_4_LC_7_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15477\,
            in2 => \N__16448\,
            in3 => \N__15465\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_4\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_3\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_5_LC_7_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16308\,
            in2 => \N__16188\,
            in3 => \N__15462\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_5\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_4\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_6_LC_7_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15459\,
            in2 => \N__17934\,
            in3 => \N__15450\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_6\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_5\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_7_LC_7_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16380\,
            in2 => \N__17247\,
            in3 => \N__15447\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_7\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_6\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_8_LC_7_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16164\,
            in2 => \N__18618\,
            in3 => \N__15444\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_8\,
            ltout => OPEN,
            carryin => \bfn_7_24_0_\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_9_LC_7_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15441\,
            in2 => \N__17220\,
            in3 => \N__15432\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_9\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_8\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_10_LC_7_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15537\,
            in2 => \N__17838\,
            in3 => \N__15528\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_10\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_9\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_11_LC_7_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15525\,
            in2 => \N__19266\,
            in3 => \N__15516\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_11\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_10\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_12_LC_7_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16389\,
            in2 => \N__19296\,
            in3 => \N__15513\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_12\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_11\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_13_LC_7_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18156\,
            in2 => \N__15792\,
            in3 => \N__15510\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_13\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_12\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_2_14_LC_7_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17583\,
            in2 => \N__15585\,
            in3 => \N__15507\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_14\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_13\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_15_LC_7_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16476\,
            in2 => \N__15576\,
            in3 => \N__15504\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_15\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_14\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_16_LC_7_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17757\,
            in2 => \_gnd_net_\,
            in3 => \N__15501\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_16\,
            ltout => OPEN,
            carryin => \bfn_7_25_0_\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_17_LC_7_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15498\,
            in2 => \_gnd_net_\,
            in3 => \N__15489\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_17\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_16\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_18_LC_7_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__20875\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15486\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNISRB55_14_LC_7_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010110010110"
        )
    port map (
            in0 => \N__17715\,
            in1 => \N__21461\,
            in2 => \N__21512\,
            in3 => \N__16317\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un1_init_pulses_0_axb_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNINK8A6_14_LC_7_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__15588\,
            in3 => \N__17579\,
            lcout => \ppm_encoder_1.init_pulses_RNINK8A6Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNIN4HJ_12_LC_7_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000001010"
        )
    port map (
            in0 => \N__20104\,
            in1 => \N__19043\,
            in2 => \N__19373\,
            in3 => \N__20218\,
            lcout => \ppm_encoder_1.un2_throttle_iv_0_1_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIJJM71_15_LC_7_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__21813\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16472\,
            lcout => \ppm_encoder_1.init_pulses_RNIJJM71Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_RNI3HMS_11_LC_7_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__20103\,
            in1 => \N__20217\,
            in2 => \_gnd_net_\,
            in3 => \N__19406\,
            lcout => \ppm_encoder_1.N_403\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_0_LC_7_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111111001101"
        )
    port map (
            in0 => \N__21230\,
            in1 => \N__23513\,
            in2 => \N__16363\,
            in3 => \N__21929\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23810\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_esr_RNIUAMB2_14_LC_7_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000100"
        )
    port map (
            in0 => \N__22121\,
            in1 => \N__21880\,
            in2 => \N__15552\,
            in3 => \N__16404\,
            lcout => \ppm_encoder_1.N_304\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIFN3K_2_LC_7_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__20235\,
            in1 => \N__20119\,
            in2 => \_gnd_net_\,
            in3 => \N__19830\,
            lcout => \ppm_encoder_1.N_443\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_1_rep2_LC_7_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110000000110"
        )
    port map (
            in0 => \N__21928\,
            in1 => \N__20236\,
            in2 => \N__23532\,
            in3 => \N__21231\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23810\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m2_i_0_LC_7_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010101010"
        )
    port map (
            in0 => \N__21882\,
            in1 => \N__19745\,
            in2 => \_gnd_net_\,
            in3 => \N__20349\,
            lcout => \ppm_encoder_1.N_114\,
            ltout => \ppm_encoder_1.N_114_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_0_rep2_LC_7_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011001111"
        )
    port map (
            in0 => \N__20120\,
            in1 => \N__23523\,
            in2 => \N__15678\,
            in3 => \N__21233\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23810\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_10_LC_7_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010011100000000"
        )
    port map (
            in0 => \N__21881\,
            in1 => \N__15675\,
            in2 => \N__15651\,
            in3 => \N__22122\,
            lcout => \ppm_encoder_1.N_383\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_2_rep2_LC_7_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000001100"
        )
    port map (
            in0 => \N__20350\,
            in1 => \N__18289\,
            in2 => \N__23533\,
            in3 => \N__21232\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23810\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_57_c_RNIFNBA1_LC_7_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__19769\,
            in1 => \N__24558\,
            in2 => \N__20815\,
            in3 => \N__24411\,
            lcout => \ppm_encoder_1.N_348\,
            ltout => \ppm_encoder_1.N_348_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_14_LC_7_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110010"
        )
    port map (
            in0 => \N__16843\,
            in1 => \N__18321\,
            in2 => \N__15621\,
            in3 => \N__18102\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.init_pulses_18_i_0_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_14_LC_7_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000110100001100"
        )
    port map (
            in0 => \N__15606\,
            in1 => \N__15618\,
            in2 => \N__15609\,
            in3 => \N__17716\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23803\,
            ce => 'H',
            sr => \N__23378\
        );

    \ppm_encoder_1.init_pulses_RNO_1_14_LC_7_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000101000100"
        )
    port map (
            in0 => \N__21229\,
            in1 => \N__20348\,
            in2 => \N__21773\,
            in3 => \N__21602\,
            lcout => \ppm_encoder_1.init_pulses_18_i_a2_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_3_rep2_RNIMOAF1_LC_7_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101100101"
        )
    port map (
            in0 => \N__20347\,
            in1 => \N__19770\,
            in2 => \N__21620\,
            in3 => \N__21228\,
            lcout => \ppm_encoder_1.N_241\,
            ltout => \ppm_encoder_1.N_241_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_16_LC_7_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__16791\,
            in1 => \N__15600\,
            in2 => \N__15591\,
            in3 => \N__18369\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23803\,
            ce => 'H',
            sr => \N__23378\
        );

    \ppm_encoder_1.elevator_RNIDBNT_13_LC_7_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010001000"
        )
    port map (
            in0 => \N__15806\,
            in1 => \N__20241\,
            in2 => \N__15741\,
            in3 => \N__20128\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.pulses2count_9_0_o2_0_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNI06LN1_13_LC_7_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111000"
        )
    port map (
            in0 => \N__15866\,
            in1 => \N__21907\,
            in2 => \N__15849\,
            in3 => \N__22110\,
            lcout => \ppm_encoder_1.N_303\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_13_LC_7_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__15807\,
            in1 => \N__15846\,
            in2 => \N__17564\,
            in3 => \N__15822\,
            lcout => \ppm_encoder_1.aileronZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23796\,
            ce => 'H',
            sr => \N__23384\
        );

    \ppm_encoder_1.rudder_RNIAAE02_13_LC_7_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__20659\,
            in1 => \N__20362\,
            in2 => \_gnd_net_\,
            in3 => \N__17061\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un2_throttle_iv_0_0_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIJ94E4_13_LC_7_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101011010101001"
        )
    port map (
            in0 => \N__21349\,
            in1 => \N__21287\,
            in2 => \N__15798\,
            in3 => \N__17714\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un1_init_pulses_0_axb_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIC11J5_13_LC_7_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__15795\,
            in3 => \N__18145\,
            lcout => \ppm_encoder_1.init_pulses_RNIC11J5Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_13_LC_7_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__15740\,
            in1 => \N__15780\,
            in2 => \N__17565\,
            in3 => \N__15753\,
            lcout => \ppm_encoder_1.elevatorZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23796\,
            ce => 'H',
            sr => \N__23384\
        );

    \ppm_encoder_1.elevator_RNIL2HJ_11_LC_7_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000001100"
        )
    port map (
            in0 => \N__18457\,
            in1 => \N__20127\,
            in2 => \N__19988\,
            in3 => \N__20240\,
            lcout => \ppm_encoder_1.un2_throttle_iv_0_1_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_11_LC_7_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101101011001100"
        )
    port map (
            in0 => \N__15720\,
            in1 => \N__18458\,
            in2 => \N__15693\,
            in3 => \N__17534\,
            lcout => \ppm_encoder_1.elevatorZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23791\,
            ce => 'H',
            sr => \N__23392\
        );

    \ppm_encoder_1.throttle_11_LC_7_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101011001010"
        )
    port map (
            in0 => \N__19984\,
            in1 => \N__16023\,
            in2 => \N__17559\,
            in3 => \N__16005\,
            lcout => \ppm_encoder_1.throttleZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23791\,
            ce => 'H',
            sr => \N__23392\
        );

    \ppm_encoder_1.aileron_12_LC_8_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__15996\,
            in1 => \N__15972\,
            in2 => \N__17552\,
            in3 => \N__19081\,
            lcout => \ppm_encoder_1.aileronZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23842\,
            ce => 'H',
            sr => \N__23344\
        );

    \ppm_encoder_1.throttle_2_LC_8_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17520\,
            in2 => \_gnd_net_\,
            in3 => \N__20614\,
            lcout => \ppm_encoder_1.throttleZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23842\,
            ce => 'H',
            sr => \N__23344\
        );

    \ppm_encoder_1.throttle_RNI3LTK_8_LC_8_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__18427\,
            in1 => \N__18759\,
            in2 => \_gnd_net_\,
            in3 => \N__18885\,
            lcout => \ppm_encoder_1.N_418\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNIJO941_8_LC_8_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000010000000"
        )
    port map (
            in0 => \N__18886\,
            in1 => \N__18589\,
            in2 => \N__18781\,
            in3 => \N__18571\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.N_417_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.rudder_RNI17FJ2_8_LC_8_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__18550\,
            in1 => \N__15957\,
            in2 => \N__15951\,
            in3 => \N__19597\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un2_throttle_iv_0_1_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIGLDI4_8_LC_8_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001101001"
        )
    port map (
            in0 => \N__22692\,
            in1 => \N__17705\,
            in2 => \N__15948\,
            in3 => \N__17049\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_8_LC_8_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__15945\,
            in1 => \N__15933\,
            in2 => \N__17561\,
            in3 => \N__18572\,
            lcout => \ppm_encoder_1.aileronZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23836\,
            ce => 'H',
            sr => \N__23347\
        );

    \ppm_encoder_1.throttle_8_LC_8_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011110010101010"
        )
    port map (
            in0 => \N__18428\,
            in1 => \N__15912\,
            in2 => \N__15894\,
            in3 => \N__17548\,
            lcout => \ppm_encoder_1.throttleZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23836\,
            ce => 'H',
            sr => \N__23347\
        );

    \ppm_encoder_1.elevator_8_LC_8_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__16155\,
            in1 => \N__16140\,
            in2 => \N__17562\,
            in3 => \N__18590\,
            lcout => \ppm_encoder_1.elevatorZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23836\,
            ce => 'H',
            sr => \N__23347\
        );

    \ppm_encoder_1.elevator_esr_5_LC_8_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16113\,
            lcout => \ppm_encoder_1.elevatorZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23831\,
            ce => \N__16243\,
            sr => \N__23351\
        );

    \ppm_encoder_1.rudder_esr_4_LC_8_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16098\,
            lcout => \ppm_encoder_1.rudderZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23831\,
            ce => \N__16243\,
            sr => \N__23351\
        );

    \ppm_encoder_1.throttle_esr_4_LC_8_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16074\,
            lcout => \ppm_encoder_1.throttleZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23831\,
            ce => \N__16243\,
            sr => \N__23351\
        );

    \ppm_encoder_1.throttle_esr_5_LC_8_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__16050\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \ppm_encoder_1.throttleZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23831\,
            ce => \N__16243\,
            sr => \N__23351\
        );

    \ppm_encoder_1.aileron_esr_RNITLTI_5_LC_8_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000100010"
        )
    port map (
            in0 => \N__17879\,
            in1 => \N__16287\,
            in2 => \N__16038\,
            in3 => \N__17188\,
            lcout => \ppm_encoder_1.pulses2count_9_i_o2_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.rudder_esr_RNI4IR61_5_LC_8_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001011110011"
        )
    port map (
            in0 => \N__18741\,
            in1 => \N__19554\,
            in2 => \N__22310\,
            in3 => \N__18902\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un1_init_pulses_0_axb_5_1_sn_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_esr_RNI8RGL2_5_LC_8_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110011111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16302\,
            in2 => \N__16029\,
            in3 => \N__18920\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un1_init_pulses_0_axb_5_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIK6FK4_5_LC_8_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101101001"
        )
    port map (
            in0 => \N__22569\,
            in1 => \N__17711\,
            in2 => \N__16026\,
            in3 => \N__17045\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un1_init_pulses_0_axb_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIT8FS5_5_LC_8_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16184\,
            in2 => \N__16311\,
            in3 => \_gnd_net_\,
            lcout => \ppm_encoder_1.init_pulses_RNIT8FS5Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_esr_RNI7JNR_5_LC_8_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010101010"
        )
    port map (
            in0 => \N__18932\,
            in1 => \N__22303\,
            in2 => \_gnd_net_\,
            in3 => \N__19553\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_axb_5_1_rn_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_esr_5_LC_8_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16296\,
            lcout => \ppm_encoder_1.aileronZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23826\,
            ce => \N__16254\,
            sr => \N__23356\
        );

    \ppm_encoder_1.rudder_esr_5_LC_8_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16281\,
            lcout => \ppm_encoder_1.rudderZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23826\,
            ce => \N__16254\,
            sr => \N__23356\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_LC_8_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110000000110"
        )
    port map (
            in0 => \N__21974\,
            in1 => \N__18775\,
            in2 => \N__23534\,
            in3 => \N__21055\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23821\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNI92081_5_LC_8_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011010011110000"
        )
    port map (
            in0 => \N__21054\,
            in1 => \N__17807\,
            in2 => \N__22576\,
            in3 => \N__19603\,
            lcout => \ppm_encoder_1.N_252_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNITQDQ5_8_LC_8_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18611\,
            in2 => \_gnd_net_\,
            in3 => \N__16173\,
            lcout => \ppm_encoder_1.init_pulses_RNITQDQ5Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIHO7D_1_LC_8_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__17864\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17181\,
            lcout => \ppm_encoder_1.N_235\,
            ltout => \ppm_encoder_1.N_235_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNII7Q51_3_LC_8_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101011"
        )
    port map (
            in0 => \N__19860\,
            in1 => \N__19815\,
            in2 => \N__16158\,
            in3 => \N__21053\,
            lcout => \ppm_encoder_1.N_246\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIUBDK6_7_LC_8_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17234\,
            in2 => \_gnd_net_\,
            in3 => \N__17199\,
            lcout => \ppm_encoder_1.init_pulses_RNIUBDK6Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_0_LC_8_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101011110011"
        )
    port map (
            in0 => \N__17183\,
            in1 => \N__16370\,
            in2 => \N__23535\,
            in3 => \N__21056\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23821\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI6LFQ_1_LC_8_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001111010011"
        )
    port map (
            in0 => \N__17865\,
            in1 => \N__19859\,
            in2 => \N__19826\,
            in3 => \N__17182\,
            lcout => \ppm_encoder_1.N_305\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_RNI4IMS_12_LC_8_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001010"
        )
    port map (
            in0 => \N__20243\,
            in1 => \_gnd_net_\,
            in2 => \N__19088\,
            in3 => \N__20133\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.N_407_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.rudder_RNIIORA2_12_LC_8_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111110"
        )
    port map (
            in0 => \N__16338\,
            in1 => \N__20398\,
            in2 => \N__16332\,
            in3 => \N__18494\,
            lcout => \ppm_encoder_1.un2_throttle_iv_0_2_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNIUETK_2_LC_8_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__20615\,
            in1 => \N__20132\,
            in2 => \_gnd_net_\,
            in3 => \N__18740\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un1_init_pulses_0_axb_2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNI7NRJ2_2_LC_8_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101101001"
        )
    port map (
            in0 => \N__20540\,
            in1 => \N__17687\,
            in2 => \N__16329\,
            in3 => \N__17036\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un1_init_pulses_0_axb_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIE48O3_2_LC_8_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16326\,
            in3 => \N__18040\,
            lcout => \ppm_encoder_1.init_pulses_RNIE48O3Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.rudder_esr_RNIKMK32_14_LC_8_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__21540\,
            in1 => \N__20399\,
            in2 => \_gnd_net_\,
            in3 => \N__17037\,
            lcout => \ppm_encoder_1.un2_throttle_iv_0_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNI81081_4_LC_8_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001101100"
        )
    port map (
            in0 => \N__17805\,
            in1 => \N__22639\,
            in2 => \N__19620\,
            in3 => \N__21083\,
            lcout => \ppm_encoder_1.N_251_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_3_rep1_LC_8_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010100000001"
        )
    port map (
            in0 => \N__23512\,
            in1 => \N__21167\,
            in2 => \N__18654\,
            in3 => \N__17806\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_3_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23816\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIPNS41_13_LC_8_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101001011110000"
        )
    port map (
            in0 => \N__19713\,
            in1 => \N__21062\,
            in2 => \N__21336\,
            in3 => \N__19626\,
            lcout => \ppm_encoder_1.N_259_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_esr_RNI14O81_14_LC_8_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000100010"
        )
    port map (
            in0 => \N__20222\,
            in1 => \N__16428\,
            in2 => \N__16419\,
            in3 => \N__20115\,
            lcout => \ppm_encoder_1.pulses2count_9_i_o2_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNICOM64_12_LC_8_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001110010110"
        )
    port map (
            in0 => \N__16398\,
            in1 => \N__17669\,
            in2 => \N__19337\,
            in3 => \N__17058\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un1_init_pulses_0_axb_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNI5FJB5_12_LC_8_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16392\,
            in3 => \N__19295\,
            lcout => \ppm_encoder_1.init_pulses_RNI5FJB5Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIDCUU1_6_LC_8_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010110010110"
        )
    port map (
            in0 => \N__17668\,
            in1 => \N__21064\,
            in2 => \N__19180\,
            in3 => \N__17748\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un1_init_pulses_3_axb_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNI69BV2_6_LC_8_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16383\,
            in3 => \N__17916\,
            lcout => \ppm_encoder_1.init_pulses_RNI69BV2Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIPSC01_6_LC_8_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001101010101010"
        )
    port map (
            in0 => \N__19170\,
            in1 => \N__21061\,
            in2 => \N__17813\,
            in3 => \N__19822\,
            lcout => \ppm_encoder_1.N_253_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNI5UV71_1_LC_8_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111101000000"
        )
    port map (
            in0 => \N__21063\,
            in1 => \N__17802\,
            in2 => \N__19632\,
            in3 => \N__17304\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIKON03_13_LC_8_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18131\,
            in2 => \_gnd_net_\,
            in3 => \N__16530\,
            lcout => \ppm_encoder_1.init_pulses_RNIKON03Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_13_LC_8_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__16786\,
            in1 => \N__18111\,
            in2 => \N__16878\,
            in3 => \N__16518\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23804\,
            ce => 'H',
            sr => \N__23379\
        );

    \ppm_encoder_1.init_pulses_17_LC_8_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0011000100100000"
        )
    port map (
            in0 => \N__16863\,
            in1 => \N__16789\,
            in2 => \N__18354\,
            in3 => \N__16509\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23804\,
            ce => 'H',
            sr => \N__23379\
        );

    \ppm_encoder_1.init_pulses_18_LC_8_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__16788\,
            in1 => \N__18336\,
            in2 => \N__16880\,
            in3 => \N__16503\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23804\,
            ce => 'H',
            sr => \N__23379\
        );

    \ppm_encoder_1.init_pulses_1_LC_8_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0010001100100000"
        )
    port map (
            in0 => \N__18069\,
            in1 => \N__16790\,
            in2 => \N__16881\,
            in3 => \N__16497\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23804\,
            ce => 'H',
            sr => \N__23379\
        );

    \ppm_encoder_1.init_pulses_15_LC_8_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__16787\,
            in1 => \N__18378\,
            in2 => \N__16879\,
            in3 => \N__16485\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23804\,
            ce => 'H',
            sr => \N__23379\
        );

    \ppm_encoder_1.init_pulses_RNISPS41_15_LC_8_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001111000"
        )
    port map (
            in0 => \N__19746\,
            in1 => \N__20342\,
            in2 => \N__21817\,
            in3 => \N__21145\,
            lcout => \ppm_encoder_1.N_245_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIF6081_9_LC_8_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001110011001100"
        )
    port map (
            in0 => \N__21211\,
            in1 => \N__24147\,
            in2 => \N__19765\,
            in3 => \N__20343\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_9_LC_8_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__16782\,
            in1 => \N__18213\,
            in2 => \N__16877\,
            in3 => \N__16461\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23797\,
            ce => 'H',
            sr => \N__23385\
        );

    \ppm_encoder_1.init_pulses_RNINKS41_10_LC_8_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001110011001100"
        )
    port map (
            in0 => \N__21212\,
            in1 => \N__22512\,
            in2 => \N__19766\,
            in3 => \N__20344\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_10_LC_8_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__16780\,
            in1 => \N__16596\,
            in2 => \N__16875\,
            in3 => \N__18198\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23797\,
            ce => 'H',
            sr => \N__23385\
        );

    \ppm_encoder_1.init_pulses_RNIOLS41_0_11_LC_8_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001110011001100"
        )
    port map (
            in0 => \N__21213\,
            in1 => \N__20014\,
            in2 => \N__19767\,
            in3 => \N__20345\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_11_LC_8_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000101100001000"
        )
    port map (
            in0 => \N__18180\,
            in1 => \N__16853\,
            in2 => \N__16800\,
            in3 => \N__16587\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23797\,
            ce => 'H',
            sr => \N__23385\
        );

    \ppm_encoder_1.init_pulses_RNIPMS41_0_12_LC_8_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001110011001100"
        )
    port map (
            in0 => \N__21214\,
            in1 => \N__19318\,
            in2 => \N__19768\,
            in3 => \N__20346\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_12_LC_8_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__16781\,
            in1 => \N__18165\,
            in2 => \N__16876\,
            in3 => \N__16578\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23797\,
            ce => 'H',
            sr => \N__23385\
        );

    \ppm_encoder_1.init_pulses_2_LC_8_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__16794\,
            in1 => \N__18018\,
            in2 => \N__16919\,
            in3 => \N__16569\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23792\,
            ce => 'H',
            sr => \N__23393\
        );

    \ppm_encoder_1.init_pulses_3_LC_8_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011011000"
        )
    port map (
            in0 => \N__16910\,
            in1 => \N__17997\,
            in2 => \N__16557\,
            in3 => \N__16799\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23792\,
            ce => 'H',
            sr => \N__23393\
        );

    \ppm_encoder_1.init_pulses_5_LC_8_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__16795\,
            in1 => \N__17952\,
            in2 => \N__16920\,
            in3 => \N__16542\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23792\,
            ce => 'H',
            sr => \N__23393\
        );

    \ppm_encoder_1.init_pulses_6_LC_8_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001100100000"
        )
    port map (
            in0 => \N__17895\,
            in1 => \N__16797\,
            in2 => \N__16922\,
            in3 => \N__16947\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23792\,
            ce => 'H',
            sr => \N__23393\
        );

    \ppm_encoder_1.init_pulses_7_LC_8_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__16796\,
            in1 => \N__18243\,
            in2 => \N__16921\,
            in3 => \N__16935\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23792\,
            ce => 'H',
            sr => \N__23393\
        );

    \ppm_encoder_1.init_pulses_8_LC_8_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0011000100100000"
        )
    port map (
            in0 => \N__16914\,
            in1 => \N__16798\,
            in2 => \N__18231\,
            in3 => \N__16722\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23792\,
            ce => 'H',
            sr => \N__23393\
        );

    \CONSTANT_ONE_LUT4_LC_9_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.rudder_8_LC_9_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011110000"
        )
    port map (
            in0 => \N__16710\,
            in1 => \N__16698\,
            in2 => \N__18555\,
            in3 => \N__17459\,
            lcout => \ppm_encoder_1.rudderZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23827\,
            ce => 'H',
            sr => \N__23357\
        );

    \ppm_encoder_1.throttle_7_LC_9_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__16674\,
            in1 => \N__16656\,
            in2 => \N__17509\,
            in3 => \N__18534\,
            lcout => \ppm_encoder_1.throttleZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23827\,
            ce => 'H',
            sr => \N__23357\
        );

    \ppm_encoder_1.rudder_7_LC_9_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011110000"
        )
    port map (
            in0 => \N__16638\,
            in1 => \N__16623\,
            in2 => \N__22283\,
            in3 => \N__17458\,
            lcout => \ppm_encoder_1.rudderZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23827\,
            ce => 'H',
            sr => \N__23357\
        );

    \ppm_encoder_1.rudder_RNITHN71_7_LC_9_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010011110101"
        )
    port map (
            in0 => \N__19552\,
            in1 => \N__18739\,
            in2 => \N__22279\,
            in3 => \N__18901\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un2_throttle_iv_0_sn_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNI5QED3_7_LC_9_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__18512\,
            in1 => \_gnd_net_\,
            in2 => \N__16599\,
            in3 => \N__17133\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un2_throttle_0_0_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIJ7DC5_7_LC_9_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100110010110"
        )
    port map (
            in0 => \N__19467\,
            in1 => \N__17703\,
            in2 => \N__17202\,
            in3 => \N__17029\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNIFL141_7_LC_9_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101100000000"
        )
    port map (
            in0 => \N__17184\,
            in1 => \N__17087\,
            in2 => \N__17151\,
            in3 => \N__17872\,
            lcout => \ppm_encoder_1.pulses2count_9_i_o2_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNIPIL11_7_LC_9_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011101010101"
        )
    port map (
            in0 => \N__18532\,
            in1 => \N__22269\,
            in2 => \_gnd_net_\,
            in3 => \N__19551\,
            lcout => \ppm_encoder_1.un2_throttle_iv_0_rn_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_7_LC_9_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__17127\,
            in1 => \N__17112\,
            in2 => \N__17535\,
            in3 => \N__17088\,
            lcout => \ppm_encoder_1.aileronZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23822\,
            ce => 'H',
            sr => \N__23361\
        );

    \ppm_encoder_1.init_pulses_RNI4LRJ2_1_LC_9_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001110010110"
        )
    port map (
            in0 => \N__17067\,
            in1 => \N__17306\,
            in2 => \N__17704\,
            in3 => \N__17027\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un1_init_pulses_0_axb_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIOC8K3_1_LC_9_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17079\,
            in3 => \N__17276\,
            lcout => \ppm_encoder_1.init_pulses_RNIOC8K3Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNISDTK_1_LC_9_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__20770\,
            in1 => \N__18735\,
            in2 => \_gnd_net_\,
            in3 => \N__18899\,
            lcout => \ppm_encoder_1.N_426\,
            ltout => \ppm_encoder_1.N_426_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNI6NRJ2_3_LC_9_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110001110011100"
        )
    port map (
            in0 => \N__17028\,
            in1 => \N__20586\,
            in2 => \N__16962\,
            in3 => \N__17666\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un1_init_pulses_0_axb_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNISG8K3_3_LC_9_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16959\,
            in3 => \N__17258\,
            lcout => \ppm_encoder_1.init_pulses_RNISG8K3Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_1_LC_9_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17563\,
            in2 => \_gnd_net_\,
            in3 => \N__20771\,
            lcout => \ppm_encoder_1.throttleZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23817\,
            ce => 'H',
            sr => \N__23365\
        );

    \ppm_encoder_1.init_pulses_RNIKNC01_1_LC_9_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011100001000"
        )
    port map (
            in0 => \N__17803\,
            in1 => \N__19820\,
            in2 => \N__21130\,
            in3 => \N__17305\,
            lcout => \ppm_encoder_1.N_248_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIMPC01_3_LC_9_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001111000"
        )
    port map (
            in0 => \N__19821\,
            in1 => \N__17804\,
            in2 => \N__20591\,
            in3 => \N__21060\,
            lcout => \ppm_encoder_1.N_250_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIB4081_7_LC_9_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011010011110000"
        )
    port map (
            in0 => \N__21085\,
            in1 => \N__19593\,
            in2 => \N__19475\,
            in3 => \N__17811\,
            lcout => \ppm_encoder_1.N_254_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.PPM_STATE_fast_RNICIAB_0_LC_9_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19425\,
            in3 => \N__22835\,
            lcout => \ppm_encoder_1.PPM_STATE_fast_RNICIABZ0Z_0\,
            ltout => \ppm_encoder_1.PPM_STATE_fast_RNICIABZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIE6081_9_LC_9_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010011010101010"
        )
    port map (
            in0 => \N__24157\,
            in1 => \N__19686\,
            in2 => \N__17223\,
            in3 => \N__19592\,
            lcout => \ppm_encoder_1.N_246_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIK17J_3_LC_9_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110111"
        )
    port map (
            in0 => \N__19858\,
            in1 => \N__19816\,
            in2 => \N__24405\,
            in3 => \N__22836\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIK17JZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_3_LC_9_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000000010001"
        )
    port map (
            in0 => \N__23506\,
            in1 => \N__18640\,
            in2 => \N__19866\,
            in3 => \N__21204\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23811\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_2_LC_9_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001000010000"
        )
    port map (
            in0 => \N__21202\,
            in1 => \N__23507\,
            in2 => \N__18290\,
            in3 => \N__19817\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23811\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_1_LC_9_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110000000110"
        )
    port map (
            in0 => \N__21973\,
            in1 => \N__17871\,
            in2 => \N__23531\,
            in3 => \N__21203\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23811\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIMKS41_10_LC_9_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001101100"
        )
    port map (
            in0 => \N__19591\,
            in1 => \N__22525\,
            in2 => \N__19706\,
            in3 => \N__21084\,
            lcout => \ppm_encoder_1.N_256_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNI70081_3_LC_9_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100011011001100"
        )
    port map (
            in0 => \N__17812\,
            in1 => \N__20587\,
            in2 => \N__21169\,
            in3 => \N__19630\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIVM131_0_16_LC_9_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001111000"
        )
    port map (
            in0 => \N__21772\,
            in1 => \N__24004\,
            in2 => \N__21271\,
            in3 => \N__21099\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_axb_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNI98UU1_2_LC_9_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100101010110"
        )
    port map (
            in0 => \N__20532\,
            in1 => \N__17744\,
            in2 => \N__21168\,
            in3 => \N__17667\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un1_init_pulses_3_axb_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIGLA33_2_LC_9_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17586\,
            in3 => \N__18039\,
            lcout => \ppm_encoder_1.init_pulses_RNIGLA33Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIROS41_14_LC_9_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001110011001100"
        )
    port map (
            in0 => \N__21097\,
            in1 => \N__21507\,
            in2 => \N__19714\,
            in3 => \N__20391\,
            lcout => \ppm_encoder_1.N_260_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIA2081_5_LC_9_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001111000"
        )
    port map (
            in0 => \N__19631\,
            in1 => \N__19701\,
            in2 => \N__22577\,
            in3 => \N__21098\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.PPM_STATE_fast_RNI4RFR_0_LC_9_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001111000"
        )
    port map (
            in0 => \N__19862\,
            in1 => \N__19818\,
            in2 => \N__20539\,
            in3 => \N__19424\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.PPM_STATE_fast_RNI4RFRZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNI7DC41_2_LC_9_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20531\,
            in2 => \N__18090\,
            in3 => \N__22837\,
            lcout => \ppm_encoder_1.N_249_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIUUR33_0_LC_9_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18087\,
            in2 => \N__20440\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_26_0_\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_1_LC_9_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18075\,
            in2 => \_gnd_net_\,
            in3 => \N__18063\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_1\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_0\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_2_LC_9_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18060\,
            in2 => \N__18047\,
            in3 => \N__18006\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_2\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_1\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_3_LC_9_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18003\,
            in2 => \_gnd_net_\,
            in3 => \N__17988\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_3\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_2\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_4_LC_9_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17985\,
            in2 => \_gnd_net_\,
            in3 => \N__17961\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_4\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_3\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_5_LC_9_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17958\,
            in2 => \_gnd_net_\,
            in3 => \N__17943\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_5\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_4\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_6_LC_9_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17940\,
            in2 => \N__17929\,
            in3 => \N__17886\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_6\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_5\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_7_LC_9_26_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19431\,
            in2 => \_gnd_net_\,
            in3 => \N__18234\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_7\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_6\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_8_LC_9_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18666\,
            in2 => \_gnd_net_\,
            in3 => \N__18222\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_8\,
            ltout => OPEN,
            carryin => \bfn_9_27_0_\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_9_LC_9_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18219\,
            in2 => \_gnd_net_\,
            in3 => \N__18207\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_9\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_8\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_10_LC_9_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18204\,
            in2 => \_gnd_net_\,
            in3 => \N__18192\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_10\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_9\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_11_LC_9_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18189\,
            in3 => \N__18174\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_11\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_10\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_12_LC_9_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18171\,
            in2 => \_gnd_net_\,
            in3 => \N__18159\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_12\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_11\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_13_LC_9_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18152\,
            in2 => \N__18120\,
            in3 => \N__18105\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_13\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_12\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_init_pulses_3_cry_13_THRU_LUT4_0_LC_9_27_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18317\,
            in3 => \N__18093\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_cry_13_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_13\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_15_LC_9_27_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20625\,
            in2 => \_gnd_net_\,
            in3 => \N__18372\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_15\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_14\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_16_LC_9_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18327\,
            in2 => \_gnd_net_\,
            in3 => \N__18357\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_16\,
            ltout => OPEN,
            carryin => \bfn_9_28_0_\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_17_LC_9_28_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18300\,
            in2 => \_gnd_net_\,
            in3 => \N__18342\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_17\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_16\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_18_LC_9_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19968\,
            in2 => \_gnd_net_\,
            in3 => \N__18339\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_2_LC_9_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001000010000"
        )
    port map (
            in0 => \N__21218\,
            in1 => \N__23522\,
            in2 => \N__18273\,
            in3 => \N__23961\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23788\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIVM131_16_LC_9_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011010011110000"
        )
    port map (
            in0 => \N__21216\,
            in1 => \N__23959\,
            in2 => \N__21272\,
            in3 => \N__21685\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNITK131_14_LC_9_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001101100"
        )
    port map (
            in0 => \N__21684\,
            in1 => \N__21511\,
            in2 => \N__24002\,
            in3 => \N__21215\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNI0O131_17_LC_9_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011010011110000"
        )
    port map (
            in0 => \N__21217\,
            in1 => \N__23960\,
            in2 => \N__20926\,
            in3 => \N__21686\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m6_0_0_LC_9_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011110001000"
        )
    port map (
            in0 => \N__22097\,
            in1 => \N__21965\,
            in2 => \N__21734\,
            in3 => \N__20396\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_ns_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m9_0_i_LC_9_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011100001111"
        )
    port map (
            in0 => \N__22096\,
            in1 => \N__21964\,
            in2 => \N__21733\,
            in3 => \N__20395\,
            lcout => \ppm_encoder_1.N_204\,
            ltout => \ppm_encoder_1.N_204_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_3_LC_9_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010000000101"
        )
    port map (
            in0 => \N__23511\,
            in1 => \N__21702\,
            in2 => \N__18597\,
            in3 => \N__21219\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23785\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_2_8_LC_10_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000001110000"
        )
    port map (
            in0 => \N__18594\,
            in1 => \N__20159\,
            in2 => \N__20273\,
            in3 => \N__18576\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.N_379_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_8_LC_10_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20419\,
            in2 => \N__18558\,
            in3 => \N__18551\,
            lcout => \ppm_encoder_1.pulses2count_9_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_7_LC_10_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010111001100"
        )
    port map (
            in0 => \N__18533\,
            in1 => \N__18516\,
            in2 => \N__18789\,
            in3 => \N__18903\,
            lcout => \ppm_encoder_1.N_302\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_3_12_LC_10_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__20420\,
            in1 => \N__18501\,
            in2 => \N__20274\,
            in3 => \N__20160\,
            lcout => \ppm_encoder_1.N_396\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_11_LC_10_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__22116\,
            in1 => \N__21975\,
            in2 => \N__18387\,
            in3 => \N__18468\,
            lcout => \ppm_encoder_1.pulses2count_9_0_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_8_LC_10_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110100"
        )
    port map (
            in0 => \N__22117\,
            in1 => \N__21976\,
            in2 => \N__18444\,
            in3 => \N__18435\,
            lcout => \ppm_encoder_1.pulses2count_9_i_1_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_3_11_LC_10_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__20158\,
            in1 => \N__18414\,
            in2 => \N__20421\,
            in3 => \N__20272\,
            lcout => \ppm_encoder_1.N_391\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_12_LC_10_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__22118\,
            in1 => \N__21991\,
            in2 => \N__19092\,
            in3 => \N__24025\,
            lcout => \ppm_encoder_1.N_393\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_RNIHVID1_1_LC_10_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011110100"
        )
    port map (
            in0 => \N__21993\,
            in1 => \N__20418\,
            in2 => \N__21786\,
            in3 => \N__22120\,
            lcout => \ppm_encoder_1.pulses2count_9_0_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_12_LC_10_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__22119\,
            in1 => \N__21992\,
            in2 => \N__19059\,
            in3 => \N__19047\,
            lcout => \ppm_encoder_1.pulses2count_9_0_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_2_9_LC_10_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__20257\,
            in1 => \N__20157\,
            in2 => \_gnd_net_\,
            in3 => \N__19014\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.N_327_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_9_LC_10_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111110"
        )
    port map (
            in0 => \N__18984\,
            in1 => \N__24024\,
            in2 => \N__18972\,
            in3 => \N__18969\,
            lcout => \ppm_encoder_1.pulses2count_9_i_0_1_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_5_LC_10_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001011100"
        )
    port map (
            in0 => \N__18939\,
            in1 => \N__18921\,
            in2 => \N__18900\,
            in3 => \N__18787\,
            lcout => \ppm_encoder_1.N_300\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNID5081_0_8_LC_10_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001111000"
        )
    port map (
            in0 => \N__19690\,
            in1 => \N__19623\,
            in2 => \N__22703\,
            in3 => \N__21089\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_3_rep2_LC_10_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001100000001"
        )
    port map (
            in0 => \N__21090\,
            in1 => \N__23520\,
            in2 => \N__18653\,
            in3 => \N__19691\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_3_repZ0Z2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23805\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNID5081_8_LC_10_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001111000"
        )
    port map (
            in0 => \N__19688\,
            in1 => \N__19622\,
            in2 => \N__22702\,
            in3 => \N__21087\,
            lcout => \ppm_encoder_1.N_255_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_2_12_LC_10_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__20828\,
            in1 => \N__19336\,
            in2 => \N__24253\,
            in3 => \N__19374\,
            lcout => \ppm_encoder_1.pulses2count_9_0_2_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIPMS41_12_LC_10_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001111000"
        )
    port map (
            in0 => \N__19689\,
            in1 => \N__20407\,
            in2 => \N__19338\,
            in3 => \N__21088\,
            lcout => \ppm_encoder_1.N_258_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIOLS41_11_LC_10_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001111000"
        )
    port map (
            in0 => \N__19687\,
            in1 => \N__20406\,
            in2 => \N__20039\,
            in3 => \N__21086\,
            lcout => \ppm_encoder_1.N_257_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_6_LC_10_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011101100"
        )
    port map (
            in0 => \N__20408\,
            in1 => \N__21781\,
            in2 => \N__21609\,
            in3 => \N__19239\,
            lcout => \ppm_encoder_1.pulses2count_9_0_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_21_c_RNO_LC_10_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__19143\,
            in1 => \N__22384\,
            in2 => \N__19128\,
            in3 => \N__22327\,
            lcout => \ppm_encoder_1.counter24_0_I_21_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_6_LC_10_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111011101110"
        )
    port map (
            in0 => \N__19209\,
            in1 => \N__19203\,
            in2 => \N__19188\,
            in3 => \N__24236\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23799\,
            ce => \N__23569\,
            sr => \N__23371\
        );

    \ppm_encoder_1.pulses2count_esr_7_LC_10_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001100000001"
        )
    port map (
            in0 => \N__24235\,
            in1 => \N__19137\,
            in2 => \N__22251\,
            in3 => \N__19471\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23799\,
            ce => \N__23569\,
            sr => \N__23371\
        );

    \ppm_encoder_1.pulses2count_esr_12_LC_10_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__21407\,
            in1 => \N__19119\,
            in2 => \N__19113\,
            in3 => \N__19101\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23799\,
            ce => \N__23569\,
            sr => \N__23371\
        );

    \ppm_encoder_1.init_pulses_RNILB4M_0_LC_10_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011010011110000"
        )
    port map (
            in0 => \N__24393\,
            in1 => \N__19861\,
            in2 => \N__22235\,
            in3 => \N__19819\,
            lcout => \ppm_encoder_1.init_pulses_RNILB4MZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIC4081_7_LC_10_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001111000"
        )
    port map (
            in0 => \N__19705\,
            in1 => \N__19621\,
            in2 => \N__19479\,
            in3 => \N__21100\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.PPM_STATE_fast_0_LC_10_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000001"
        )
    port map (
            in0 => \N__22840\,
            in1 => \N__24529\,
            in2 => \N__22872\,
            in3 => \N__24579\,
            lcout => \ppm_encoder_1.PPM_STATE_fastZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23794\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter_RNII3AF_1_LC_10_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__24345\,
            in1 => \N__22186\,
            in2 => \N__22469\,
            in3 => \N__22839\,
            lcout => \ppm_encoder_1.un1_PPM_STATE_0_sqmuxa_0_i_0_a2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter_RNIS9KG_2_LC_10_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__20753\,
            in1 => \N__20732\,
            in2 => \N__22770\,
            in3 => \N__22733\,
            lcout => \ppm_encoder_1.un1_PPM_STATE_0_sqmuxa_0_i_0_a2_16_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.PPM_STATE_0_LC_10_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000001011"
        )
    port map (
            in0 => \N__24578\,
            in1 => \N__22868\,
            in2 => \N__24534\,
            in3 => \N__22841\,
            lcout => \ppm_encoder_1.PPM_STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23794\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.PPM_STATE_1_LC_10_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__24394\,
            in1 => \N__24528\,
            in2 => \_gnd_net_\,
            in3 => \N__24577\,
            lcout => \ppm_encoder_1.PPM_STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23794\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.ppm_output_reg_RNO_1_LC_10_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__24346\,
            in1 => \N__22194\,
            in2 => \N__22470\,
            in3 => \N__24401\,
            lcout => \ppm_encoder_1.un1_PPM_STATE_1_sqmuxa_i_i_a2_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_11_LC_10_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__22072\,
            in1 => \N__21942\,
            in2 => \N__24086\,
            in3 => \N__19410\,
            lcout => \ppm_encoder_1.N_388\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIMR0V_0_LC_10_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__22231\,
            in1 => \N__20466\,
            in2 => \_gnd_net_\,
            in3 => \N__22838\,
            lcout => \ppm_encoder_1.N_247_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_1_rep2_RNI1UMR_LC_10_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__20414\,
            in1 => \N__20255\,
            in2 => \_gnd_net_\,
            in3 => \N__20143\,
            lcout => \ppm_encoder_1.N_441\,
            ltout => \ppm_encoder_1.N_441_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_2_11_LC_10_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__20816\,
            in1 => \N__20032\,
            in2 => \N__19995\,
            in3 => \N__19992\,
            lcout => \ppm_encoder_1.pulses2count_9_0_2_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter_RNIM3KG_18_LC_10_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__21450\,
            in1 => \N__22990\,
            in2 => \N__22428\,
            in3 => \N__22155\,
            lcout => \ppm_encoder_1.un1_PPM_STATE_0_sqmuxa_0_i_0_a2_2_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_3_18_LC_10_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001101100"
        )
    port map (
            in0 => \N__21761\,
            in1 => \N__20885\,
            in2 => \N__24005\,
            in3 => \N__21221\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_2_10_LC_10_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__22059\,
            in1 => \N__21980\,
            in2 => \_gnd_net_\,
            in3 => \N__19962\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.N_385_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_10_LC_10_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111100"
        )
    port map (
            in0 => \N__19932\,
            in1 => \N__19902\,
            in2 => \N__19890\,
            in3 => \N__23981\,
            lcout => \ppm_encoder_1.pulses2count_9_i_1_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_1_LC_10_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010000100110000"
        )
    port map (
            in0 => \N__21222\,
            in1 => \N__23521\,
            in2 => \N__22098\,
            in3 => \N__21981\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23786\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_2_4_LC_10_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__22058\,
            in1 => \N__21979\,
            in2 => \_gnd_net_\,
            in3 => \N__19887\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.N_371_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_4_LC_10_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111110"
        )
    port map (
            in0 => \N__20700\,
            in1 => \N__23980\,
            in2 => \N__20688\,
            in3 => \N__20685\,
            lcout => \ppm_encoder_1.pulses2count_9_i_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_13_LC_10_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011101100"
        )
    port map (
            in0 => \N__23982\,
            in1 => \N__21762\,
            in2 => \N__21621\,
            in3 => \N__20664\,
            lcout => \ppm_encoder_1.pulses2count_9_0_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_RNIIFQ91_0_1_LC_10_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101010101010"
        )
    port map (
            in0 => \N__21703\,
            in1 => \N__22068\,
            in2 => \N__24003\,
            in3 => \N__21966\,
            lcout => \ppm_encoder_1.N_247\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIUL131_15_LC_10_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001111000"
        )
    port map (
            in0 => \N__21687\,
            in1 => \N__23962\,
            in2 => \N__21830\,
            in3 => \N__21220\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_2_LC_11_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000110"
        )
    port map (
            in0 => \N__22123\,
            in1 => \N__21977\,
            in2 => \N__24085\,
            in3 => \N__20619\,
            lcout => \ppm_encoder_1.N_360\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_3_LC_11_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111011111010"
        )
    port map (
            in0 => \N__20472\,
            in1 => \N__24255\,
            in2 => \N__20502\,
            in3 => \N__20592\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23806\,
            ce => \N__23564\,
            sr => \N__23366\
        );

    \ppm_encoder_1.pulses2count_esr_2_LC_11_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001010001"
        )
    port map (
            in0 => \N__20556\,
            in1 => \N__24260\,
            in2 => \N__20547\,
            in3 => \N__20501\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23800\,
            ce => \N__23567\,
            sr => \N__23372\
        );

    \ppm_encoder_1.counter24_0_I_9_c_RNO_LC_11_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__20731\,
            in1 => \N__20487\,
            in2 => \N__20481\,
            in3 => \N__20752\,
            lcout => \ppm_encoder_1.counter24_0_I_9_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_3_LC_11_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011000000010"
        )
    port map (
            in0 => \N__22124\,
            in1 => \N__21978\,
            in2 => \N__24089\,
            in3 => \N__20777\,
            lcout => \ppm_encoder_1.N_365\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_1_LC_11_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111011111010"
        )
    port map (
            in0 => \N__21408\,
            in1 => \N__20829\,
            in2 => \N__20793\,
            in3 => \N__20778\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23800\,
            ce => \N__23567\,
            sr => \N__23372\
        );

    \ppm_encoder_1.counter_0_LC_11_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22154\,
            in2 => \N__21227\,
            in3 => \N__21201\,
            lcout => \ppm_encoder_1.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_11_24_0_\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_0\,
            clk => \N__23795\,
            ce => 'H',
            sr => \N__21423\
        );

    \ppm_encoder_1.counter_1_LC_11_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22187\,
            in2 => \_gnd_net_\,
            in3 => \N__20757\,
            lcout => \ppm_encoder_1.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_0\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_1\,
            clk => \N__23795\,
            ce => 'H',
            sr => \N__21423\
        );

    \ppm_encoder_1.counter_2_LC_11_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20754\,
            in2 => \_gnd_net_\,
            in3 => \N__20736\,
            lcout => \ppm_encoder_1.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_1\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_2\,
            clk => \N__23795\,
            ce => 'H',
            sr => \N__21423\
        );

    \ppm_encoder_1.counter_3_LC_11_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20733\,
            in2 => \_gnd_net_\,
            in3 => \N__20715\,
            lcout => \ppm_encoder_1.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_2\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_3\,
            clk => \N__23795\,
            ce => 'H',
            sr => \N__21423\
        );

    \ppm_encoder_1.counter_4_LC_11_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21449\,
            in2 => \_gnd_net_\,
            in3 => \N__20712\,
            lcout => \ppm_encoder_1.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_3\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_4\,
            clk => \N__23795\,
            ce => 'H',
            sr => \N__21423\
        );

    \ppm_encoder_1.counter_5_LC_11_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22368\,
            in2 => \_gnd_net_\,
            in3 => \N__20709\,
            lcout => \ppm_encoder_1.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_4\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_5\,
            clk => \N__23795\,
            ce => 'H',
            sr => \N__21423\
        );

    \ppm_encoder_1.counter_6_LC_11_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22329\,
            in2 => \_gnd_net_\,
            in3 => \N__20706\,
            lcout => \ppm_encoder_1.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_5\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_6\,
            clk => \N__23795\,
            ce => 'H',
            sr => \N__21423\
        );

    \ppm_encoder_1.counter_7_LC_11_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22386\,
            in2 => \_gnd_net_\,
            in3 => \N__20703\,
            lcout => \ppm_encoder_1.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_6\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_7\,
            clk => \N__23795\,
            ce => 'H',
            sr => \N__21423\
        );

    \ppm_encoder_1.counter_8_LC_11_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24299\,
            in2 => \_gnd_net_\,
            in3 => \N__20856\,
            lcout => \ppm_encoder_1.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_11_25_0_\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_8\,
            clk => \N__23790\,
            ce => 'H',
            sr => \N__21422\
        );

    \ppm_encoder_1.counter_9_LC_11_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24347\,
            in2 => \_gnd_net_\,
            in3 => \N__20853\,
            lcout => \ppm_encoder_1.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_8\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_9\,
            clk => \N__23790\,
            ce => 'H',
            sr => \N__21422\
        );

    \ppm_encoder_1.counter_10_LC_11_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22427\,
            in2 => \_gnd_net_\,
            in3 => \N__20850\,
            lcout => \ppm_encoder_1.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_9\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_10\,
            clk => \N__23790\,
            ce => 'H',
            sr => \N__21422\
        );

    \ppm_encoder_1.counter_11_LC_11_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22468\,
            in2 => \_gnd_net_\,
            in3 => \N__20847\,
            lcout => \ppm_encoder_1.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_10\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_11\,
            clk => \N__23790\,
            ce => 'H',
            sr => \N__21422\
        );

    \ppm_encoder_1.counter_12_LC_11_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23019\,
            in2 => \_gnd_net_\,
            in3 => \N__20844\,
            lcout => \ppm_encoder_1.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_11\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_12\,
            clk => \N__23790\,
            ce => 'H',
            sr => \N__21422\
        );

    \ppm_encoder_1.counter_13_LC_11_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22938\,
            in2 => \_gnd_net_\,
            in3 => \N__20841\,
            lcout => \ppm_encoder_1.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_12\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_13\,
            clk => \N__23790\,
            ce => 'H',
            sr => \N__21422\
        );

    \ppm_encoder_1.counter_14_LC_11_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22349\,
            in2 => \_gnd_net_\,
            in3 => \N__20838\,
            lcout => \ppm_encoder_1.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_13\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_14\,
            clk => \N__23790\,
            ce => 'H',
            sr => \N__21422\
        );

    \ppm_encoder_1.counter_15_LC_11_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22968\,
            in2 => \_gnd_net_\,
            in3 => \N__20835\,
            lcout => \ppm_encoder_1.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_14\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_15\,
            clk => \N__23790\,
            ce => 'H',
            sr => \N__21422\
        );

    \ppm_encoder_1.counter_16_LC_11_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22734\,
            in2 => \_gnd_net_\,
            in3 => \N__20832\,
            lcout => \ppm_encoder_1.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_11_26_0_\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_16\,
            clk => \N__23787\,
            ce => 'H',
            sr => \N__21421\
        );

    \ppm_encoder_1.counter_17_LC_11_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22766\,
            in2 => \_gnd_net_\,
            in3 => \N__21429\,
            lcout => \ppm_encoder_1.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_16\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_17\,
            clk => \N__23787\,
            ce => 'H',
            sr => \N__21421\
        );

    \ppm_encoder_1.counter_18_LC_11_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22994\,
            in2 => \_gnd_net_\,
            in3 => \N__21426\,
            lcout => \ppm_encoder_1.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23787\,
            ce => 'H',
            sr => \N__21421\
        );

    \ppm_encoder_1.pulses2count_esr_11_LC_11_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__21394\,
            in1 => \N__21381\,
            in2 => \N__21375\,
            in3 => \N__21366\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23784\,
            ce => \N__23570\,
            sr => \N__23396\
        );

    \ppm_encoder_1.pulses2count_esr_13_LC_11_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__24225\,
            in1 => \N__21350\,
            in2 => \N__21303\,
            in3 => \N__21294\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23784\,
            ce => \N__23570\,
            sr => \N__23396\
        );

    \ppm_encoder_1.pulses2count_esr_16_LC_11_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__24017\,
            in1 => \N__21622\,
            in2 => \N__21276\,
            in3 => \N__21760\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23782\,
            ce => \N__23571\,
            sr => \N__23401\
        );

    \ppm_encoder_1.PPM_STATE_fast_RNI9VGK_0_LC_12_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23490\,
            in2 => \_gnd_net_\,
            in3 => \N__21234\,
            lcout => \ppm_encoder_1.N_238_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_17_LC_12_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__24068\,
            in1 => \N__20930\,
            in2 => \N__21624\,
            in3 => \N__21777\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23798\,
            ce => \N__23562\,
            sr => \N__23373\
        );

    \ppm_encoder_1.pulses2count_esr_18_LC_12_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__21776\,
            in1 => \N__21614\,
            in2 => \N__20889\,
            in3 => \N__24069\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23798\,
            ce => \N__23562\,
            sr => \N__23373\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_5_LC_12_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011101110"
        )
    port map (
            in0 => \N__24067\,
            in1 => \N__21775\,
            in2 => \N__21623\,
            in3 => \N__22311\,
            lcout => \ppm_encoder_1.pulses2count_9_i_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_7_LC_12_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010101110"
        )
    port map (
            in0 => \N__21774\,
            in1 => \N__24066\,
            in2 => \N__22287\,
            in3 => \N__21610\,
            lcout => \ppm_encoder_1.pulses2count_9_i_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_0_LC_12_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111010"
        )
    port map (
            in0 => \N__21989\,
            in1 => \N__24073\,
            in2 => \N__22133\,
            in3 => \N__22236\,
            lcout => \ppm_encoder_1.pulses2count_9_0_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_1_c_RNO_LC_12_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__22185\,
            in1 => \N__23889\,
            in2 => \N__22164\,
            in3 => \N__22150\,
            lcout => \ppm_encoder_1.counter24_0_I_1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_RNIIFQ91_1_LC_12_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011101010"
        )
    port map (
            in0 => \N__21778\,
            in1 => \N__22125\,
            in2 => \N__24087\,
            in3 => \N__21990\,
            lcout => \ppm_encoder_1.N_244\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_15_LC_12_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__21619\,
            in1 => \N__21780\,
            in2 => \N__21831\,
            in3 => \N__24077\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23793\,
            ce => \N__23563\,
            sr => \N__23380\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_14_LC_12_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011111010"
        )
    port map (
            in0 => \N__21779\,
            in1 => \N__21618\,
            in2 => \N__24088\,
            in3 => \N__21539\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.pulses2count_9_i_0_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_14_LC_12_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000001011"
        )
    port map (
            in0 => \N__21513\,
            in1 => \N__24261\,
            in2 => \N__21471\,
            in3 => \N__21468\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23793\,
            ce => \N__23563\,
            sr => \N__23380\
        );

    \ppm_encoder_1.counter24_0_I_15_c_RNO_LC_12_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__22366\,
            in1 => \N__22608\,
            in2 => \N__22539\,
            in3 => \N__21445\,
            lcout => \ppm_encoder_1.counter24_0_I_15_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_4_LC_12_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100000001"
        )
    port map (
            in0 => \N__22656\,
            in1 => \N__24259\,
            in2 => \N__24125\,
            in3 => \N__22644\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23789\,
            ce => \N__23566\,
            sr => \N__23386\
        );

    \ppm_encoder_1.pulses2count_esr_5_LC_12_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001100000001"
        )
    port map (
            in0 => \N__24257\,
            in1 => \N__22602\,
            in2 => \N__22590\,
            in3 => \N__22578\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23789\,
            ce => \N__23566\,
            sr => \N__23386\
        );

    \ppm_encoder_1.pulses2count_esr_10_LC_12_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001010001"
        )
    port map (
            in0 => \N__24118\,
            in1 => \N__24258\,
            in2 => \N__22530\,
            in3 => \N__22488\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23789\,
            ce => \N__23566\,
            sr => \N__23386\
        );

    \ppm_encoder_1.counter24_0_I_33_c_RNO_LC_12_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__22476\,
            in1 => \N__22461\,
            in2 => \N__22440\,
            in3 => \N__22423\,
            lcout => \ppm_encoder_1.counter24_0_I_33_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_57_c_RNIJMMD_LC_12_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__24554\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24407\,
            lcout => \ppm_encoder_1.counter24_0_I_57_c_RNIJMMDZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_45_c_RNO_LC_12_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__22966\,
            in1 => \N__22407\,
            in2 => \N__22398\,
            in3 => \N__22345\,
            lcout => \ppm_encoder_1.counter24_0_I_45_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter_RNIGV08_5_LC_12_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22385\,
            in2 => \_gnd_net_\,
            in3 => \N__22367\,
            lcout => \ppm_encoder_1.un1_PPM_STATE_0_sqmuxa_0_i_0_a2_2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter_RNIUBKG_6_LC_12_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__23018\,
            in1 => \N__24298\,
            in2 => \N__22350\,
            in3 => \N__22328\,
            lcout => \ppm_encoder_1.un1_PPM_STATE_0_sqmuxa_0_i_0_a2_16_4\,
            ltout => \ppm_encoder_1.un1_PPM_STATE_0_sqmuxa_0_i_0_a2_16_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter_RNI09RH2_1_LC_12_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22895\,
            in1 => \N__23055\,
            in2 => \N__23046\,
            in3 => \N__22920\,
            lcout => \ppm_encoder_1.N_330\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_39_c_RNO_LC_12_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__23043\,
            in1 => \N__22936\,
            in2 => \N__23031\,
            in3 => \N__23017\,
            lcout => \ppm_encoder_1.counter24_0_I_39_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_57_c_RNO_LC_12_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23004\,
            in2 => \_gnd_net_\,
            in3 => \N__22995\,
            lcout => \ppm_encoder_1.counter24_0_I_57_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter_RNIKF811_13_LC_12_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__22974\,
            in1 => \N__22967\,
            in2 => \N__22950\,
            in3 => \N__22937\,
            lcout => \ppm_encoder_1.un1_PPM_STATE_0_sqmuxa_0_i_0_a2_2\,
            ltout => \ppm_encoder_1.un1_PPM_STATE_0_sqmuxa_0_i_0_a2_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.ppm_output_reg_RNO_0_LC_12_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22914\,
            in1 => \N__22905\,
            in2 => \N__22899\,
            in3 => \N__22896\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.N_431_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.ppm_output_reg_LC_12_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010001110101011"
        )
    port map (
            in0 => \N__22787\,
            in1 => \N__22862\,
            in2 => \N__22851\,
            in3 => \N__22848\,
            lcout => ppm_output_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23783\,
            ce => 'H',
            sr => \N__23397\
        );

    \ppm_encoder_1.counter24_0_I_51_c_RNO_LC_12_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__22776\,
            in1 => \N__22762\,
            in2 => \N__22746\,
            in3 => \N__22732\,
            lcout => \ppm_encoder_1.counter24_0_I_51_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_8_LC_13_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001100000001"
        )
    port map (
            in0 => \N__24254\,
            in1 => \N__22716\,
            in2 => \N__24126\,
            in3 => \N__22704\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23807\,
            ce => \N__23565\,
            sr => \N__23381\
        );

    \ppm_encoder_1.pulses2count_esr_9_LC_13_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001010001"
        )
    port map (
            in0 => \N__24273\,
            in1 => \N__24256\,
            in2 => \N__24165\,
            in3 => \N__24117\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23801\,
            ce => \N__23568\,
            sr => \N__23387\
        );

    \ppm_encoder_1.pulses2count_esr_0_LC_13_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__24116\,
            in1 => \N__24096\,
            in2 => \_gnd_net_\,
            in3 => \N__24078\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23801\,
            ce => \N__23568\,
            sr => \N__23387\
        );

    \ppm_encoder_1.counter24_0_I_1_c_LC_13_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23094\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_13_24_0_\,
            carryout => \ppm_encoder_1.counter24_0_data_tmp_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_9_c_LC_13_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23088\,
            in2 => \N__24747\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ppm_encoder_1.counter24_0_data_tmp_0\,
            carryout => \ppm_encoder_1.counter24_0_data_tmp_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_15_c_LC_13_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23076\,
            in2 => \N__24741\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ppm_encoder_1.counter24_0_data_tmp_1\,
            carryout => \ppm_encoder_1.counter24_0_data_tmp_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_21_c_LC_13_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23070\,
            in2 => \N__24744\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ppm_encoder_1.counter24_0_data_tmp_2\,
            carryout => \ppm_encoder_1.counter24_0_data_tmp_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_27_c_LC_13_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24279\,
            in2 => \N__24742\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ppm_encoder_1.counter24_0_data_tmp_3\,
            carryout => \ppm_encoder_1.counter24_0_data_tmp_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_33_c_LC_13_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23061\,
            in2 => \N__24745\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ppm_encoder_1.counter24_0_data_tmp_4\,
            carryout => \ppm_encoder_1.counter24_0_data_tmp_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_39_c_LC_13_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24801\,
            in2 => \N__24743\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ppm_encoder_1.counter24_0_data_tmp_5\,
            carryout => \ppm_encoder_1.counter24_0_data_tmp_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_45_c_LC_13_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24795\,
            in2 => \N__24746\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ppm_encoder_1.counter24_0_data_tmp_6\,
            carryout => \ppm_encoder_1.counter24_0_data_tmp_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_51_c_LC_13_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24712\,
            in2 => \N__24789\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_13_25_0_\,
            carryout => \ppm_encoder_1.counter24_0_data_tmp_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_57_c_LC_13_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24777\,
            in2 => \N__24748\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ppm_encoder_1.counter24_0_data_tmp_8\,
            carryout => \ppm_encoder_1.counter24_0_N_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_N_2_THRU_LUT4_0_LC_13_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24582\,
            lcout => \ppm_encoder_1.counter24_0_N_2_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_57_c_RNIGCO83_LC_13_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111010"
        )
    port map (
            in0 => \N__24569\,
            in1 => \N__24550\,
            in2 => \N__24533\,
            in3 => \N__24406\,
            lcout => \ppm_encoder_1.counter24_0_I_57_c_RNIGCOZ0Z83\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_27_c_RNO_LC_13_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__24348\,
            in1 => \N__24321\,
            in2 => \N__24312\,
            in3 => \N__24300\,
            lcout => \ppm_encoder_1.counter24_0_I_27_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
